module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[11:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[63:0] pcr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  reg [2:0] state;
  wire[2:0] T363;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire[3:0] rx_cmd;
  reg [3:0] cmd;
  wire[3:0] T19;
  wire T20;
  wire T21;
  reg [14:0] rx_count;
  wire[14:0] T364;
  wire[14:0] T22;
  wire[14:0] T23;
  wire[14:0] T24;
  wire T25;
  wire T26;
  wire[12:0] T365;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T27;
  wire[11:0] T28;
  wire[63:0] rx_shifter_in;
  wire[47:0] T29;
  reg [63:0] rx_shifter;
  wire[63:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire nack;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire bad_mem_packet;
  wire T43;
  wire[2:0] T44;
  reg [39:0] addr;
  wire[39:0] T45;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire[39:0] T50;
  wire T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T366;
  wire[14:0] T56;
  wire[14:0] T57;
  wire[14:0] T58;
  wire T59;
  wire T60;
  wire[3:0] next_cmd;
  wire T61;
  wire[12:0] rx_word_count;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire rx_done;
  wire T66;
  wire T67;
  wire T68;
  wire[2:0] T69;
  wire T70;
  wire[12:0] T367;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire rx_word_done;
  wire T75;
  wire[1:0] T76;
  wire T77;
  wire T78;
  wire cnt_done;
  wire T79;
  reg [1:0] cnt;
  wire[1:0] T368;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire[2:0] T90;
  wire T91;
  wire T92;
  reg [8:0] pos;
  wire[8:0] T93;
  wire[8:0] T94;
  wire[8:0] T95;
  wire[8:0] T96;
  wire[8:0] T97;
  wire[8:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire[2:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[2:0] T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire tx_done;
  wire T113;
  wire T114;
  wire T115;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire[12:0] T369;
  wire T119;
  wire T120;
  wire[1:0] tx_subword_count;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[11:0] pcr_addr;
  wire T127;
  wire T128;
  wire[1:0] pcr_coreid;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire[2:0] T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire T138;
  wire T139;
  wire[2:0] T140;
  wire[63:0] T141;
  wire T142;
  wire[2:0] T143;
  wire[2:0] T144;
  wire[5:0] T145;
  wire[5:0] scr_addr;
  wire T146;
  wire T147;
  wire[16:0] T148;
  wire[16:0] T149;
  wire[16:0] T150;
  wire[16:0] T151;
  wire[15:0] T152;
  wire T153;
  wire[2:0] T154;
  wire[2:0] T155;
  wire[2:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire[127:0] T160;
  wire[127:0] T161;
  wire[127:0] T162;
  wire[127:0] mem_req_data;
  wire[63:0] T163;
  wire[2:0] T164;
  wire[63:0] T165;
  wire[2:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire[1:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire[25:0] T173;
  wire[25:0] T174;
  wire[25:0] T370;
  wire[36:0] init_addr;
  wire[39:0] T175;
  wire[25:0] T176;
  wire[25:0] T371;
  wire T177;
  wire T178;
  wire T179;
  reg  R180;
  wire T372;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[63:0] T185;
  reg [63:0] rtc;
  wire[63:0] T373;
  wire[63:0] T186;
  wire[63:0] T187;
  wire rtc_tick;
  reg [6:0] R188;
  wire[6:0] T374;
  wire[6:0] T189;
  wire[6:0] T190;
  wire T191;
  wire T192;
  reg  R193;
  wire T375;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg  R198;
  wire T376;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[11:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  reg  R213;
  wire T377;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire[15:0] T378;
  wire[63:0] T218;
  wire[5:0] T219;
  wire[1:0] T220;
  wire[63:0] tx_data;
  wire[63:0] T221;
  wire[63:0] T222;
  reg [63:0] pcrReadData;
  wire[63:0] T223;
  wire[63:0] T224;
  wire[63:0] T225;
  wire[63:0] T379;
  wire[63:0] T226;
  wire[63:0] T227;
  wire[63:0] T228;
  wire[63:0] T229;
  wire[63:0] T230;
  wire[63:0] T231;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T232;
  wire[5:0] T233;
  wire[63:0] T234;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T235;
  wire T236;
  wire[63:0] T237;
  wire[63:0] T238;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T239;
  wire[63:0] T240;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T241;
  wire T242;
  wire T243;
  wire[63:0] T244;
  wire[63:0] T245;
  wire[63:0] T246;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T247;
  wire[63:0] T248;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T249;
  wire T250;
  wire[63:0] T251;
  wire[63:0] T252;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T253;
  wire[63:0] T254;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire[63:0] T259;
  wire[63:0] T260;
  wire[63:0] T261;
  wire[63:0] T262;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T263;
  wire[63:0] T264;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T265;
  wire T266;
  wire[63:0] T267;
  wire[63:0] T268;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T269;
  wire[63:0] T270;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T271;
  wire T272;
  wire T273;
  wire[63:0] T274;
  wire[63:0] T275;
  wire[63:0] T276;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T277;
  wire[63:0] T278;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T279;
  wire T280;
  wire[63:0] T281;
  wire[63:0] T282;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T283;
  wire[63:0] T284;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire[63:0] T290;
  wire[63:0] T291;
  wire[63:0] T292;
  wire[63:0] T293;
  wire[63:0] T294;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T295;
  wire[63:0] T296;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T297;
  wire T298;
  wire[63:0] T299;
  wire[63:0] T300;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T301;
  wire[63:0] T302;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T303;
  wire T304;
  wire T305;
  wire[63:0] T306;
  wire[63:0] T307;
  wire[63:0] T308;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T309;
  wire[63:0] T310;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T311;
  wire T312;
  wire[63:0] T313;
  wire[63:0] T314;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T315;
  wire[63:0] T316;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[63:0] T321;
  wire[63:0] T322;
  wire[63:0] T323;
  wire[63:0] T324;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T325;
  wire[63:0] T326;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T327;
  wire T328;
  wire[63:0] T329;
  wire[63:0] T330;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T331;
  wire[63:0] T332;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T333;
  wire T334;
  wire T335;
  wire[63:0] T336;
  wire[63:0] T337;
  wire[63:0] T338;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T339;
  wire[63:0] T340;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T341;
  wire T342;
  wire[63:0] T343;
  wire[63:0] T344;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T345;
  wire[63:0] T346;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire[63:0] tx_header;
  wire[15:0] T356;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T357;
  reg [7:0] seqno;
  wire[7:0] T358;
  wire[7:0] T359;
  wire T360;
  wire T361;
  wire T362;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    state = {1{$random}};
    cmd = {1{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    rx_shifter = {2{$random}};
    addr = {2{$random}};
    tx_count = {1{$random}};
    cnt = {1{$random}};
    pos = {1{$random}};
    R180 = {1{$random}};
    rtc = {2{$random}};
    R188 = {1{$random}};
    R193 = {1{$random}};
    R198 = {1{$random}};
    R213 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_cpu_0_ipi_rep_bits = {1{$random}};
//  assign io_cpu_0_id = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_scr_wdata = pcr_wdata;
  assign pcr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_data[7'h7f:7'h40];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 3'h5;
  assign T363 = reset ? 3'h0 : T4;
  assign T4 = T132 ? 3'h7 : T5;
  assign T5 = T130 ? 3'h7 : T6;
  assign T6 = T125 ? 3'h7 : T7;
  assign T7 = T122 ? 3'h2 : T8;
  assign T8 = T112 ? T108 : T9;
  assign T9 = T106 ? T102 : T10;
  assign T10 = T100 ? T90 : T11;
  assign T11 = T88 ? 3'h5 : T12;
  assign T12 = T78 ? 3'h6 : T13;
  assign T13 = T65 ? T14 : state;
  assign T14 = T64 ? 3'h3 : T15;
  assign T15 = T63 ? 3'h4 : T16;
  assign T16 = T17 ? 3'h1 : 3'h7;
  assign T17 = T62 | T18;
  assign T18 = rx_cmd == 4'h3;
  assign rx_cmd = T61 ? next_cmd : cmd;
  assign T19 = T20 ? next_cmd : cmd;
  assign T20 = T60 & T21;
  assign T21 = rx_count == 15'h3;
  assign T364 = reset ? 15'h0 : T22;
  assign T22 = T25 ? 15'h0 : T23;
  assign T23 = T60 ? T24 : rx_count;
  assign T24 = rx_count + 15'h1;
  assign T25 = T112 & T26;
  assign T26 = tx_word_count == T365;
  assign T365 = {1'h0, tx_size};
  assign tx_size = T31 ? size : 12'h0;
  assign T27 = T20 ? T28 : size;
  assign T28 = rx_shifter_in[4'hf:3'h4];
  assign rx_shifter_in = {io_host_in_bits, T29};
  assign T29 = rx_shifter[6'h3f:5'h10];
  assign T30 = T60 ? rx_shifter_in : rx_shifter;
  assign T31 = T37 & T32;
  assign T32 = T34 | T33;
  assign T33 = cmd == 4'h3;
  assign T34 = T36 | T35;
  assign T35 = cmd == 4'h2;
  assign T36 = cmd == 4'h0;
  assign T37 = nack ^ 1'h1;
  assign nack = T53 ? bad_mem_packet : T38;
  assign T38 = T40 ? T39 : 1'h1;
  assign T39 = size != 12'h1;
  assign T40 = T42 | T41;
  assign T41 = cmd == 4'h3;
  assign T42 = cmd == 4'h2;
  assign bad_mem_packet = T51 | T43;
  assign T43 = T44 != 3'h0;
  assign T44 = addr[2'h2:1'h0];
  assign T45 = T106 ? T50 : T46;
  assign T46 = T100 ? T49 : T47;
  assign T47 = T20 ? T48 : addr;
  assign T48 = rx_shifter_in[6'h3f:5'h18];
  assign T49 = addr + 40'h8;
  assign T50 = addr + 40'h8;
  assign T51 = T52 != 3'h0;
  assign T52 = size[2'h2:1'h0];
  assign T53 = T55 | T54;
  assign T54 = cmd == 4'h1;
  assign T55 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T366 = reset ? 15'h0 : T56;
  assign T56 = T25 ? 15'h0 : T57;
  assign T57 = T59 ? T58 : tx_count;
  assign T58 = tx_count + 15'h1;
  assign T59 = io_host_out_valid & io_host_out_ready;
  assign T60 = io_host_in_valid & io_host_in_ready;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign T61 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T62 = rx_cmd == 4'h2;
  assign T63 = rx_cmd == 4'h1;
  assign T64 = rx_cmd == 4'h0;
  assign T65 = T77 & rx_done;
  assign rx_done = rx_word_done & T66;
  assign T66 = T74 ? T71 : T67;
  assign T67 = T70 | T68;
  assign T68 = T69 == 3'h0;
  assign T69 = rx_word_count[2'h2:1'h0];
  assign T70 = rx_word_count == T367;
  assign T367 = {1'h0, size};
  assign T71 = T73 & T72;
  assign T72 = next_cmd != 4'h3;
  assign T73 = next_cmd != 4'h1;
  assign T74 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T75;
  assign T75 = T76 == 2'h3;
  assign T76 = rx_count[1'h1:1'h0];
  assign T77 = state == 3'h0;
  assign T78 = T87 & cnt_done;
  assign cnt_done = T82 & T79;
  assign T79 = cnt == 2'h3;
  assign T368 = reset ? 2'h0 : T80;
  assign T80 = T82 ? T81 : cnt;
  assign T81 = cnt + 2'h1;
  assign T82 = T85 | T83;
  assign T83 = T84 & io_mem_grant_valid;
  assign T84 = state == 3'h5;
  assign T85 = T86 & io_mem_acquire_ready;
  assign T86 = state == 3'h4;
  assign T87 = state == 3'h4;
  assign T88 = T89 & io_mem_acquire_ready;
  assign T89 = state == 3'h3;
  assign T90 = T91 ? 3'h7 : 3'h0;
  assign T91 = T99 | T92;
  assign T92 = pos == 9'h1;
  assign T93 = T106 ? T98 : T94;
  assign T94 = T100 ? T97 : T95;
  assign T95 = T20 ? T96 : pos;
  assign T96 = rx_shifter_in[4'hf:3'h7];
  assign T97 = pos - 9'h1;
  assign T98 = pos - 9'h1;
  assign T99 = cmd == 4'h0;
  assign T100 = T101 & io_mem_grant_valid;
  assign T101 = state == 3'h6;
  assign T102 = T103 ? 3'h7 : 3'h0;
  assign T103 = T105 | T104;
  assign T104 = pos == 9'h1;
  assign T105 = cmd == 4'h0;
  assign T106 = T107 & cnt_done;
  assign T107 = state == 3'h5;
  assign T108 = T109 ? 3'h3 : 3'h0;
  assign T109 = T111 & T110;
  assign T110 = pos != 9'h0;
  assign T111 = cmd == 4'h0;
  assign T112 = T121 & tx_done;
  assign tx_done = T119 & T113;
  assign T113 = T118 | T114;
  assign T114 = T117 & T115;
  assign T115 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T116 - 3'h1;
  assign T116 = tx_word_count[2'h2:1'h0];
  assign T117 = 13'h0 < tx_word_count;
  assign T118 = tx_word_count == T369;
  assign T369 = {1'h0, tx_size};
  assign T119 = io_host_out_ready & T120;
  assign T120 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T121 = state == 3'h7;
  assign T122 = T124 & T123;
  assign T123 = io_cpu_0_pcr_req_ready & io_cpu_0_pcr_req_valid;
  assign T124 = state == 3'h1;
  assign T125 = T127 & T126;
  assign T126 = pcr_addr == 12'h782;
  assign pcr_addr = addr[4'hb:1'h0];
  assign T127 = T129 & T128;
  assign T128 = pcr_coreid == 2'h0;
  assign pcr_coreid = addr[5'h15:5'h14];
  assign T129 = state == 3'h1;
  assign T130 = T131 & io_cpu_0_pcr_rep_valid;
  assign T131 = state == 3'h2;
  assign T132 = T134 & T133;
  assign T133 = pcr_coreid == 2'h3;
  assign T134 = state == 3'h1;
  assign T135 = {io_mem_grant_bits_addr_beat, 1'h1};
  assign T137 = io_mem_grant_bits_data[6'h3f:1'h0];
  assign T138 = T139 & io_mem_grant_valid;
  assign T139 = state == 3'h5;
  assign T140 = {io_mem_grant_bits_addr_beat, 1'h0};
  assign T142 = rx_word_done & io_host_in_ready;
  assign T143 = T144 - 3'h1;
  assign T144 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T145;
  assign T145 = scr_addr;
  assign scr_addr = addr[3'h5:1'h0];
  assign io_scr_wen = T146;
  assign T146 = T132 ? T147 : 1'h0;
  assign T147 = cmd == 4'h3;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_union = T148;
  assign T148 = T153 ? T150 : T149;
  assign T149 = 17'h1c1;
  assign T150 = T151;
  assign T151 = {T152, 1'h1};
  assign T152 = 16'hffff;
  assign T153 = cmd == 4'h1;
  assign io_mem_acquire_bits_a_type = T154;
  assign T154 = T153 ? T156 : T155;
  assign T155 = 3'h1;
  assign T156 = 3'h3;
  assign io_mem_acquire_bits_is_builtin_type = T157;
  assign T157 = T153 ? T159 : T158;
  assign T158 = 1'h1;
  assign T159 = 1'h1;
  assign io_mem_acquire_bits_data = T160;
  assign T160 = T153 ? T162 : T161;
  assign T161 = 128'h0;
  assign T162 = mem_req_data;
  assign mem_req_data = {T165, T163};
  assign T163 = packet_ram[T164];
  assign T164 = {cnt, 1'h0};
  assign T165 = packet_ram[T166];
  assign T166 = {cnt, 1'h1};
  assign io_mem_acquire_bits_addr_beat = T167;
  assign T167 = T153 ? T169 : T168;
  assign T168 = 2'h0;
  assign T169 = cnt;
  assign io_mem_acquire_bits_client_xact_id = T170;
  assign T170 = T153 ? T172 : T171;
  assign T171 = 1'h0;
  assign T172 = 1'h0;
  assign io_mem_acquire_bits_addr_block = T173;
  assign T173 = T153 ? T176 : T174;
  assign T174 = T370;
  assign T370 = init_addr[5'h19:1'h0];
  assign init_addr = T175 >> 2'h3;
  assign T175 = addr;
  assign T176 = T371;
  assign T371 = init_addr[5'h19:1'h0];
  assign io_mem_acquire_valid = T177;
  assign T177 = T179 | T178;
  assign T178 = state == 3'h4;
  assign T179 = state == 3'h3;
  assign io_cpu_0_ipi_rep_valid = R180;
  assign T372 = reset ? 1'h0 : T181;
  assign T181 = T183 ? 1'h1 : T182;
  assign T182 = io_cpu_0_ipi_rep_ready ? 1'h0 : R180;
  assign T183 = io_cpu_0_ipi_req_valid & T184;
  assign T184 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = T185;
  assign T185 = T191 ? rtc : pcr_wdata;
  assign T373 = reset ? 64'h0 : T186;
  assign T186 = rtc_tick ? T187 : rtc;
  assign T187 = rtc + 64'h1;
  assign rtc_tick = R188 == 7'h63;
  assign T374 = reset ? 7'h0 : T189;
  assign T189 = rtc_tick ? 7'h0 : T190;
  assign T190 = R188 + 7'h1;
  assign T191 = T196 & T192;
  assign T192 = R193 ^ 1'h1;
  assign T375 = reset ? 1'h0 : T194;
  assign T194 = T191 ? io_cpu_0_pcr_req_ready : T195;
  assign T195 = io_cpu_0_pcr_rep_valid ? 1'h0 : R193;
  assign T196 = T201 & T197;
  assign T197 = R198 ^ 1'h1;
  assign T376 = reset ? 1'h0 : T199;
  assign T199 = T191 ? io_cpu_0_pcr_req_ready : T200;
  assign T200 = rtc_tick ? 1'h0 : R198;
  assign T201 = T203 & T202;
  assign T202 = state != 3'h2;
  assign T203 = state != 3'h1;
  assign io_cpu_0_pcr_req_bits_addr = T204;
  assign T204 = T191 ? 12'h782 : pcr_addr;
  assign io_cpu_0_pcr_req_bits_rw = T205;
  assign T205 = T191 ? 1'h1 : T206;
  assign T206 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T207;
  assign T207 = T191 ? 1'h1 : T208;
  assign T208 = R193 ? 1'h0 : T209;
  assign T209 = T211 & T210;
  assign T210 = pcr_addr != 12'h782;
  assign T211 = T212 & T128;
  assign T212 = state == 3'h1;
  assign io_cpu_0_reset = R213;
  assign T377 = reset ? 1'h1 : T214;
  assign T214 = T216 ? T215 : R213;
  assign T215 = pcr_wdata[1'h0:1'h0];
  assign T216 = T125 & T217;
  assign T217 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T378;
  assign T378 = T218[4'hf:1'h0];
  assign T218 = tx_data >> T219;
  assign T219 = {T220, 4'h0};
  assign T220 = tx_count[1'h1:1'h0];
  assign tx_data = T360 ? tx_header : T221;
  assign T221 = T353 ? pcrReadData : T222;
  assign T222 = packet_ram[packet_ram_raddr];
  assign T223 = T132 ? T226 : T224;
  assign T224 = T130 ? io_cpu_0_pcr_rep_bits : T225;
  assign T225 = T125 ? T379 : pcrReadData;
  assign T379 = {63'h0, R213};
  assign T226 = T352 ? T290 : T227;
  assign T227 = T289 ? T259 : T228;
  assign T228 = T258 ? T244 : T229;
  assign T229 = T243 ? T237 : T230;
  assign T230 = T236 ? T234 : T231;
  assign T231 = T232 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T232 = T233[1'h0:1'h0];
  assign T233 = scr_addr;
  assign T234 = T235 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T235 = T233[1'h0:1'h0];
  assign T236 = T233[1'h1:1'h1];
  assign T237 = T242 ? T240 : T238;
  assign T238 = T239 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T239 = T233[1'h0:1'h0];
  assign T240 = T241 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T241 = T233[1'h0:1'h0];
  assign T242 = T233[1'h1:1'h1];
  assign T243 = T233[2'h2:2'h2];
  assign T244 = T257 ? T251 : T245;
  assign T245 = T250 ? T248 : T246;
  assign T246 = T247 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T247 = T233[1'h0:1'h0];
  assign T248 = T249 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T249 = T233[1'h0:1'h0];
  assign T250 = T233[1'h1:1'h1];
  assign T251 = T256 ? T254 : T252;
  assign T252 = T253 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T253 = T233[1'h0:1'h0];
  assign T254 = T255 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T255 = T233[1'h0:1'h0];
  assign T256 = T233[1'h1:1'h1];
  assign T257 = T233[2'h2:2'h2];
  assign T258 = T233[2'h3:2'h3];
  assign T259 = T288 ? T274 : T260;
  assign T260 = T273 ? T267 : T261;
  assign T261 = T266 ? T264 : T262;
  assign T262 = T263 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T263 = T233[1'h0:1'h0];
  assign T264 = T265 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T265 = T233[1'h0:1'h0];
  assign T266 = T233[1'h1:1'h1];
  assign T267 = T272 ? T270 : T268;
  assign T268 = T269 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T269 = T233[1'h0:1'h0];
  assign T270 = T271 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T271 = T233[1'h0:1'h0];
  assign T272 = T233[1'h1:1'h1];
  assign T273 = T233[2'h2:2'h2];
  assign T274 = T287 ? T281 : T275;
  assign T275 = T280 ? T278 : T276;
  assign T276 = T277 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T277 = T233[1'h0:1'h0];
  assign T278 = T279 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T279 = T233[1'h0:1'h0];
  assign T280 = T233[1'h1:1'h1];
  assign T281 = T286 ? T284 : T282;
  assign T282 = T283 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T283 = T233[1'h0:1'h0];
  assign T284 = T285 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T285 = T233[1'h0:1'h0];
  assign T286 = T233[1'h1:1'h1];
  assign T287 = T233[2'h2:2'h2];
  assign T288 = T233[2'h3:2'h3];
  assign T289 = T233[3'h4:3'h4];
  assign T290 = T351 ? T321 : T291;
  assign T291 = T320 ? T306 : T292;
  assign T292 = T305 ? T299 : T293;
  assign T293 = T298 ? T296 : T294;
  assign T294 = T295 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T295 = T233[1'h0:1'h0];
  assign T296 = T297 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T297 = T233[1'h0:1'h0];
  assign T298 = T233[1'h1:1'h1];
  assign T299 = T304 ? T302 : T300;
  assign T300 = T301 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T301 = T233[1'h0:1'h0];
  assign T302 = T303 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T303 = T233[1'h0:1'h0];
  assign T304 = T233[1'h1:1'h1];
  assign T305 = T233[2'h2:2'h2];
  assign T306 = T319 ? T313 : T307;
  assign T307 = T312 ? T310 : T308;
  assign T308 = T309 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T309 = T233[1'h0:1'h0];
  assign T310 = T311 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T311 = T233[1'h0:1'h0];
  assign T312 = T233[1'h1:1'h1];
  assign T313 = T318 ? T316 : T314;
  assign T314 = T315 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T315 = T233[1'h0:1'h0];
  assign T316 = T317 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T317 = T233[1'h0:1'h0];
  assign T318 = T233[1'h1:1'h1];
  assign T319 = T233[2'h2:2'h2];
  assign T320 = T233[2'h3:2'h3];
  assign T321 = T350 ? T336 : T322;
  assign T322 = T335 ? T329 : T323;
  assign T323 = T328 ? T326 : T324;
  assign T324 = T325 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T325 = T233[1'h0:1'h0];
  assign T326 = T327 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T327 = T233[1'h0:1'h0];
  assign T328 = T233[1'h1:1'h1];
  assign T329 = T334 ? T332 : T330;
  assign T330 = T331 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T331 = T233[1'h0:1'h0];
  assign T332 = T333 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T333 = T233[1'h0:1'h0];
  assign T334 = T233[1'h1:1'h1];
  assign T335 = T233[2'h2:2'h2];
  assign T336 = T349 ? T343 : T337;
  assign T337 = T342 ? T340 : T338;
  assign T338 = T339 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T339 = T233[1'h0:1'h0];
  assign T340 = T341 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T341 = T233[1'h0:1'h0];
  assign T342 = T233[1'h1:1'h1];
  assign T343 = T348 ? T346 : T344;
  assign T344 = T345 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T345 = T233[1'h0:1'h0];
  assign T346 = T347 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T347 = T233[1'h0:1'h0];
  assign T348 = T233[1'h1:1'h1];
  assign T349 = T233[2'h2:2'h2];
  assign T350 = T233[2'h3:2'h3];
  assign T351 = T233[3'h4:3'h4];
  assign T352 = T233[3'h5:3'h5];
  assign T353 = T355 | T354;
  assign T354 = cmd == 4'h3;
  assign T355 = cmd == 4'h2;
  assign tx_header = {T357, T356};
  assign T356 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T357 = {addr, seqno};
  assign T358 = T20 ? T359 : seqno;
  assign T359 = rx_shifter_in[5'h17:5'h10];
  assign T360 = tx_word_count == 13'h0;
  assign io_host_out_valid = T361;
  assign T361 = state == 3'h7;
  assign io_host_in_ready = T362;
  assign T362 = state == 3'h0;

  always @(posedge clk) begin
    if (T2)
      packet_ram[T135] <= T1;
    if(reset) begin
      state <= 3'h0;
    end else if(T132) begin
      state <= 3'h7;
    end else if(T130) begin
      state <= 3'h7;
    end else if(T125) begin
      state <= 3'h7;
    end else if(T122) begin
      state <= 3'h2;
    end else if(T112) begin
      state <= T108;
    end else if(T106) begin
      state <= T102;
    end else if(T100) begin
      state <= T90;
    end else if(T88) begin
      state <= 3'h5;
    end else if(T78) begin
      state <= 3'h6;
    end else if(T65) begin
      state <= T14;
    end
    if(T20) begin
      cmd <= next_cmd;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T25) begin
      rx_count <= 15'h0;
    end else if(T60) begin
      rx_count <= T24;
    end
    if(T20) begin
      size <= T28;
    end
    if(T60) begin
      rx_shifter <= rx_shifter_in;
    end
    if(T106) begin
      addr <= T50;
    end else if(T100) begin
      addr <= T49;
    end else if(T20) begin
      addr <= T48;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T25) begin
      tx_count <= 15'h0;
    end else if(T59) begin
      tx_count <= T58;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T82) begin
      cnt <= T81;
    end
    if(T106) begin
      pos <= T98;
    end else if(T100) begin
      pos <= T97;
    end else if(T20) begin
      pos <= T96;
    end
    if (T138)
      packet_ram[T140] <= T137;
    if (T142)
      packet_ram[T143] <= rx_shifter_in;
    if(reset) begin
      R180 <= 1'h0;
    end else if(T183) begin
      R180 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R180 <= 1'h0;
    end
    if(reset) begin
      rtc <= 64'h0;
    end else if(rtc_tick) begin
      rtc <= T187;
    end
    if(reset) begin
      R188 <= 7'h0;
    end else if(rtc_tick) begin
      R188 <= 7'h0;
    end else begin
      R188 <= T190;
    end
    if(reset) begin
      R193 <= 1'h0;
    end else if(T191) begin
      R193 <= io_cpu_0_pcr_req_ready;
    end else if(io_cpu_0_pcr_rep_valid) begin
      R193 <= 1'h0;
    end
    if(reset) begin
      R198 <= 1'h0;
    end else if(T191) begin
      R198 <= io_cpu_0_pcr_req_ready;
    end else if(rtc_tick) begin
      R198 <= 1'h0;
    end
    if(reset) begin
      R213 <= 1'h1;
    end else if(T216) begin
      R213 <= T215;
    end
    if(T132) begin
      pcrReadData <= T226;
    end else if(T130) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T125) begin
      pcrReadData <= T379;
    end
    if(T20) begin
      seqno <= T359;
    end
  end
endmodule

module ClientTileLinkIOWrapper_0(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input  io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[127:0] io_in_grant_bits_data,
    output io_in_grant_bits_client_xact_id,
    output[2:0] io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output[127:0] io_out_acquire_bits_data,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [127:0] io_out_grant_bits_data,
    input  io_out_grant_bits_client_xact_id,
    input [2:0] io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[25:0] io_out_release_bits_addr_block
    //output io_out_release_bits_client_xact_id
    //output[1:0] io_out_release_bits_addr_beat
    //output[127:0] io_out_release_bits_data
    //output[2:0] io_out_release_bits_r_type
    //output io_out_release_bits_voluntary
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module FinishQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_fin_manager_xact_id,
    input [1:0] io_enq_bits_dst,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_fin_manager_xact_id,
    output[1:0] io_deq_bits_dst,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[4:0] T11;
  reg [4:0] ram [1:0];
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[2:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_dst = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_fin_manager_xact_id, io_enq_bits_dst};
  assign io_deq_bits_fin_manager_xact_id = T15;
  assign T15 = T11[3'h4:2'h2];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module FinishUnit_0(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [127:0] io_grant_bits_payload_data,
    input  io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[127:0] io_refill_bits_data,
    output io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h0;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue_0 FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input  io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[127:0] io_client_grant_bits_data,
    output io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [25:0] io_client_release_bits_addr_block,
    input  io_client_release_bits_client_xact_id,
    input [1:0] io_client_release_bits_addr_beat,
    input [127:0] io_client_release_bits_data,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[25:0] io_network_release_bits_payload_addr_block,
    output io_network_release_bits_payload_client_xact_id,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[127:0] io_network_release_bits_payload_data,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary
);

  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[127:0] rel_with_header_bits_payload_data;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h0;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h0;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_0 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input  io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [127:0] io_enq_bits_payload_data,
    input  io_enq_bits_payload_is_builtin_type,
    input [2:0] io_enq_bits_payload_a_type,
    input [16:0] io_enq_bits_payload_union,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[127:0] io_deq_bits_payload_data,
    output io_deq_bits_payload_is_builtin_type,
    output[2:0] io_deq_bits_payload_a_type,
    output[16:0] io_deq_bits_payload_union,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T33;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T34;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T35;
  wire T8;
  wire T9;
  wire[16:0] T10;
  wire[181:0] T11;
  reg [181:0] ram [1:0];
  wire[181:0] T12;
  wire[181:0] T13;
  wire[181:0] T14;
  wire[150:0] T15;
  wire[20:0] T16;
  wire[19:0] T17;
  wire[129:0] T18;
  wire[30:0] T19;
  wire[26:0] T20;
  wire[3:0] T21;
  wire[2:0] T22;
  wire T23;
  wire[127:0] T24;
  wire[1:0] T25;
  wire T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire empty;
  wire T31;
  wire T32;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T33 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T34 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T35 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_union = T10;
  assign T10 = T11[5'h10:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T19, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_payload_is_builtin_type, T17};
  assign T17 = {io_enq_bits_payload_a_type, io_enq_bits_payload_union};
  assign T18 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_data};
  assign T19 = {T21, T20};
  assign T20 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T21 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_a_type = T22;
  assign T22 = T11[5'h13:5'h11];
  assign io_deq_bits_payload_is_builtin_type = T23;
  assign T23 = T11[5'h14:5'h14];
  assign io_deq_bits_payload_data = T24;
  assign T24 = T11[8'h94:5'h15];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h96:8'h95];
  assign io_deq_bits_payload_client_xact_id = T26;
  assign T26 = T11[8'h97:8'h97];
  assign io_deq_bits_payload_addr_block = T27;
  assign T27 = T11[8'hb1:8'h98];
  assign io_deq_bits_header_dst = T28;
  assign T28 = T11[8'hb3:8'hb2];
  assign io_deq_bits_header_src = T29;
  assign T29 = T11[8'hb5:8'hb4];
  assign io_deq_valid = T30;
  assign T30 = empty ^ 1'h1;
  assign empty = ptr_match & T31;
  assign T31 = maybe_full ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_p_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T23;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T24;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[27:0] T15;
  wire[3:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_p_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_p_type};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T11[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T11[5'h1d:5'h1c];
  assign io_deq_bits_header_src = T19;
  assign T19 = T11[5'h1f:5'h1e];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input  io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [127:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_enq_bits_payload_voluntary,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[127:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type,
    output io_deq_bits_payload_voluntary,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire T10;
  wire[164:0] T11;
  reg [164:0] ram [1:0];
  wire[164:0] T12;
  wire[164:0] T13;
  wire[164:0] T14;
  wire[133:0] T15;
  wire[3:0] T16;
  wire[129:0] T17;
  wire[30:0] T18;
  wire[26:0] T19;
  wire[3:0] T20;
  wire[2:0] T21;
  wire[127:0] T22;
  wire[1:0] T23;
  wire T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_voluntary = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_r_type, io_enq_bits_payload_voluntary};
  assign T17 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_data};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T21;
  assign T21 = T11[2'h3:1'h1];
  assign io_deq_bits_payload_data = T22;
  assign T22 = T11[8'h83:3'h4];
  assign io_deq_bits_payload_addr_beat = T23;
  assign T23 = T11[8'h85:8'h84];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[8'h86:8'h86];
  assign io_deq_bits_payload_addr_block = T25;
  assign T25 = T11[8'ha0:8'h87];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'ha2:8'ha1];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'ha4:8'ha3];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [127:0] io_enq_bits_payload_data,
    input  io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_manager_xact_id,
    input  io_enq_bits_payload_is_builtin_type,
    input [3:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[127:0] io_deq_bits_payload_data,
    output io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_manager_xact_id,
    output io_deq_bits_payload_is_builtin_type,
    output[3:0] io_deq_bits_payload_g_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire[142:0] T11;
  reg [142:0] ram [1:0];
  wire[142:0] T12;
  wire[142:0] T13;
  wire[142:0] T14;
  wire[8:0] T15;
  wire[4:0] T16;
  wire[3:0] T17;
  wire[133:0] T18;
  wire[129:0] T19;
  wire[3:0] T20;
  wire T21;
  wire[2:0] T22;
  wire T23;
  wire[127:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_g_type = T10;
  assign T10 = T11[2'h3:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_is_builtin_type, io_enq_bits_payload_g_type};
  assign T17 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_manager_xact_id};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_data};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_is_builtin_type = T21;
  assign T21 = T11[3'h4:3'h4];
  assign io_deq_bits_payload_manager_xact_id = T22;
  assign T22 = T11[3'h7:3'h5];
  assign io_deq_bits_payload_client_xact_id = T23;
  assign T23 = T11[4'h8:4'h8];
  assign io_deq_bits_payload_data = T24;
  assign T24 = T11[8'h88:4'h9];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h8a:8'h89];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'h8c:8'h8b];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'h8e:8'h8d];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_manager_xact_id,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[6:0] T11;
  reg [6:0] ram [1:0];
  wire[6:0] T12;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[4:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_manager_xact_id = T10;
  assign T10 = T11[2'h2:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_header_src, T15};
  assign T15 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T16;
  assign T16 = T11[3'h4:2'h3];
  assign io_deq_bits_header_src = T17;
  assign T17 = T11[3'h6:3'h5];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module TileLinkEnqueuer_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input  io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_grant_bits_payload_client_xact_id,
    output[2:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [2:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [25:0] io_client_release_bits_payload_addr_block,
    input  io_client_release_bits_payload_client_xact_id,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [127:0] io_client_release_bits_payload_data,
    input [2:0] io_client_release_bits_payload_r_type,
    input  io_client_release_bits_payload_voluntary,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_grant_bits_payload_client_xact_id,
    input [2:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[2:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output io_manager_release_bits_payload_client_xact_id,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[127:0] io_manager_release_bits_payload_data,
    output[2:0] io_manager_release_bits_payload_r_type,
    output io_manager_release_bits_payload_voluntary
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire Queue_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire[127:0] Queue_io_deq_bits_payload_data;
  wire Queue_io_deq_bits_payload_is_builtin_type;
  wire[2:0] Queue_io_deq_bits_payload_a_type;
  wire[16:0] Queue_io_deq_bits_payload_union;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[1:0] Queue_1_io_deq_bits_header_src;
  wire[1:0] Queue_1_io_deq_bits_header_dst;
  wire[25:0] Queue_1_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_1_io_deq_bits_payload_p_type;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[1:0] Queue_2_io_deq_bits_header_src;
  wire[1:0] Queue_2_io_deq_bits_header_dst;
  wire[25:0] Queue_2_io_deq_bits_payload_addr_block;
  wire Queue_2_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_2_io_deq_bits_payload_addr_beat;
  wire[127:0] Queue_2_io_deq_bits_payload_data;
  wire[2:0] Queue_2_io_deq_bits_payload_r_type;
  wire Queue_2_io_deq_bits_payload_voluntary;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_header_src;
  wire[1:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_payload_addr_beat;
  wire[127:0] Queue_3_io_deq_bits_payload_data;
  wire Queue_3_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_3_io_deq_bits_payload_manager_xact_id;
  wire Queue_3_io_deq_bits_payload_is_builtin_type;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[2:0] Queue_4_io_deq_bits_payload_manager_xact_id;


  assign io_manager_release_bits_payload_voluntary = Queue_2_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_2_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_2_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_2_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_header_dst = Queue_2_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_2_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_2_io_deq_valid;
  assign io_manager_probe_ready = Queue_1_io_enq_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = Queue_4_io_deq_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_finish_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_finish_valid = Queue_4_io_deq_valid;
  assign io_manager_grant_ready = Queue_3_io_enq_ready;
  assign io_manager_acquire_bits_payload_union = Queue_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = Queue_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_acquire_valid = Queue_io_deq_valid;
  assign io_client_release_ready = Queue_2_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = Queue_1_io_deq_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = Queue_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = Queue_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_header_src = Queue_1_io_deq_bits_header_src;
  assign io_client_probe_valid = Queue_1_io_deq_valid;
  assign io_client_finish_ready = Queue_4_io_enq_ready;
  assign io_client_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_client_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_client_grant_valid = Queue_3_io_deq_valid;
  assign io_client_acquire_ready = Queue_io_enq_ready;
  Queue_5 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_acquire_valid ),
       .io_enq_bits_header_src( io_client_acquire_bits_header_src ),
       .io_enq_bits_header_dst( io_client_acquire_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_acquire_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_acquire_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_acquire_bits_payload_addr_beat ),
       .io_enq_bits_payload_data( io_client_acquire_bits_payload_data ),
       .io_enq_bits_payload_is_builtin_type( io_client_acquire_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_a_type( io_client_acquire_bits_payload_a_type ),
       .io_enq_bits_payload_union( io_client_acquire_bits_payload_union ),
       .io_deq_ready( io_manager_acquire_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data ),
       .io_deq_bits_payload_is_builtin_type( Queue_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_a_type( Queue_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_union( Queue_io_deq_bits_payload_union )
       //.io_count(  )
  );
  Queue_6 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( io_manager_probe_valid ),
       .io_enq_bits_header_src( io_manager_probe_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_probe_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_manager_probe_bits_payload_addr_block ),
       .io_enq_bits_payload_p_type( io_manager_probe_bits_payload_p_type ),
       .io_deq_ready( io_client_probe_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_1_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_p_type( Queue_1_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
  Queue_7 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_2_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_2_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_2_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_data( Queue_2_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_2_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_voluntary( Queue_2_io_deq_bits_payload_voluntary )
       //.io_count(  )
  );
  Queue_8 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( io_manager_grant_valid ),
       .io_enq_bits_header_src( io_manager_grant_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_grant_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_manager_grant_bits_payload_addr_beat ),
       .io_enq_bits_payload_data( io_manager_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( io_manager_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( io_manager_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_is_builtin_type( io_manager_grant_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_g_type( io_manager_grant_bits_payload_g_type ),
       .io_deq_ready( io_client_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_3_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_3_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_is_builtin_type( Queue_3_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type )
       //.io_count(  )
  );
  Queue_9 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( io_client_finish_valid ),
       .io_enq_bits_header_src( io_client_finish_bits_header_src ),
       .io_enq_bits_header_dst( io_client_finish_bits_header_dst ),
       .io_enq_bits_payload_manager_xact_id( io_client_finish_bits_payload_manager_xact_id ),
       .io_deq_ready( io_manager_finish_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_4_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
endmodule

module FinishUnit_1(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [127:0] io_grant_bits_payload_data,
    input  io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[127:0] io_refill_bits_data,
    output io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue_0 FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input  io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[127:0] io_client_grant_bits_data,
    output io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [25:0] io_client_release_bits_addr_block,
    input  io_client_release_bits_client_xact_id,
    input [1:0] io_client_release_bits_addr_beat,
    input [127:0] io_client_release_bits_data,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[25:0] io_network_release_bits_payload_addr_block,
    output io_network_release_bits_payload_client_xact_id,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[127:0] io_network_release_bits_payload_data,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary
);

  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[127:0] rel_with_header_bits_payload_data;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h1;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h1;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_1 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module FinishUnit_2(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [127:0] io_grant_bits_payload_data,
    input  io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[127:0] io_refill_bits_data,
    output io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T33;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T33 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h2;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T27;
  assign T27 = T28 & io_refill_ready;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue_0 FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_2(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input  io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[127:0] io_client_grant_bits_data,
    output io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [25:0] io_client_release_bits_addr_block,
    input  io_client_release_bits_client_xact_id,
    input [1:0] io_client_release_bits_addr_beat,
    input [127:0] io_client_release_bits_data,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[25:0] io_network_release_bits_payload_addr_block,
    output io_network_release_bits_payload_client_xact_id,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[127:0] io_network_release_bits_payload_data,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary
);

  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[127:0] rel_with_header_bits_payload_data;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h2;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h2;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_2 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module ManagerTileLinkNetworkPort_0(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output[127:0] io_manager_acquire_bits_data,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output[1:0] io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [127:0] io_manager_grant_bits_data,
    input  io_manager_grant_bits_client_xact_id,
    input [2:0] io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input [1:0] io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[2:0] io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input [1:0] io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[25:0] io_manager_release_bits_addr_block,
    output io_manager_release_bits_client_xact_id,
    output[1:0] io_manager_release_bits_addr_beat,
    output[127:0] io_manager_release_bits_data,
    output[2:0] io_manager_release_bits_r_type,
    output io_manager_release_bits_voluntary,
    output[1:0] io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input [1:0] io_network_acquire_bits_header_src,
    input [1:0] io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input  io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output[1:0] io_network_grant_bits_header_src,
    output[1:0] io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[127:0] io_network_grant_bits_payload_data,
    output io_network_grant_bits_payload_client_xact_id,
    output[2:0] io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input [1:0] io_network_finish_bits_header_src,
    input [1:0] io_network_finish_bits_header_dst,
    input [2:0] io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output[1:0] io_network_probe_bits_header_src,
    output[1:0] io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input [1:0] io_network_release_bits_header_src,
    input [1:0] io_network_release_bits_header_dst,
    input [25:0] io_network_release_bits_payload_addr_block,
    input  io_network_release_bits_payload_client_xact_id,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [127:0] io_network_release_bits_payload_data,
    input [2:0] io_network_release_bits_payload_r_type,
    input  io_network_release_bits_payload_voluntary
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire[3:0] T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire[127:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[127:0] T19;
  wire[1:0] T20;
  wire T21;
  wire[25:0] T22;
  wire T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire[16:0] T28;
  wire[2:0] T29;
  wire T30;
  wire[127:0] T31;
  wire[1:0] T32;
  wire T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = io_manager_probe_bits_client_id;
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 2'h0;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_g_type = T7;
  assign T7 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T8;
  assign T8 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T9;
  assign T9 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T10;
  assign T10 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_data = T11;
  assign T11 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = io_manager_grant_bits_client_id;
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 2'h0;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src;
  assign io_manager_release_bits_voluntary = T17;
  assign T17 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_r_type = T18;
  assign T18 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_data = T19;
  assign T19 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_addr_beat = T20;
  assign T20 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_bits_client_xact_id = T21;
  assign T21 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T22;
  assign T22 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src;
  assign io_manager_acquire_bits_union = T28;
  assign T28 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T29;
  assign T29 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T30;
  assign T30 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_data = T31;
  assign T31 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input  io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [127:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_enq_bits_payload_voluntary,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[127:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type,
    output io_deq_bits_payload_voluntary,
    output io_count
);

  wire T23;
  wire[1:0] T0;
  reg  full;
  wire T24;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire T3;
  wire[164:0] T4;
  reg [164:0] ram [0:0];
  wire[164:0] T5;
  wire[164:0] T6;
  wire[164:0] T7;
  wire[133:0] T8;
  wire[3:0] T9;
  wire[129:0] T10;
  wire[30:0] T11;
  wire[26:0] T12;
  wire[3:0] T13;
  wire[2:0] T14;
  wire[127:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[25:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire empty;
  wire T22;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T23;
  assign T23 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T24 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_voluntary = T3;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_payload_r_type, io_enq_bits_payload_voluntary};
  assign T10 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_data};
  assign T11 = {T13, T12};
  assign T12 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T13 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T14;
  assign T14 = T4[2'h3:1'h1];
  assign io_deq_bits_payload_data = T15;
  assign T15 = T4[8'h83:3'h4];
  assign io_deq_bits_payload_addr_beat = T16;
  assign T16 = T4[8'h85:8'h84];
  assign io_deq_bits_payload_client_xact_id = T17;
  assign T17 = T4[8'h86:8'h86];
  assign io_deq_bits_payload_addr_block = T18;
  assign T18 = T4[8'ha0:8'h87];
  assign io_deq_bits_header_dst = T19;
  assign T19 = T4[8'ha2:8'ha1];
  assign io_deq_bits_header_src = T20;
  assign T20 = T4[8'ha4:8'ha3];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module TileLinkEnqueuer_2(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input  io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_grant_bits_payload_client_xact_id,
    output[2:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [2:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [25:0] io_client_release_bits_payload_addr_block,
    input  io_client_release_bits_payload_client_xact_id,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [127:0] io_client_release_bits_payload_data,
    input [2:0] io_client_release_bits_payload_r_type,
    input  io_client_release_bits_payload_voluntary,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_grant_bits_payload_client_xact_id,
    input [2:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[2:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output io_manager_release_bits_payload_client_xact_id,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[127:0] io_manager_release_bits_payload_data,
    output[2:0] io_manager_release_bits_payload_r_type,
    output io_manager_release_bits_payload_voluntary
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire Queue_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire[127:0] Queue_io_deq_bits_payload_data;
  wire[2:0] Queue_io_deq_bits_payload_r_type;
  wire Queue_io_deq_bits_payload_voluntary;


  assign io_manager_release_bits_payload_voluntary = Queue_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_io_deq_valid;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_client_release_ready = Queue_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_acquire_ready = io_manager_acquire_ready;
  Queue_10 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_voluntary( Queue_io_deq_bits_payload_voluntary )
       //.io_count(  )
  );
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input  io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [127:0] io_in_2_bits_payload_data,
    input  io_in_2_bits_payload_is_builtin_type,
    input [2:0] io_in_2_bits_payload_a_type,
    input [16:0] io_in_2_bits_payload_union,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input  io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [127:0] io_in_1_bits_payload_data,
    input  io_in_1_bits_payload_is_builtin_type,
    input [2:0] io_in_1_bits_payload_a_type,
    input [16:0] io_in_1_bits_payload_union,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input  io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [127:0] io_in_0_bits_payload_data,
    input  io_in_0_bits_payload_is_builtin_type,
    input [2:0] io_in_0_bits_payload_a_type,
    input [16:0] io_in_0_bits_payload_union,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output io_out_bits_payload_client_xact_id,
    output[1:0] io_out_bits_payload_addr_beat,
    output[127:0] io_out_bits_payload_data,
    output io_out_bits_payload_is_builtin_type,
    output[2:0] io_out_bits_payload_a_type,
    output[16:0] io_out_bits_payload_union,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T107;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T108;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  locked;
  wire T109;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  reg [1:0] R26;
  wire[1:0] T110;
  wire[1:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire T30;
  wire[1:0] T31;
  wire T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[127:0] T41;
  wire[127:0] T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[25:0] T53;
  wire[25:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R26 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T107 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T108 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T20 & T18;
  assign T18 = io_out_bits_payload_is_builtin_type & T19;
  assign T19 = 3'h3 == io_out_bits_payload_a_type;
  assign T20 = io_out_ready & io_out_valid;
  assign T109 = reset ? 1'h0 : T21;
  assign T21 = T23 ? 1'h0 : T22;
  assign T22 = T15 ? 1'h1 : locked;
  assign T23 = T20 & T24;
  assign T24 = T25 == 2'h0;
  assign T25 = R26 + 2'h1;
  assign T110 = reset ? 2'h0 : T27;
  assign T27 = T17 ? T25 : R26;
  assign io_out_bits_payload_union = T28;
  assign T28 = T32 ? io_in_2_bits_payload_union : T29;
  assign T29 = T30 ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign T30 = T31[1'h0:1'h0];
  assign T31 = chosen;
  assign T32 = T31[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T33;
  assign T33 = T36 ? io_in_2_bits_payload_a_type : T34;
  assign T34 = T35 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T35 = T31[1'h0:1'h0];
  assign T36 = T31[1'h1:1'h1];
  assign io_out_bits_payload_is_builtin_type = T37;
  assign T37 = T40 ? io_in_2_bits_payload_is_builtin_type : T38;
  assign T38 = T39 ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign T39 = T31[1'h0:1'h0];
  assign T40 = T31[1'h1:1'h1];
  assign io_out_bits_payload_data = T41;
  assign T41 = T44 ? io_in_2_bits_payload_data : T42;
  assign T42 = T43 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T43 = T31[1'h0:1'h0];
  assign T44 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T45;
  assign T45 = T48 ? io_in_2_bits_payload_addr_beat : T46;
  assign T46 = T47 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T47 = T31[1'h0:1'h0];
  assign T48 = T31[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T49;
  assign T49 = T52 ? io_in_2_bits_payload_client_xact_id : T50;
  assign T50 = T51 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T51 = T31[1'h0:1'h0];
  assign T52 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T53;
  assign T53 = T56 ? io_in_2_bits_payload_addr_block : T54;
  assign T54 = T55 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T55 = T31[1'h0:1'h0];
  assign T56 = T31[1'h1:1'h1];
  assign io_out_bits_header_dst = T57;
  assign T57 = T60 ? io_in_2_bits_header_dst : T58;
  assign T58 = T59 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T59 = T31[1'h0:1'h0];
  assign T60 = T31[1'h1:1'h1];
  assign io_out_bits_header_src = T61;
  assign T61 = T64 ? io_in_2_bits_header_src : T62;
  assign T62 = T63 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T63 = T31[1'h0:1'h0];
  assign T64 = T31[1'h1:1'h1];
  assign io_out_valid = T65;
  assign T65 = T68 ? io_in_2_valid : T66;
  assign T66 = T67 ? io_in_1_valid : io_in_0_valid;
  assign T67 = T31[1'h0:1'h0];
  assign T68 = T31[1'h1:1'h1];
  assign io_in_0_ready = T69;
  assign T69 = T70 & io_out_ready;
  assign T70 = locked ? T82 : T71;
  assign T71 = T81 | T72;
  assign T72 = T73 ^ 1'h1;
  assign T73 = T76 | T74;
  assign T74 = io_in_2_valid & T75;
  assign T75 = last_grant < 2'h2;
  assign T76 = T79 | T77;
  assign T77 = io_in_1_valid & T78;
  assign T78 = last_grant < 2'h1;
  assign T79 = io_in_0_valid & T80;
  assign T80 = last_grant < 2'h0;
  assign T81 = last_grant < 2'h0;
  assign T82 = lockIdx == 2'h0;
  assign io_in_1_ready = T83;
  assign T83 = T84 & io_out_ready;
  assign T84 = locked ? T93 : T85;
  assign T85 = T90 | T86;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | io_in_0_valid;
  assign T88 = T89 | T74;
  assign T89 = T79 | T77;
  assign T90 = T92 & T91;
  assign T91 = last_grant < 2'h1;
  assign T92 = T79 ^ 1'h1;
  assign T93 = lockIdx == 2'h1;
  assign io_in_2_ready = T94;
  assign T94 = T95 & io_out_ready;
  assign T95 = locked ? T106 : T96;
  assign T96 = T102 | T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T99 | io_in_1_valid;
  assign T99 = T100 | io_in_0_valid;
  assign T100 = T101 | T74;
  assign T101 = T79 | T77;
  assign T102 = T104 & T103;
  assign T103 = last_grant < 2'h2;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T79 | T77;
  assign T106 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T23) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R26 <= 2'h0;
    end else if(T17) begin
      R26 <= T25;
    end
  end
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input  io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [127:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    input  io_in_2_bits_payload_voluntary,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input  io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [127:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    input  io_in_1_bits_payload_voluntary,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input  io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [127:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_in_0_bits_payload_voluntary,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output io_out_bits_payload_client_xact_id,
    output[1:0] io_out_bits_payload_addr_beat,
    output[127:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output io_out_bits_payload_voluntary,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T106;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T107;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg  locked;
  wire T108;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T109;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire[127:0] T40;
  wire[127:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[25:0] T52;
  wire[25:0] T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R29 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T106 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T107 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T23 & T18;
  assign T18 = T20 | T19;
  assign T19 = 3'h2 == io_out_bits_payload_r_type;
  assign T20 = T22 | T21;
  assign T21 = 3'h1 == io_out_bits_payload_r_type;
  assign T22 = 3'h0 == io_out_bits_payload_r_type;
  assign T23 = io_out_ready & io_out_valid;
  assign T108 = reset ? 1'h0 : T24;
  assign T24 = T26 ? 1'h0 : T25;
  assign T25 = T15 ? 1'h1 : locked;
  assign T26 = T23 & T27;
  assign T27 = T28 == 2'h0;
  assign T28 = R29 + 2'h1;
  assign T109 = reset ? 2'h0 : T30;
  assign T30 = T17 ? T28 : R29;
  assign io_out_bits_payload_voluntary = T31;
  assign T31 = T35 ? io_in_2_bits_payload_voluntary : T32;
  assign T32 = T33 ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign T33 = T34[1'h0:1'h0];
  assign T34 = chosen;
  assign T35 = T34[1'h1:1'h1];
  assign io_out_bits_payload_r_type = T36;
  assign T36 = T39 ? io_in_2_bits_payload_r_type : T37;
  assign T37 = T38 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T38 = T34[1'h0:1'h0];
  assign T39 = T34[1'h1:1'h1];
  assign io_out_bits_payload_data = T40;
  assign T40 = T43 ? io_in_2_bits_payload_data : T41;
  assign T41 = T42 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T42 = T34[1'h0:1'h0];
  assign T43 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T44;
  assign T44 = T47 ? io_in_2_bits_payload_addr_beat : T45;
  assign T45 = T46 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T46 = T34[1'h0:1'h0];
  assign T47 = T34[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T48;
  assign T48 = T51 ? io_in_2_bits_payload_client_xact_id : T49;
  assign T49 = T50 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T50 = T34[1'h0:1'h0];
  assign T51 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T52;
  assign T52 = T55 ? io_in_2_bits_payload_addr_block : T53;
  assign T53 = T54 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T54 = T34[1'h0:1'h0];
  assign T55 = T34[1'h1:1'h1];
  assign io_out_bits_header_dst = T56;
  assign T56 = T59 ? io_in_2_bits_header_dst : T57;
  assign T57 = T58 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T58 = T34[1'h0:1'h0];
  assign T59 = T34[1'h1:1'h1];
  assign io_out_bits_header_src = T60;
  assign T60 = T63 ? io_in_2_bits_header_src : T61;
  assign T61 = T62 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T62 = T34[1'h0:1'h0];
  assign T63 = T34[1'h1:1'h1];
  assign io_out_valid = T64;
  assign T64 = T67 ? io_in_2_valid : T65;
  assign T65 = T66 ? io_in_1_valid : io_in_0_valid;
  assign T66 = T34[1'h0:1'h0];
  assign T67 = T34[1'h1:1'h1];
  assign io_in_0_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = locked ? T81 : T70;
  assign T70 = T80 | T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T75 | T73;
  assign T73 = io_in_2_valid & T74;
  assign T74 = last_grant < 2'h2;
  assign T75 = T78 | T76;
  assign T76 = io_in_1_valid & T77;
  assign T77 = last_grant < 2'h1;
  assign T78 = io_in_0_valid & T79;
  assign T79 = last_grant < 2'h0;
  assign T80 = last_grant < 2'h0;
  assign T81 = lockIdx == 2'h0;
  assign io_in_1_ready = T82;
  assign T82 = T83 & io_out_ready;
  assign T83 = locked ? T92 : T84;
  assign T84 = T89 | T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T87 | io_in_0_valid;
  assign T87 = T88 | T73;
  assign T88 = T78 | T76;
  assign T89 = T91 & T90;
  assign T90 = last_grant < 2'h1;
  assign T91 = T78 ^ 1'h1;
  assign T92 = lockIdx == 2'h1;
  assign io_in_2_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = locked ? T105 : T95;
  assign T95 = T101 | T96;
  assign T96 = T97 ^ 1'h1;
  assign T97 = T98 | io_in_1_valid;
  assign T98 = T99 | io_in_0_valid;
  assign T99 = T100 | T73;
  assign T100 = T78 | T76;
  assign T101 = T103 & T102;
  assign T102 = last_grant < 2'h2;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T78 | T76;
  assign T105 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T26) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R29 <= 2'h0;
    end else if(T17) begin
      R29 <= T28;
    end
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_manager_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_payload_manager_xact_id = T9;
  assign T9 = T13 ? io_in_2_bits_payload_manager_xact_id : T10;
  assign T10 = T11 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_header_dst = T14;
  assign T14 = T17 ? io_in_2_bits_header_dst : T15;
  assign T15 = T16 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_header_src = T18;
  assign T18 = T21 ? io_in_2_bits_header_src : T19;
  assign T19 = T20 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module RocketChipTileLinkArbiter_0(input clk, input reset,
    output io_clients_2_acquire_ready,
    input  io_clients_2_acquire_valid,
    input [25:0] io_clients_2_acquire_bits_addr_block,
    input  io_clients_2_acquire_bits_client_xact_id,
    input [1:0] io_clients_2_acquire_bits_addr_beat,
    input [127:0] io_clients_2_acquire_bits_data,
    input  io_clients_2_acquire_bits_is_builtin_type,
    input [2:0] io_clients_2_acquire_bits_a_type,
    input [16:0] io_clients_2_acquire_bits_union,
    input  io_clients_2_grant_ready,
    output io_clients_2_grant_valid,
    output[1:0] io_clients_2_grant_bits_addr_beat,
    output[127:0] io_clients_2_grant_bits_data,
    output io_clients_2_grant_bits_client_xact_id,
    output[2:0] io_clients_2_grant_bits_manager_xact_id,
    output io_clients_2_grant_bits_is_builtin_type,
    output[3:0] io_clients_2_grant_bits_g_type,
    input  io_clients_2_probe_ready,
    output io_clients_2_probe_valid,
    output[25:0] io_clients_2_probe_bits_addr_block,
    output[1:0] io_clients_2_probe_bits_p_type,
    output io_clients_2_release_ready,
    input  io_clients_2_release_valid,
    input [25:0] io_clients_2_release_bits_addr_block,
    input  io_clients_2_release_bits_client_xact_id,
    input [1:0] io_clients_2_release_bits_addr_beat,
    input [127:0] io_clients_2_release_bits_data,
    input [2:0] io_clients_2_release_bits_r_type,
    input  io_clients_2_release_bits_voluntary,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [25:0] io_clients_1_acquire_bits_addr_block,
    input  io_clients_1_acquire_bits_client_xact_id,
    input [1:0] io_clients_1_acquire_bits_addr_beat,
    input [127:0] io_clients_1_acquire_bits_data,
    input  io_clients_1_acquire_bits_is_builtin_type,
    input [2:0] io_clients_1_acquire_bits_a_type,
    input [16:0] io_clients_1_acquire_bits_union,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_addr_beat,
    output[127:0] io_clients_1_grant_bits_data,
    output io_clients_1_grant_bits_client_xact_id,
    output[2:0] io_clients_1_grant_bits_manager_xact_id,
    output io_clients_1_grant_bits_is_builtin_type,
    output[3:0] io_clients_1_grant_bits_g_type,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[25:0] io_clients_1_probe_bits_addr_block,
    output[1:0] io_clients_1_probe_bits_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [25:0] io_clients_1_release_bits_addr_block,
    input  io_clients_1_release_bits_client_xact_id,
    input [1:0] io_clients_1_release_bits_addr_beat,
    input [127:0] io_clients_1_release_bits_data,
    input [2:0] io_clients_1_release_bits_r_type,
    input  io_clients_1_release_bits_voluntary,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [25:0] io_clients_0_acquire_bits_addr_block,
    input  io_clients_0_acquire_bits_client_xact_id,
    input [1:0] io_clients_0_acquire_bits_addr_beat,
    input [127:0] io_clients_0_acquire_bits_data,
    input  io_clients_0_acquire_bits_is_builtin_type,
    input [2:0] io_clients_0_acquire_bits_a_type,
    input [16:0] io_clients_0_acquire_bits_union,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_addr_beat,
    output[127:0] io_clients_0_grant_bits_data,
    output io_clients_0_grant_bits_client_xact_id,
    output[2:0] io_clients_0_grant_bits_manager_xact_id,
    output io_clients_0_grant_bits_is_builtin_type,
    output[3:0] io_clients_0_grant_bits_g_type,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[25:0] io_clients_0_probe_bits_addr_block,
    output[1:0] io_clients_0_probe_bits_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [25:0] io_clients_0_release_bits_addr_block,
    input  io_clients_0_release_bits_client_xact_id,
    input [1:0] io_clients_0_release_bits_addr_beat,
    input [127:0] io_clients_0_release_bits_data,
    input [2:0] io_clients_0_release_bits_r_type,
    input  io_clients_0_release_bits_voluntary,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[25:0] io_managers_0_acquire_bits_addr_block,
    output io_managers_0_acquire_bits_client_xact_id,
    output[1:0] io_managers_0_acquire_bits_addr_beat,
    output[127:0] io_managers_0_acquire_bits_data,
    output io_managers_0_acquire_bits_is_builtin_type,
    output[2:0] io_managers_0_acquire_bits_a_type,
    output[16:0] io_managers_0_acquire_bits_union,
    output[1:0] io_managers_0_acquire_bits_client_id,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_addr_beat,
    input [127:0] io_managers_0_grant_bits_data,
    input  io_managers_0_grant_bits_client_xact_id,
    input [2:0] io_managers_0_grant_bits_manager_xact_id,
    input  io_managers_0_grant_bits_is_builtin_type,
    input [3:0] io_managers_0_grant_bits_g_type,
    input [1:0] io_managers_0_grant_bits_client_id,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output[2:0] io_managers_0_finish_bits_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [25:0] io_managers_0_probe_bits_addr_block,
    input [1:0] io_managers_0_probe_bits_p_type,
    input [1:0] io_managers_0_probe_bits_client_id,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[25:0] io_managers_0_release_bits_addr_block,
    output io_managers_0_release_bits_client_xact_id,
    output[1:0] io_managers_0_release_bits_addr_beat,
    output[127:0] io_managers_0_release_bits_data,
    output[2:0] io_managers_0_release_bits_r_type,
    output io_managers_0_release_bits_voluntary,
    output[1:0] io_managers_0_release_bits_client_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_io_manager_finish_valid;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_io_manager_release_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_io_network_grant_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type;
  wire ManagerTileLinkNetworkPort_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_io_network_probe_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_io_network_release_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[1:0] LockingRRArbiter_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_payload_union;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire LockingRRArbiter_1_io_out_bits_payload_voluntary;
  wire RRArbiter_io_in_2_ready;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[1:0] RRArbiter_io_out_bits_header_src;
  wire[1:0] RRArbiter_io_out_bits_header_dst;
  wire[2:0] RRArbiter_io_out_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_acquire_ready;
  wire TileLinkEnqueuer_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_io_client_finish_ready;
  wire TileLinkEnqueuer_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_io_client_release_ready;
  wire TileLinkEnqueuer_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_io_manager_grant_ready;
  wire TileLinkEnqueuer_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_manager_probe_ready;
  wire TileLinkEnqueuer_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  wire TileLinkEnqueuer_1_io_client_acquire_ready;
  wire TileLinkEnqueuer_1_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_1_io_client_finish_ready;
  wire TileLinkEnqueuer_1_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_1_io_client_release_ready;
  wire TileLinkEnqueuer_1_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_1_io_manager_grant_ready;
  wire TileLinkEnqueuer_1_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_manager_probe_ready;
  wire TileLinkEnqueuer_1_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  wire TileLinkEnqueuer_2_io_client_acquire_ready;
  wire TileLinkEnqueuer_2_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_2_io_client_finish_ready;
  wire TileLinkEnqueuer_2_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_2_io_client_release_ready;
  wire TileLinkEnqueuer_2_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block;
  wire TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_2_io_manager_grant_ready;
  wire TileLinkEnqueuer_2_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_manager_probe_ready;
  wire TileLinkEnqueuer_2_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block;
  wire TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary;
  wire TileLinkEnqueuer_3_io_client_acquire_ready;
  wire TileLinkEnqueuer_3_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_3_io_client_finish_ready;
  wire TileLinkEnqueuer_3_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_3_io_client_release_ready;
  wire TileLinkEnqueuer_3_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block;
  wire TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_3_io_manager_grant_ready;
  wire TileLinkEnqueuer_3_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_manager_probe_ready;
  wire TileLinkEnqueuer_3_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block;
  wire TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary;
  wire ClientTileLinkNetworkPort_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  wire ClientTileLinkNetworkPort_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_io_client_release_ready;
  wire ClientTileLinkNetworkPort_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union;
  wire ClientTileLinkNetworkPort_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_data;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary;
  wire ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_2_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  wire ClientTileLinkNetworkPort_2_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_2_io_client_release_ready;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire ClientTileLinkNetworkPort_2_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_2_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_2_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;


  assign T0 = T5 ? TileLinkEnqueuer_2_io_manager_probe_ready : T1;
  assign T1 = T4 ? TileLinkEnqueuer_1_io_manager_probe_ready : T2;
  assign T2 = T3 ? TileLinkEnqueuer_io_manager_probe_ready : 1'h0;
  assign T3 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h0;
  assign T4 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h1;
  assign T5 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h2;
  assign T6 = T11 ? TileLinkEnqueuer_2_io_manager_grant_ready : T7;
  assign T7 = T10 ? TileLinkEnqueuer_1_io_manager_grant_ready : T8;
  assign T8 = T9 ? TileLinkEnqueuer_io_manager_grant_ready : 1'h0;
  assign T9 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h0;
  assign T10 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h1;
  assign T11 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h2;
  assign T12 = T5 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T13 = T11 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T14 = T4 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T15 = T10 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T16 = T3 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T17 = T9 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_io_manager_release_valid;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_io_manager_probe_ready;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_io_manager_finish_valid;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_io_manager_grant_ready;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  assign io_clients_0_release_ready = ClientTileLinkNetworkPort_io_client_release_ready;
  assign io_clients_0_probe_bits_p_type = ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  assign io_clients_0_probe_bits_addr_block = ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  assign io_clients_0_probe_valid = ClientTileLinkNetworkPort_io_client_probe_valid;
  assign io_clients_0_grant_bits_g_type = ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  assign io_clients_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  assign io_clients_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  assign io_clients_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  assign io_clients_0_grant_bits_data = ClientTileLinkNetworkPort_io_client_grant_bits_data;
  assign io_clients_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  assign io_clients_0_grant_valid = ClientTileLinkNetworkPort_io_client_grant_valid;
  assign io_clients_0_acquire_ready = ClientTileLinkNetworkPort_io_client_acquire_ready;
  assign io_clients_1_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_1_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_1_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_1_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_1_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_1_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_1_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_1_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_1_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_1_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_1_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_1_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_2_release_ready = ClientTileLinkNetworkPort_2_io_client_release_ready;
  assign io_clients_2_probe_bits_p_type = ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  assign io_clients_2_probe_bits_addr_block = ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  assign io_clients_2_probe_valid = ClientTileLinkNetworkPort_2_io_client_probe_valid;
  assign io_clients_2_grant_bits_g_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  assign io_clients_2_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  assign io_clients_2_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  assign io_clients_2_grant_bits_client_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  assign io_clients_2_grant_bits_data = ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  assign io_clients_2_grant_bits_addr_beat = ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  assign io_clients_2_grant_valid = ClientTileLinkNetworkPort_2_io_client_grant_valid;
  assign io_clients_2_acquire_ready = ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  ClientTileLinkNetworkPort_0 ClientTileLinkNetworkPort(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_0_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_0_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_0_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_0_acquire_bits_addr_beat ),
       .io_client_acquire_bits_data( io_clients_0_acquire_bits_data ),
       .io_client_acquire_bits_is_builtin_type( io_clients_0_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_0_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_0_acquire_bits_union ),
       .io_client_grant_ready( io_clients_0_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_io_client_grant_bits_data ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_io_client_grant_bits_g_type ),
       .io_client_probe_ready( io_clients_0_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_io_client_release_ready ),
       .io_client_release_valid( io_clients_0_release_valid ),
       .io_client_release_bits_addr_block( io_clients_0_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_0_release_bits_client_xact_id ),
       .io_client_release_bits_addr_beat( io_clients_0_release_bits_addr_beat ),
       .io_client_release_bits_data( io_clients_0_release_bits_data ),
       .io_client_release_bits_r_type( io_clients_0_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_0_release_bits_voluntary ),
       .io_network_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_network_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_0_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_manager_grant_valid( T17 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_finish_ready( RRArbiter_io_in_0_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_manager_probe_valid( T16 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary )
  );
  ClientTileLinkNetworkPort_1 ClientTileLinkNetworkPort_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_1_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_1_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_1_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_1_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_1_acquire_bits_addr_beat ),
       .io_client_acquire_bits_data( io_clients_1_acquire_bits_data ),
       .io_client_acquire_bits_is_builtin_type( io_clients_1_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_1_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_1_acquire_bits_union ),
       .io_client_grant_ready( io_clients_1_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_1_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_1_io_client_grant_bits_data ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type ),
       .io_client_probe_ready( io_clients_1_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_1_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_1_io_client_release_ready ),
       .io_client_release_valid( io_clients_1_release_valid ),
       .io_client_release_bits_addr_block( io_clients_1_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_1_release_bits_client_xact_id ),
       .io_client_release_bits_addr_beat( io_clients_1_release_bits_addr_beat ),
       .io_client_release_bits_data( io_clients_1_release_bits_data ),
       .io_client_release_bits_r_type( io_clients_1_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_1_release_bits_voluntary ),
       .io_network_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_network_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_1_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_manager_grant_valid( T15 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_finish_ready( RRArbiter_io_in_1_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_manager_probe_valid( T14 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary )
  );
  ClientTileLinkNetworkPort_2 ClientTileLinkNetworkPort_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_2_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_2_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_2_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_2_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_2_acquire_bits_addr_beat ),
       .io_client_acquire_bits_data( io_clients_2_acquire_bits_data ),
       .io_client_acquire_bits_is_builtin_type( io_clients_2_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_2_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_2_acquire_bits_union ),
       .io_client_grant_ready( io_clients_2_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_2_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_2_io_client_grant_bits_data ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type ),
       .io_client_probe_ready( io_clients_2_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_2_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_2_io_client_release_ready ),
       .io_client_release_valid( io_clients_2_release_valid ),
       .io_client_release_bits_addr_block( io_clients_2_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_2_release_bits_client_xact_id ),
       .io_client_release_bits_addr_beat( io_clients_2_release_bits_addr_beat ),
       .io_client_release_bits_data( io_clients_2_release_bits_data ),
       .io_client_release_bits_r_type( io_clients_2_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_2_release_bits_voluntary ),
       .io_network_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_network_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_2_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_2_io_manager_grant_ready ),
       .io_manager_grant_valid( T13 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_finish_ready( RRArbiter_io_in_2_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_2_io_manager_probe_ready ),
       .io_manager_probe_valid( T12 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary )
  );
  ManagerTileLinkNetworkPort_0 ManagerTileLinkNetworkPort(
       .io_manager_acquire_ready( io_managers_0_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_0_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_0_grant_bits_addr_beat ),
       .io_manager_grant_bits_data( io_managers_0_grant_bits_data ),
       .io_manager_grant_bits_client_xact_id( io_managers_0_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_0_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_0_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_0_grant_bits_g_type ),
       .io_manager_grant_bits_client_id( io_managers_0_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_0_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_0_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_0_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_0_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_0_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_0_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_io_manager_release_valid ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_io_manager_release_bits_data ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_io_manager_release_bits_r_type ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_network_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_3(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_client_acquire_valid( LockingRRArbiter_io_out_valid ),
       .io_client_acquire_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_client_acquire_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_client_grant_ready( T6 ),
       .io_client_grant_valid( TileLinkEnqueuer_3_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_client_finish_valid( RRArbiter_io_out_valid ),
       .io_client_finish_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_client_finish_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id ),
       .io_client_probe_ready( T0 ),
       .io_client_probe_valid( TileLinkEnqueuer_3_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_client_release_valid( LockingRRArbiter_1_io_out_valid ),
       .io_client_release_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_client_release_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_client_release_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary )
  );
  LockingRRArbiter_0 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_in_2_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_in_1_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_in_0_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data ),
       .io_in_2_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_in_2_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_in_1_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_in_1_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_in_0_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_in_0_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary )
       //.io_chosen(  )
  );
  RRArbiter_1 RRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( RRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module BroadcastVoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [3:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [9:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[25:0] io_inner_probe_bits_addr_block
    //output[1:0] io_inner_probe_bits_p_type
    //output[1:0] io_inner_probe_bits_client_id
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [3:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[9:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T133;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire oacq_data_done;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] R18;
  wire[1:0] T134;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[9:0] T33;
  wire[9:0] T135;
  wire[1:0] T34;
  wire T35;
  wire[2:0] T36;
  wire T37;
  wire[3:0] T38;
  wire[3:0] T39;
  wire[3:0] T40;
  reg [3:0] data_buffer_0;
  wire[3:0] T41;
  wire[3:0] T42;
  wire T43;
  wire T44;
  wire[3:0] T45;
  wire[1:0] T46;
  wire T47;
  reg  collect_irel_data;
  wire T136;
  wire T48;
  wire T49;
  wire T50;
  wire irel_data_done;
  wire T51;
  wire T52;
  wire T53;
  reg [1:0] R54;
  wire[1:0] T137;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire[1:0] T71;
  reg [3:0] data_buffer_1;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T80;
  reg [3:0] data_buffer_2;
  wire[3:0] T81;
  wire[3:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg [3:0] data_buffer_3;
  wire[3:0] T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire[1:0] T95;
  wire[2:0] T96;
  wire[25:0] T97;
  reg [25:0] xact_addr_block;
  wire[25:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  reg [3:0] irel_data_valid;
  wire[3:0] T138;
  wire[3:0] T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T139;
  wire T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[1:0] T123;
  reg [1:0] xact_client_id;
  wire[1:0] T124;
  wire[3:0] T125;
  wire T126;
  wire[2:0] T127;
  wire T128;
  reg  xact_client_xact_id;
  wire T129;
  wire[3:0] T130;
  wire[1:0] T131;
  wire T132;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    R18 = {1{$random}};
    data_buffer_0 = {1{$random}};
    collect_irel_data = {1{$random}};
    R54 = {1{$random}};
    data_buffer_1 = {1{$random}};
    data_buffer_2 = {1{$random}};
    data_buffer_3 = {1{$random}};
    xact_addr_block = {1{$random}};
    irel_data_valid = {1{$random}};
    xact_client_id = {1{$random}};
    xact_client_xact_id = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_inner_probe_bits_client_id = {1{$random}};
//  assign io_inner_probe_bits_p_type = {1{$random}};
//  assign io_inner_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_has_release_match = io_inner_release_bits_voluntary;
  assign io_has_acquire_match = 1'h0;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = T0;
  assign T0 = T1 ? io_inner_grant_ready : 1'h0;
  assign T1 = 2'h2 == state;
  assign T133 = reset ? 2'h0 : T2;
  assign T2 = T31 ? 2'h0 : T3;
  assign T3 = T29 ? T25 : T4;
  assign T4 = T14 ? 2'h2 : T5;
  assign T5 = T12 ? T6 : state;
  assign T6 = T7 ? 2'h1 : 2'h3;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_inner_release_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_inner_release_bits_r_type;
  assign T11 = 3'h0 == io_inner_release_bits_r_type;
  assign T12 = T13 & io_inner_release_valid;
  assign T13 = 2'h0 == state;
  assign T14 = T24 & oacq_data_done;
  assign oacq_data_done = T22 ? T16 : T15;
  assign T15 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T16 = T21 & T17;
  assign T17 = R18 == 2'h3;
  assign T134 = reset ? 2'h0 : T19;
  assign T19 = T21 ? T20 : R18;
  assign T20 = R18 + 2'h1;
  assign T21 = T15 & T22;
  assign T22 = io_outer_acquire_bits_is_builtin_type & T23;
  assign T23 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T24 = 2'h1 == state;
  assign T25 = T26 ? 2'h3 : 2'h0;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_inner_grant_bits_is_builtin_type & T28;
  assign T28 = io_inner_grant_bits_g_type == 4'h0;
  assign T29 = T1 & T30;
  assign T30 = io_inner_grant_ready & io_inner_grant_valid;
  assign T31 = T32 & io_inner_finish_valid;
  assign T32 = 2'h3 == state;
  assign io_outer_acquire_bits_union = T33;
  assign T33 = T135;
  assign T135 = {8'h0, T34};
  assign T34 = {T35, 1'h1};
  assign T35 = 1'h1;
  assign io_outer_acquire_bits_a_type = T36;
  assign T36 = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T37;
  assign T37 = 1'h1;
  assign io_outer_acquire_bits_data = T38;
  assign T38 = T39;
  assign T39 = T94 ? T80 : T40;
  assign T40 = T78 ? data_buffer_1 : data_buffer_0;
  assign T41 = T68 ? io_inner_release_bits_data : T42;
  assign T42 = T43 ? io_inner_release_bits_data : data_buffer_0;
  assign T43 = T47 & T44;
  assign T44 = T45[1'h0:1'h0];
  assign T45 = 1'h1 << T46;
  assign T46 = io_inner_release_bits_addr_beat;
  assign T47 = collect_irel_data & io_inner_release_valid;
  assign T136 = reset ? 1'h0 : T48;
  assign T48 = T12 ? T63 : T49;
  assign T49 = T50 ? 1'h0 : collect_irel_data;
  assign T50 = collect_irel_data & irel_data_done;
  assign irel_data_done = T58 ? T52 : T51;
  assign T51 = io_inner_release_ready & io_inner_release_valid;
  assign T52 = T57 & T53;
  assign T53 = R54 == 2'h3;
  assign T137 = reset ? 2'h0 : T55;
  assign T55 = T57 ? T56 : R54;
  assign T56 = R54 + 2'h1;
  assign T57 = T51 & T58;
  assign T58 = T60 | T59;
  assign T59 = 3'h2 == io_inner_release_bits_r_type;
  assign T60 = T62 | T61;
  assign T61 = 3'h1 == io_inner_release_bits_r_type;
  assign T62 = 3'h0 == io_inner_release_bits_r_type;
  assign T63 = T65 | T64;
  assign T64 = 3'h2 == io_inner_release_bits_r_type;
  assign T65 = T67 | T66;
  assign T66 = 3'h1 == io_inner_release_bits_r_type;
  assign T67 = 3'h0 == io_inner_release_bits_r_type;
  assign T68 = T12 & T69;
  assign T69 = T70[1'h0:1'h0];
  assign T70 = 1'h1 << T71;
  assign T71 = 2'h0;
  assign T72 = T76 ? io_inner_release_bits_data : T73;
  assign T73 = T74 ? io_inner_release_bits_data : data_buffer_1;
  assign T74 = T47 & T75;
  assign T75 = T45[1'h1:1'h1];
  assign T76 = T12 & T77;
  assign T77 = T70[1'h1:1'h1];
  assign T78 = T79[1'h0:1'h0];
  assign T79 = oacq_data_cnt;
  assign oacq_data_cnt = T22 ? R18 : 2'h0;
  assign T80 = T93 ? data_buffer_3 : data_buffer_2;
  assign T81 = T85 ? io_inner_release_bits_data : T82;
  assign T82 = T83 ? io_inner_release_bits_data : data_buffer_2;
  assign T83 = T47 & T84;
  assign T84 = T45[2'h2:2'h2];
  assign T85 = T12 & T86;
  assign T86 = T70[2'h2:2'h2];
  assign T87 = T91 ? io_inner_release_bits_data : T88;
  assign T88 = T89 ? io_inner_release_bits_data : data_buffer_3;
  assign T89 = T47 & T90;
  assign T90 = T45[2'h3:2'h3];
  assign T91 = T12 & T92;
  assign T92 = T70[2'h3:2'h3];
  assign T93 = T79[1'h0:1'h0];
  assign T94 = T79[1'h1:1'h1];
  assign io_outer_acquire_bits_addr_beat = T95;
  assign T95 = oacq_data_cnt;
  assign io_outer_acquire_bits_client_xact_id = T96;
  assign T96 = 3'h0;
  assign io_outer_acquire_bits_addr_block = T97;
  assign T97 = xact_addr_block;
  assign T98 = T12 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign io_outer_acquire_valid = T99;
  assign T99 = T24 ? T100 : 1'h0;
  assign T100 = T121 | T101;
  assign T101 = T106 & T102;
  assign T102 = T103 - 1'h1;
  assign T103 = 1'h1 << T104;
  assign T104 = T105 + 2'h1;
  assign T105 = oacq_data_cnt - oacq_data_cnt;
  assign T106 = irel_data_valid >> oacq_data_cnt;
  assign T138 = reset ? 4'h0 : T107;
  assign T107 = T12 ? T115 : T108;
  assign T108 = T47 ? T109 : irel_data_valid;
  assign T109 = T113 | T110;
  assign T110 = T139 & T111;
  assign T111 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T139 = T112 ? 4'hf : 4'h0;
  assign T112 = 1'h1;
  assign T113 = irel_data_valid & T114;
  assign T114 = ~ T111;
  assign T115 = T116 << io_inner_release_bits_addr_beat;
  assign T116 = T118 | T117;
  assign T117 = 3'h2 == io_inner_release_bits_r_type;
  assign T118 = T120 | T119;
  assign T119 = 3'h1 == io_inner_release_bits_r_type;
  assign T120 = 3'h0 == io_inner_release_bits_r_type;
  assign T121 = collect_irel_data ^ 1'h1;
  assign io_inner_release_ready = T122;
  assign T122 = T13 ? 1'h1 : collect_irel_data;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = T32;
  assign io_inner_grant_bits_client_id = T123;
  assign T123 = xact_client_id;
  assign T124 = T12 ? io_inner_release_bits_client_id : xact_client_id;
  assign io_inner_grant_bits_g_type = T125;
  assign T125 = 4'h0;
  assign io_inner_grant_bits_is_builtin_type = T126;
  assign T126 = 1'h1;
  assign io_inner_grant_bits_manager_xact_id = T127;
  assign T127 = 3'h0;
  assign io_inner_grant_bits_client_xact_id = T128;
  assign T128 = xact_client_xact_id;
  assign T129 = T12 ? io_inner_release_bits_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_data = T130;
  assign T130 = 4'h0;
  assign io_inner_grant_bits_addr_beat = T131;
  assign T131 = 2'h0;
  assign io_inner_grant_valid = T132;
  assign T132 = T1 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T31) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= T25;
    end else if(T14) begin
      state <= 2'h2;
    end else if(T12) begin
      state <= T6;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T21) begin
      R18 <= T20;
    end
    if(T68) begin
      data_buffer_0 <= io_inner_release_bits_data;
    end else if(T43) begin
      data_buffer_0 <= io_inner_release_bits_data;
    end
    if(reset) begin
      collect_irel_data <= 1'h0;
    end else if(T12) begin
      collect_irel_data <= T63;
    end else if(T50) begin
      collect_irel_data <= 1'h0;
    end
    if(reset) begin
      R54 <= 2'h0;
    end else if(T57) begin
      R54 <= T56;
    end
    if(T76) begin
      data_buffer_1 <= io_inner_release_bits_data;
    end else if(T74) begin
      data_buffer_1 <= io_inner_release_bits_data;
    end
    if(T85) begin
      data_buffer_2 <= io_inner_release_bits_data;
    end else if(T83) begin
      data_buffer_2 <= io_inner_release_bits_data;
    end
    if(T91) begin
      data_buffer_3 <= io_inner_release_bits_data;
    end else if(T89) begin
      data_buffer_3 <= io_inner_release_bits_data;
    end
    if(T12) begin
      xact_addr_block <= io_inner_release_bits_addr_block;
    end
    if(reset) begin
      irel_data_valid <= 4'h0;
    end else if(T12) begin
      irel_data_valid <= T115;
    end else if(T47) begin
      irel_data_valid <= T109;
    end
    if(T12) begin
      xact_client_id <= io_inner_release_bits_client_id;
    end
    if(T12) begin
      xact_client_xact_id <= io_inner_release_bits_client_xact_id;
    end
  end
endmodule

module BroadcastAcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [3:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [9:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [3:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[9:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [2:0] state;
  wire[2:0] T361;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire pending_outer_read_;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T362;
  wire[2:0] T22;
  wire[2:0] T363;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire pending_outer_write_;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[3:0] mask_incoherent;
  wire[3:0] T364;
  wire T48;
  wire T49;
  wire[3:0] mask_self;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T365;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T366;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire pending_outer_read;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire pending_outer_write;
  wire T66;
  wire T67;
  reg [2:0] xact_a_type;
  wire[2:0] T68;
  wire T69;
  wire T70;
  wire T71;
  reg  xact_is_builtin_type;
  wire T72;
  wire T73;
  wire T74;
  reg  release_count;
  wire T367;
  wire[2:0] T368;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T369;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T370;
  wire T83;
  wire[2:0] T371;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T372;
  wire T87;
  wire T88;
  wire[2:0] T373;
  wire T89;
  wire[2:0] T374;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire oacq_data_done;
  wire T101;
  wire T102;
  wire T103;
  reg [1:0] R104;
  wire[1:0] T375;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire ignt_data_done;
  wire T127;
  wire T128;
  wire T129;
  reg [1:0] R130;
  wire[1:0] T376;
  wire[1:0] T131;
  wire[1:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[2:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  reg[0:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  xact_client_xact_id;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  reg  collect_iacq_data;
  wire T377;
  wire T157;
  wire T158;
  wire T159;
  wire iacq_data_done;
  wire T160;
  wire T161;
  wire T162;
  reg [1:0] R163;
  wire[1:0] T378;
  wire[1:0] T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  reg[0:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg [1:0] xact_client_id;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg [25:0] xact_addr_block;
  wire[25:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg  pending_ognt_ack;
  wire T379;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[9:0] T213;
  wire[9:0] T214;
  wire[9:0] T215;
  wire[9:0] outer_write_rel_union;
  wire[9:0] T380;
  wire[1:0] T216;
  wire T217;
  wire[9:0] outer_write_acq_union;
  wire[9:0] T381;
  wire[1:0] T218;
  wire T219;
  wire[9:0] outer_read_union;
  wire[2:0] T220;
  wire[2:0] T221;
  wire[2:0] T222;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[2:0] outer_read_a_type;
  wire T223;
  wire T224;
  wire T225;
  wire outer_write_rel_is_builtin_type;
  wire outer_write_acq_is_builtin_type;
  wire outer_read_is_builtin_type;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T229;
  wire[3:0] T230;
  reg [3:0] data_buffer_0;
  wire[3:0] T231;
  wire[3:0] T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire[3:0] T240;
  wire[1:0] T241;
  reg [3:0] data_buffer_1;
  wire[3:0] T242;
  wire[3:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T250;
  reg [3:0] data_buffer_2;
  wire[3:0] T251;
  wire[3:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  reg [3:0] data_buffer_3;
  wire[3:0] T257;
  wire[3:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] outer_read_data;
  wire[1:0] T265;
  wire[1:0] T266;
  wire[1:0] T267;
  wire[1:0] outer_write_rel_addr_beat;
  wire[1:0] outer_write_acq_addr_beat;
  wire[1:0] outer_read_addr_beat;
  wire[2:0] T268;
  wire[2:0] T269;
  wire[2:0] T270;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[25:0] T271;
  wire[25:0] T272;
  wire[25:0] T273;
  wire[25:0] outer_write_rel_addr_block;
  wire[25:0] outer_write_acq_addr_block;
  wire[25:0] outer_read_addr_block;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[1:0] T280;
  wire[1:0] T281;
  wire T282;
  reg [3:0] iacq_data_valid;
  wire[3:0] T382;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[3:0] T286;
  wire[3:0] T287;
  wire[3:0] T383;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire[1:0] T310;
  wire[1:0] T384;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire[25:0] T333;
  wire T334;
  wire T335;
  reg  pending_probes;
  wire T385;
  wire[3:0] T386;
  wire[3:0] T311;
  wire[3:0] T312;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire[1:0] T389;
  wire T316;
  wire[1:0] T336;
  wire[3:0] T337;
  wire[3:0] T390;
  wire[2:0] T338;
  wire[2:0] T391;
  wire[1:0] T339;
  wire T340;
  wire[2:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[2:0] T354;
  wire T355;
  wire[3:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R104 = {1{$random}};
    R130 = {1{$random}};
    T148 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R163 = {1{$random}};
    T172 = 1'b0;
    xact_client_id = {1{$random}};
    T182 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    data_buffer_0 = {1{$random}};
    data_buffer_1 = {1{$random}};
    data_buffer_2 = {1{$random}};
    data_buffer_3 = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T7 & T6;
  assign T6 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T7 = state == 3'h0;
  assign T361 = reset ? 3'h0 : T8;
  assign T8 = T146 ? 3'h0 : T9;
  assign T9 = T144 ? T140 : T10;
  assign T10 = T126 ? T122 : T11;
  assign T11 = T119 ? 3'h5 : T12;
  assign T12 = T117 ? T116 : T13;
  assign T13 = T114 ? T112 : T14;
  assign T14 = T73 ? T58 : T15;
  assign T15 = T56 ? T16 : state;
  assign T16 = T47 ? 3'h1 : T17;
  assign T17 = pending_outer_write_ ? 3'h3 : T18;
  assign T18 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T41 ? T38 : T19;
  assign T19 = T37 | T20;
  assign T20 = 4'h1 == T21;
  assign T21 = T362;
  assign T362 = {1'h0, T22};
  assign T22 = io_inner_acquire_bits_is_builtin_type ? T25 : T363;
  assign T363 = {1'h0, T23};
  assign T23 = T24 ? 2'h0 : 2'h1;
  assign T24 = io_inner_acquire_bits_a_type == 3'h0;
  assign T25 = T36 ? 3'h4 : T26;
  assign T26 = T35 ? 3'h5 : T27;
  assign T27 = T34 ? 3'h3 : T28;
  assign T28 = T33 ? 3'h3 : T29;
  assign T29 = T32 ? 3'h4 : T30;
  assign T30 = T31 ? 3'h1 : 3'h3;
  assign T31 = io_inner_acquire_bits_a_type == 3'h5;
  assign T32 = io_inner_acquire_bits_a_type == 3'h4;
  assign T33 = io_inner_acquire_bits_a_type == 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h2;
  assign T35 = io_inner_acquire_bits_a_type == 3'h1;
  assign T36 = io_inner_acquire_bits_a_type == 3'h0;
  assign T37 = 4'h0 == T21;
  assign T38 = T40 | T39;
  assign T39 = 4'h4 == T21;
  assign T40 = 4'h5 == T21;
  assign T41 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T42;
  assign T42 = T44 | T43;
  assign T43 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T46 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T47 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T364;
  assign T364 = {3'h0, T48};
  assign T48 = ~ T49;
  assign T49 = io_incoherent_0;
  assign mask_self = T53 | T50;
  assign T50 = T365 & T51;
  assign T51 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T365 = T52 ? 4'hf : 4'h0;
  assign T52 = 1'h0;
  assign T53 = T366 & T54;
  assign T54 = ~ T51;
  assign T366 = {3'h0, T55};
  assign T55 = 1'h1;
  assign T56 = T57 & io_inner_acquire_valid;
  assign T57 = 3'h0 == state;
  assign T58 = pending_outer_write ? 3'h3 : T59;
  assign T59 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T63 : T60;
  assign T60 = T62 | T61;
  assign T61 = 4'h1 == io_inner_grant_bits_g_type;
  assign T62 = 4'h0 == io_inner_grant_bits_g_type;
  assign T63 = T65 | T64;
  assign T64 = 4'h4 == io_inner_grant_bits_g_type;
  assign T65 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T66;
  assign T66 = T69 | T67;
  assign T67 = 3'h4 == xact_a_type;
  assign T68 = T56 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T69 = T71 | T70;
  assign T70 = 3'h3 == xact_a_type;
  assign T71 = 3'h2 == xact_a_type;
  assign T72 = T56 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T73 = T100 & T74;
  assign T74 = release_count == 1'h1;
  assign T367 = T368[1'h0:1'h0];
  assign T368 = reset ? 3'h0 : T75;
  assign T75 = T91 ? T374 : T76;
  assign T76 = T100 ? T373 : T77;
  assign T77 = T88 ? T78 : T369;
  assign T369 = {2'h0, release_count};
  assign T78 = T371 + T79;
  assign T79 = {1'h0, T80};
  assign T80 = T370 + T81;
  assign T81 = {1'h0, T82};
  assign T82 = mask_incoherent[2'h3:2'h3];
  assign T370 = {1'h0, T83};
  assign T83 = mask_incoherent[2'h2:2'h2];
  assign T371 = {1'h0, T84};
  assign T84 = T372 + T85;
  assign T85 = {1'h0, T86};
  assign T86 = mask_incoherent[1'h1:1'h1];
  assign T372 = {1'h0, T87};
  assign T87 = mask_incoherent[1'h0:1'h0];
  assign T88 = T56 & T47;
  assign T373 = {2'h0, T89};
  assign T89 = release_count - 1'h1;
  assign T374 = {2'h0, T90};
  assign T90 = release_count - 1'h1;
  assign T91 = T98 & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T95 | T94;
  assign T94 = 3'h2 == io_inner_release_bits_r_type;
  assign T95 = T97 | T96;
  assign T96 = 3'h1 == io_inner_release_bits_r_type;
  assign T97 = 3'h0 == io_inner_release_bits_r_type;
  assign T98 = T99 & io_inner_release_valid;
  assign T99 = 3'h1 == state;
  assign T100 = T110 & oacq_data_done;
  assign oacq_data_done = T108 ? T102 : T101;
  assign T101 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T102 = T107 & T103;
  assign T103 = R104 == 2'h3;
  assign T375 = reset ? 2'h0 : T105;
  assign T105 = T107 ? T106 : R104;
  assign T106 = R104 + 2'h1;
  assign T107 = T101 & T108;
  assign T108 = io_outer_acquire_bits_is_builtin_type & T109;
  assign T109 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T110 = T111 & io_outer_acquire_ready;
  assign T111 = T98 & T93;
  assign T112 = pending_outer_write ? 3'h3 : T113;
  assign T113 = pending_outer_read ? 3'h2 : 3'h4;
  assign T114 = T91 & T115;
  assign T115 = release_count == 1'h1;
  assign T116 = pending_outer_read ? 3'h2 : 3'h5;
  assign T117 = T118 & oacq_data_done;
  assign T118 = 3'h3 == state;
  assign T119 = T121 & T120;
  assign T120 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T121 = 3'h2 == state;
  assign T122 = T123 ? 3'h6 : 3'h0;
  assign T123 = T124 ^ 1'h1;
  assign T124 = io_inner_grant_bits_is_builtin_type & T125;
  assign T125 = io_inner_grant_bits_g_type == 4'h0;
  assign T126 = T139 & ignt_data_done;
  assign ignt_data_done = T134 ? T128 : T127;
  assign T127 = io_inner_grant_ready & io_inner_grant_valid;
  assign T128 = T133 & T129;
  assign T129 = R130 == 2'h3;
  assign T376 = reset ? 2'h0 : T131;
  assign T131 = T133 ? T132 : R130;
  assign T132 = R130 + 2'h1;
  assign T133 = T127 & T134;
  assign T134 = io_inner_grant_bits_is_builtin_type ? T138 : T135;
  assign T135 = T137 | T136;
  assign T136 = 4'h1 == io_inner_grant_bits_g_type;
  assign T137 = 4'h0 == io_inner_grant_bits_g_type;
  assign T138 = 4'h5 == io_inner_grant_bits_g_type;
  assign T139 = 3'h5 == state;
  assign T140 = T141 ? 3'h6 : 3'h0;
  assign T141 = T142 ^ 1'h1;
  assign T142 = io_inner_grant_bits_is_builtin_type & T143;
  assign T143 = io_inner_grant_bits_g_type == 4'h0;
  assign T144 = T145 & io_inner_grant_ready;
  assign T145 = 3'h4 == state;
  assign T146 = T147 & io_inner_finish_valid;
  assign T147 = 3'h6 == state;
  assign T149 = T150 | reset;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T154 & T152;
  assign T152 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T153 = T56 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T154 = T156 & T155;
  assign T155 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T156 = T171 & collect_iacq_data;
  assign T377 = reset ? 1'h0 : T157;
  assign T157 = T56 ? T169 : T158;
  assign T158 = T159 ? 1'h0 : collect_iacq_data;
  assign T159 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T167 ? T161 : T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T166 & T162;
  assign T162 = R163 == 2'h3;
  assign T378 = reset ? 2'h0 : T164;
  assign T164 = T166 ? T165 : R163;
  assign T165 = R163 + 2'h1;
  assign T166 = T160 & T167;
  assign T167 = io_inner_acquire_bits_is_builtin_type & T168;
  assign T168 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T169 = io_inner_acquire_bits_is_builtin_type & T170;
  assign T170 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T171 = state != 3'h0;
  assign T173 = T174 | reset;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T178 & T176;
  assign T176 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T177 = T56 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T178 = T180 & T179;
  assign T179 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T180 = T181 & collect_iacq_data;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T193 & T186;
  assign T186 = T188 | T187;
  assign T187 = 3'h5 == xact_a_type;
  assign T188 = T190 | T189;
  assign T189 = 3'h4 == xact_a_type;
  assign T190 = T192 | T191;
  assign T191 = 3'h2 == xact_a_type;
  assign T192 = 3'h0 == xact_a_type;
  assign T193 = T194 & xact_is_builtin_type;
  assign T194 = state != 3'h0;
  assign io_has_release_match = T195;
  assign T195 = T197 & T196;
  assign T196 = state == 3'h1;
  assign T197 = T199 & T198;
  assign T198 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T199 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T200 = T56 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T201;
  assign T201 = T202 & collect_iacq_data;
  assign T202 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T203;
  assign T203 = T205 & T204;
  assign T204 = collect_iacq_data ^ 1'h1;
  assign T205 = T207 & T206;
  assign T206 = state != 3'h0;
  assign T207 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T208;
  assign T208 = T139 ? io_inner_grant_ready : pending_ognt_ack;
  assign T379 = reset ? 1'h0 : T209;
  assign T209 = T117 ? 1'h1 : T210;
  assign T210 = T100 ? 1'h1 : T211;
  assign T211 = T212 ? 1'h0 : pending_ognt_ack;
  assign T212 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_union = T213;
  assign T213 = T121 ? outer_read_union : T214;
  assign T214 = T118 ? outer_write_acq_union : T215;
  assign T215 = T111 ? outer_write_rel_union : outer_read_union;
  assign outer_write_rel_union = T380;
  assign T380 = {8'h0, T216};
  assign T216 = {T217, 1'h1};
  assign T217 = 1'h1;
  assign outer_write_acq_union = T381;
  assign T381 = {8'h0, T218};
  assign T218 = {T219, 1'h1};
  assign T219 = 1'h1;
  assign outer_read_union = 10'h1c1;
  assign io_outer_acquire_bits_a_type = T220;
  assign T220 = T121 ? outer_read_a_type : T221;
  assign T221 = T118 ? outer_write_acq_a_type : T222;
  assign T222 = T111 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign outer_read_a_type = 3'h1;
  assign io_outer_acquire_bits_is_builtin_type = T223;
  assign T223 = T121 ? outer_read_is_builtin_type : T224;
  assign T224 = T118 ? outer_write_acq_is_builtin_type : T225;
  assign T225 = T111 ? outer_write_rel_is_builtin_type : outer_read_is_builtin_type;
  assign outer_write_rel_is_builtin_type = 1'h1;
  assign outer_write_acq_is_builtin_type = 1'h1;
  assign outer_read_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_data = T226;
  assign T226 = T121 ? outer_read_data : T227;
  assign T227 = T118 ? outer_write_acq_data : T228;
  assign T228 = T111 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_data;
  assign outer_write_acq_data = T229;
  assign T229 = T264 ? T250 : T230;
  assign T230 = T248 ? data_buffer_1 : data_buffer_0;
  assign T231 = T238 ? io_inner_acquire_bits_data : T232;
  assign T232 = T233 ? io_inner_acquire_bits_data : data_buffer_0;
  assign T233 = T237 & T234;
  assign T234 = T235[1'h0:1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = io_inner_acquire_bits_addr_beat;
  assign T237 = collect_iacq_data & io_inner_acquire_valid;
  assign T238 = T56 & T239;
  assign T239 = T240[1'h0:1'h0];
  assign T240 = 1'h1 << T241;
  assign T241 = 2'h0;
  assign T242 = T246 ? io_inner_acquire_bits_data : T243;
  assign T243 = T244 ? io_inner_acquire_bits_data : data_buffer_1;
  assign T244 = T237 & T245;
  assign T245 = T235[1'h1:1'h1];
  assign T246 = T56 & T247;
  assign T247 = T240[1'h1:1'h1];
  assign T248 = T249[1'h0:1'h0];
  assign T249 = oacq_data_cnt;
  assign oacq_data_cnt = T108 ? R104 : 2'h0;
  assign T250 = T263 ? data_buffer_3 : data_buffer_2;
  assign T251 = T255 ? io_inner_acquire_bits_data : T252;
  assign T252 = T253 ? io_inner_acquire_bits_data : data_buffer_2;
  assign T253 = T237 & T254;
  assign T254 = T235[2'h2:2'h2];
  assign T255 = T56 & T256;
  assign T256 = T240[2'h2:2'h2];
  assign T257 = T261 ? io_inner_acquire_bits_data : T258;
  assign T258 = T259 ? io_inner_acquire_bits_data : data_buffer_3;
  assign T259 = T237 & T260;
  assign T260 = T235[2'h3:2'h3];
  assign T261 = T56 & T262;
  assign T262 = T240[2'h3:2'h3];
  assign T263 = T249[1'h0:1'h0];
  assign T264 = T249[1'h1:1'h1];
  assign outer_read_data = 4'h0;
  assign io_outer_acquire_bits_addr_beat = T265;
  assign T265 = T121 ? outer_read_addr_beat : T266;
  assign T266 = T118 ? outer_write_acq_addr_beat : T267;
  assign T267 = T111 ? outer_write_rel_addr_beat : outer_read_addr_beat;
  assign outer_write_rel_addr_beat = io_inner_release_bits_addr_beat;
  assign outer_write_acq_addr_beat = oacq_data_cnt;
  assign outer_read_addr_beat = 2'h0;
  assign io_outer_acquire_bits_client_xact_id = T268;
  assign T268 = T121 ? outer_read_client_xact_id : T269;
  assign T269 = T118 ? outer_write_acq_client_xact_id : T270;
  assign T270 = T111 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h1;
  assign outer_write_acq_client_xact_id = 3'h1;
  assign outer_read_client_xact_id = 3'h1;
  assign io_outer_acquire_bits_addr_block = T271;
  assign T271 = T121 ? outer_read_addr_block : T272;
  assign T272 = T118 ? outer_write_acq_addr_block : T273;
  assign T273 = T111 ? outer_write_rel_addr_block : outer_read_addr_block;
  assign outer_write_rel_addr_block = xact_addr_block;
  assign outer_write_acq_addr_block = xact_addr_block;
  assign outer_read_addr_block = xact_addr_block;
  assign io_outer_acquire_valid = T274;
  assign T274 = T121 ? T301 : T275;
  assign T275 = T118 ? T276 : T111;
  assign T276 = T298 | T277;
  assign T277 = T282 & T278;
  assign T278 = T279 - 1'h1;
  assign T279 = 1'h1 << T280;
  assign T280 = T281 + 2'h1;
  assign T281 = oacq_data_cnt - oacq_data_cnt;
  assign T282 = iacq_data_valid >> oacq_data_cnt;
  assign T382 = reset ? 4'h0 : T283;
  assign T283 = T56 ? T291 : T284;
  assign T284 = T237 ? T285 : iacq_data_valid;
  assign T285 = T289 | T286;
  assign T286 = T383 & T287;
  assign T287 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T383 = T288 ? 4'hf : 4'h0;
  assign T288 = 1'h1;
  assign T289 = iacq_data_valid & T290;
  assign T290 = ~ T287;
  assign T291 = T292 << io_inner_acquire_bits_addr_beat;
  assign T292 = io_inner_acquire_bits_is_builtin_type & T293;
  assign T293 = T295 | T294;
  assign T294 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T295 = T297 | T296;
  assign T296 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T297 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T298 = T300 | T299;
  assign T299 = collect_iacq_data ^ 1'h1;
  assign T300 = pending_ognt_ack ^ 1'h1;
  assign T301 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T302;
  assign T302 = T99 ? T303 : 1'h0;
  assign T303 = T304 | io_outer_acquire_ready;
  assign T304 = T305 ^ 1'h1;
  assign T305 = T307 | T306;
  assign T306 = 3'h2 == io_inner_release_bits_r_type;
  assign T307 = T309 | T308;
  assign T308 = 3'h1 == io_inner_release_bits_r_type;
  assign T309 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T310;
  assign T310 = T384;
  assign T384 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T317;
  assign T317 = T318;
  assign T318 = xact_is_builtin_type ? T323 : T319;
  assign T319 = T322 ? 2'h1 : T320;
  assign T320 = T321 ? 2'h0 : 2'h2;
  assign T321 = xact_a_type == 3'h1;
  assign T322 = xact_a_type == 3'h0;
  assign T323 = T332 ? 2'h2 : T324;
  assign T324 = T331 ? 2'h0 : T325;
  assign T325 = T330 ? 2'h2 : T326;
  assign T326 = T329 ? 2'h0 : T327;
  assign T327 = T328 ? 2'h0 : 2'h2;
  assign T328 = xact_a_type == 3'h4;
  assign T329 = xact_a_type == 3'h2;
  assign T330 = xact_a_type == 3'h0;
  assign T331 = xact_a_type == 3'h3;
  assign T332 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T333;
  assign T333 = xact_addr_block;
  assign io_inner_probe_valid = T334;
  assign T334 = T99 ? T335 : 1'h0;
  assign T335 = pending_probes != 1'h0;
  assign T385 = T386[1'h0:1'h0];
  assign T386 = reset ? 4'h0 : T311;
  assign T311 = T316 ? T388 : T312;
  assign T312 = T88 ? mask_incoherent : T387;
  assign T387 = {3'h0, pending_probes};
  assign T388 = {2'h0, T313};
  assign T313 = T389 & T314;
  assign T314 = ~ T315;
  assign T315 = 1'h1 << 1'h0;
  assign T389 = {1'h0, pending_probes};
  assign T316 = T99 & io_inner_probe_ready;
  assign io_inner_finish_ready = T147;
  assign io_inner_grant_bits_client_id = T336;
  assign T336 = xact_client_id;
  assign io_inner_grant_bits_g_type = T337;
  assign T337 = T390;
  assign T390 = {1'h0, T338};
  assign T338 = xact_is_builtin_type ? T341 : T391;
  assign T391 = {1'h0, T339};
  assign T339 = T340 ? 2'h0 : 2'h1;
  assign T340 = xact_a_type == 3'h0;
  assign T341 = T352 ? 3'h4 : T342;
  assign T342 = T351 ? 3'h5 : T343;
  assign T343 = T350 ? 3'h3 : T344;
  assign T344 = T349 ? 3'h3 : T345;
  assign T345 = T348 ? 3'h4 : T346;
  assign T346 = T347 ? 3'h1 : 3'h3;
  assign T347 = xact_a_type == 3'h5;
  assign T348 = xact_a_type == 3'h4;
  assign T349 = xact_a_type == 3'h3;
  assign T350 = xact_a_type == 3'h2;
  assign T351 = xact_a_type == 3'h1;
  assign T352 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T353;
  assign T353 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T354;
  assign T354 = 3'h1;
  assign io_inner_grant_bits_client_xact_id = T355;
  assign T355 = xact_client_xact_id;
  assign io_inner_grant_bits_data = T356;
  assign T356 = 4'h0;
  assign io_inner_grant_bits_addr_beat = T357;
  assign T357 = 2'h0;
  assign io_inner_grant_valid = T358;
  assign T358 = T145 ? 1'h1 : T359;
  assign T359 = T139 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T360;
  assign T360 = T57 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics, subblock Gets/Puts, or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T172 <= 1'b1;
  if(!T173 && T172 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T148 <= 1'b1;
  if(!T149 && T148 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T146) begin
      state <= 3'h0;
    end else if(T144) begin
      state <= T140;
    end else if(T126) begin
      state <= T122;
    end else if(T119) begin
      state <= 3'h5;
    end else if(T117) begin
      state <= T116;
    end else if(T114) begin
      state <= T112;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T16;
    end
    if(T56) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T56) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T367;
    if(reset) begin
      R104 <= 2'h0;
    end else if(T107) begin
      R104 <= T106;
    end
    if(reset) begin
      R130 <= 2'h0;
    end else if(T133) begin
      R130 <= T132;
    end
    if(T56) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T56) begin
      collect_iacq_data <= T169;
    end else if(T159) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R163 <= 2'h0;
    end else if(T166) begin
      R163 <= T165;
    end
    if(T56) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T56) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T117) begin
      pending_ognt_ack <= 1'h1;
    end else if(T100) begin
      pending_ognt_ack <= 1'h1;
    end else if(T212) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T238) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T233) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T246) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T244) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T255) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T253) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T261) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T259) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T56) begin
      iacq_data_valid <= T291;
    end else if(T237) begin
      iacq_data_valid <= T285;
    end
    pending_probes <= T385;
  end
endmodule

module BroadcastAcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [3:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [9:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [3:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[9:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [2:0] state;
  wire[2:0] T361;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire pending_outer_read_;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T362;
  wire[2:0] T22;
  wire[2:0] T363;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire pending_outer_write_;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[3:0] mask_incoherent;
  wire[3:0] T364;
  wire T48;
  wire T49;
  wire[3:0] mask_self;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T365;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T366;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire pending_outer_read;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire pending_outer_write;
  wire T66;
  wire T67;
  reg [2:0] xact_a_type;
  wire[2:0] T68;
  wire T69;
  wire T70;
  wire T71;
  reg  xact_is_builtin_type;
  wire T72;
  wire T73;
  wire T74;
  reg  release_count;
  wire T367;
  wire[2:0] T368;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T369;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T370;
  wire T83;
  wire[2:0] T371;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T372;
  wire T87;
  wire T88;
  wire[2:0] T373;
  wire T89;
  wire[2:0] T374;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire oacq_data_done;
  wire T101;
  wire T102;
  wire T103;
  reg [1:0] R104;
  wire[1:0] T375;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire ignt_data_done;
  wire T127;
  wire T128;
  wire T129;
  reg [1:0] R130;
  wire[1:0] T376;
  wire[1:0] T131;
  wire[1:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[2:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  reg[0:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  xact_client_xact_id;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  reg  collect_iacq_data;
  wire T377;
  wire T157;
  wire T158;
  wire T159;
  wire iacq_data_done;
  wire T160;
  wire T161;
  wire T162;
  reg [1:0] R163;
  wire[1:0] T378;
  wire[1:0] T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  reg[0:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg [1:0] xact_client_id;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg [25:0] xact_addr_block;
  wire[25:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg  pending_ognt_ack;
  wire T379;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[9:0] T213;
  wire[9:0] T214;
  wire[9:0] T215;
  wire[9:0] outer_write_rel_union;
  wire[9:0] T380;
  wire[1:0] T216;
  wire T217;
  wire[9:0] outer_write_acq_union;
  wire[9:0] T381;
  wire[1:0] T218;
  wire T219;
  wire[9:0] outer_read_union;
  wire[2:0] T220;
  wire[2:0] T221;
  wire[2:0] T222;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[2:0] outer_read_a_type;
  wire T223;
  wire T224;
  wire T225;
  wire outer_write_rel_is_builtin_type;
  wire outer_write_acq_is_builtin_type;
  wire outer_read_is_builtin_type;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T229;
  wire[3:0] T230;
  reg [3:0] data_buffer_0;
  wire[3:0] T231;
  wire[3:0] T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire[3:0] T240;
  wire[1:0] T241;
  reg [3:0] data_buffer_1;
  wire[3:0] T242;
  wire[3:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T250;
  reg [3:0] data_buffer_2;
  wire[3:0] T251;
  wire[3:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  reg [3:0] data_buffer_3;
  wire[3:0] T257;
  wire[3:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] outer_read_data;
  wire[1:0] T265;
  wire[1:0] T266;
  wire[1:0] T267;
  wire[1:0] outer_write_rel_addr_beat;
  wire[1:0] outer_write_acq_addr_beat;
  wire[1:0] outer_read_addr_beat;
  wire[2:0] T268;
  wire[2:0] T269;
  wire[2:0] T270;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[25:0] T271;
  wire[25:0] T272;
  wire[25:0] T273;
  wire[25:0] outer_write_rel_addr_block;
  wire[25:0] outer_write_acq_addr_block;
  wire[25:0] outer_read_addr_block;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[1:0] T280;
  wire[1:0] T281;
  wire T282;
  reg [3:0] iacq_data_valid;
  wire[3:0] T382;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[3:0] T286;
  wire[3:0] T287;
  wire[3:0] T383;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire[1:0] T310;
  wire[1:0] T384;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire[25:0] T333;
  wire T334;
  wire T335;
  reg  pending_probes;
  wire T385;
  wire[3:0] T386;
  wire[3:0] T311;
  wire[3:0] T312;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire[1:0] T389;
  wire T316;
  wire[1:0] T336;
  wire[3:0] T337;
  wire[3:0] T390;
  wire[2:0] T338;
  wire[2:0] T391;
  wire[1:0] T339;
  wire T340;
  wire[2:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[2:0] T354;
  wire T355;
  wire[3:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R104 = {1{$random}};
    R130 = {1{$random}};
    T148 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R163 = {1{$random}};
    T172 = 1'b0;
    xact_client_id = {1{$random}};
    T182 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    data_buffer_0 = {1{$random}};
    data_buffer_1 = {1{$random}};
    data_buffer_2 = {1{$random}};
    data_buffer_3 = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T7 & T6;
  assign T6 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T7 = state == 3'h0;
  assign T361 = reset ? 3'h0 : T8;
  assign T8 = T146 ? 3'h0 : T9;
  assign T9 = T144 ? T140 : T10;
  assign T10 = T126 ? T122 : T11;
  assign T11 = T119 ? 3'h5 : T12;
  assign T12 = T117 ? T116 : T13;
  assign T13 = T114 ? T112 : T14;
  assign T14 = T73 ? T58 : T15;
  assign T15 = T56 ? T16 : state;
  assign T16 = T47 ? 3'h1 : T17;
  assign T17 = pending_outer_write_ ? 3'h3 : T18;
  assign T18 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T41 ? T38 : T19;
  assign T19 = T37 | T20;
  assign T20 = 4'h1 == T21;
  assign T21 = T362;
  assign T362 = {1'h0, T22};
  assign T22 = io_inner_acquire_bits_is_builtin_type ? T25 : T363;
  assign T363 = {1'h0, T23};
  assign T23 = T24 ? 2'h0 : 2'h1;
  assign T24 = io_inner_acquire_bits_a_type == 3'h0;
  assign T25 = T36 ? 3'h4 : T26;
  assign T26 = T35 ? 3'h5 : T27;
  assign T27 = T34 ? 3'h3 : T28;
  assign T28 = T33 ? 3'h3 : T29;
  assign T29 = T32 ? 3'h4 : T30;
  assign T30 = T31 ? 3'h1 : 3'h3;
  assign T31 = io_inner_acquire_bits_a_type == 3'h5;
  assign T32 = io_inner_acquire_bits_a_type == 3'h4;
  assign T33 = io_inner_acquire_bits_a_type == 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h2;
  assign T35 = io_inner_acquire_bits_a_type == 3'h1;
  assign T36 = io_inner_acquire_bits_a_type == 3'h0;
  assign T37 = 4'h0 == T21;
  assign T38 = T40 | T39;
  assign T39 = 4'h4 == T21;
  assign T40 = 4'h5 == T21;
  assign T41 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T42;
  assign T42 = T44 | T43;
  assign T43 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T46 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T47 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T364;
  assign T364 = {3'h0, T48};
  assign T48 = ~ T49;
  assign T49 = io_incoherent_0;
  assign mask_self = T53 | T50;
  assign T50 = T365 & T51;
  assign T51 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T365 = T52 ? 4'hf : 4'h0;
  assign T52 = 1'h0;
  assign T53 = T366 & T54;
  assign T54 = ~ T51;
  assign T366 = {3'h0, T55};
  assign T55 = 1'h1;
  assign T56 = T57 & io_inner_acquire_valid;
  assign T57 = 3'h0 == state;
  assign T58 = pending_outer_write ? 3'h3 : T59;
  assign T59 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T63 : T60;
  assign T60 = T62 | T61;
  assign T61 = 4'h1 == io_inner_grant_bits_g_type;
  assign T62 = 4'h0 == io_inner_grant_bits_g_type;
  assign T63 = T65 | T64;
  assign T64 = 4'h4 == io_inner_grant_bits_g_type;
  assign T65 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T66;
  assign T66 = T69 | T67;
  assign T67 = 3'h4 == xact_a_type;
  assign T68 = T56 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T69 = T71 | T70;
  assign T70 = 3'h3 == xact_a_type;
  assign T71 = 3'h2 == xact_a_type;
  assign T72 = T56 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T73 = T100 & T74;
  assign T74 = release_count == 1'h1;
  assign T367 = T368[1'h0:1'h0];
  assign T368 = reset ? 3'h0 : T75;
  assign T75 = T91 ? T374 : T76;
  assign T76 = T100 ? T373 : T77;
  assign T77 = T88 ? T78 : T369;
  assign T369 = {2'h0, release_count};
  assign T78 = T371 + T79;
  assign T79 = {1'h0, T80};
  assign T80 = T370 + T81;
  assign T81 = {1'h0, T82};
  assign T82 = mask_incoherent[2'h3:2'h3];
  assign T370 = {1'h0, T83};
  assign T83 = mask_incoherent[2'h2:2'h2];
  assign T371 = {1'h0, T84};
  assign T84 = T372 + T85;
  assign T85 = {1'h0, T86};
  assign T86 = mask_incoherent[1'h1:1'h1];
  assign T372 = {1'h0, T87};
  assign T87 = mask_incoherent[1'h0:1'h0];
  assign T88 = T56 & T47;
  assign T373 = {2'h0, T89};
  assign T89 = release_count - 1'h1;
  assign T374 = {2'h0, T90};
  assign T90 = release_count - 1'h1;
  assign T91 = T98 & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T95 | T94;
  assign T94 = 3'h2 == io_inner_release_bits_r_type;
  assign T95 = T97 | T96;
  assign T96 = 3'h1 == io_inner_release_bits_r_type;
  assign T97 = 3'h0 == io_inner_release_bits_r_type;
  assign T98 = T99 & io_inner_release_valid;
  assign T99 = 3'h1 == state;
  assign T100 = T110 & oacq_data_done;
  assign oacq_data_done = T108 ? T102 : T101;
  assign T101 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T102 = T107 & T103;
  assign T103 = R104 == 2'h3;
  assign T375 = reset ? 2'h0 : T105;
  assign T105 = T107 ? T106 : R104;
  assign T106 = R104 + 2'h1;
  assign T107 = T101 & T108;
  assign T108 = io_outer_acquire_bits_is_builtin_type & T109;
  assign T109 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T110 = T111 & io_outer_acquire_ready;
  assign T111 = T98 & T93;
  assign T112 = pending_outer_write ? 3'h3 : T113;
  assign T113 = pending_outer_read ? 3'h2 : 3'h4;
  assign T114 = T91 & T115;
  assign T115 = release_count == 1'h1;
  assign T116 = pending_outer_read ? 3'h2 : 3'h5;
  assign T117 = T118 & oacq_data_done;
  assign T118 = 3'h3 == state;
  assign T119 = T121 & T120;
  assign T120 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T121 = 3'h2 == state;
  assign T122 = T123 ? 3'h6 : 3'h0;
  assign T123 = T124 ^ 1'h1;
  assign T124 = io_inner_grant_bits_is_builtin_type & T125;
  assign T125 = io_inner_grant_bits_g_type == 4'h0;
  assign T126 = T139 & ignt_data_done;
  assign ignt_data_done = T134 ? T128 : T127;
  assign T127 = io_inner_grant_ready & io_inner_grant_valid;
  assign T128 = T133 & T129;
  assign T129 = R130 == 2'h3;
  assign T376 = reset ? 2'h0 : T131;
  assign T131 = T133 ? T132 : R130;
  assign T132 = R130 + 2'h1;
  assign T133 = T127 & T134;
  assign T134 = io_inner_grant_bits_is_builtin_type ? T138 : T135;
  assign T135 = T137 | T136;
  assign T136 = 4'h1 == io_inner_grant_bits_g_type;
  assign T137 = 4'h0 == io_inner_grant_bits_g_type;
  assign T138 = 4'h5 == io_inner_grant_bits_g_type;
  assign T139 = 3'h5 == state;
  assign T140 = T141 ? 3'h6 : 3'h0;
  assign T141 = T142 ^ 1'h1;
  assign T142 = io_inner_grant_bits_is_builtin_type & T143;
  assign T143 = io_inner_grant_bits_g_type == 4'h0;
  assign T144 = T145 & io_inner_grant_ready;
  assign T145 = 3'h4 == state;
  assign T146 = T147 & io_inner_finish_valid;
  assign T147 = 3'h6 == state;
  assign T149 = T150 | reset;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T154 & T152;
  assign T152 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T153 = T56 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T154 = T156 & T155;
  assign T155 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T156 = T171 & collect_iacq_data;
  assign T377 = reset ? 1'h0 : T157;
  assign T157 = T56 ? T169 : T158;
  assign T158 = T159 ? 1'h0 : collect_iacq_data;
  assign T159 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T167 ? T161 : T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T166 & T162;
  assign T162 = R163 == 2'h3;
  assign T378 = reset ? 2'h0 : T164;
  assign T164 = T166 ? T165 : R163;
  assign T165 = R163 + 2'h1;
  assign T166 = T160 & T167;
  assign T167 = io_inner_acquire_bits_is_builtin_type & T168;
  assign T168 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T169 = io_inner_acquire_bits_is_builtin_type & T170;
  assign T170 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T171 = state != 3'h0;
  assign T173 = T174 | reset;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T178 & T176;
  assign T176 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T177 = T56 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T178 = T180 & T179;
  assign T179 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T180 = T181 & collect_iacq_data;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T193 & T186;
  assign T186 = T188 | T187;
  assign T187 = 3'h5 == xact_a_type;
  assign T188 = T190 | T189;
  assign T189 = 3'h4 == xact_a_type;
  assign T190 = T192 | T191;
  assign T191 = 3'h2 == xact_a_type;
  assign T192 = 3'h0 == xact_a_type;
  assign T193 = T194 & xact_is_builtin_type;
  assign T194 = state != 3'h0;
  assign io_has_release_match = T195;
  assign T195 = T197 & T196;
  assign T196 = state == 3'h1;
  assign T197 = T199 & T198;
  assign T198 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T199 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T200 = T56 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T201;
  assign T201 = T202 & collect_iacq_data;
  assign T202 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T203;
  assign T203 = T205 & T204;
  assign T204 = collect_iacq_data ^ 1'h1;
  assign T205 = T207 & T206;
  assign T206 = state != 3'h0;
  assign T207 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T208;
  assign T208 = T139 ? io_inner_grant_ready : pending_ognt_ack;
  assign T379 = reset ? 1'h0 : T209;
  assign T209 = T117 ? 1'h1 : T210;
  assign T210 = T100 ? 1'h1 : T211;
  assign T211 = T212 ? 1'h0 : pending_ognt_ack;
  assign T212 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_union = T213;
  assign T213 = T121 ? outer_read_union : T214;
  assign T214 = T118 ? outer_write_acq_union : T215;
  assign T215 = T111 ? outer_write_rel_union : outer_read_union;
  assign outer_write_rel_union = T380;
  assign T380 = {8'h0, T216};
  assign T216 = {T217, 1'h1};
  assign T217 = 1'h1;
  assign outer_write_acq_union = T381;
  assign T381 = {8'h0, T218};
  assign T218 = {T219, 1'h1};
  assign T219 = 1'h1;
  assign outer_read_union = 10'h1c1;
  assign io_outer_acquire_bits_a_type = T220;
  assign T220 = T121 ? outer_read_a_type : T221;
  assign T221 = T118 ? outer_write_acq_a_type : T222;
  assign T222 = T111 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign outer_read_a_type = 3'h1;
  assign io_outer_acquire_bits_is_builtin_type = T223;
  assign T223 = T121 ? outer_read_is_builtin_type : T224;
  assign T224 = T118 ? outer_write_acq_is_builtin_type : T225;
  assign T225 = T111 ? outer_write_rel_is_builtin_type : outer_read_is_builtin_type;
  assign outer_write_rel_is_builtin_type = 1'h1;
  assign outer_write_acq_is_builtin_type = 1'h1;
  assign outer_read_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_data = T226;
  assign T226 = T121 ? outer_read_data : T227;
  assign T227 = T118 ? outer_write_acq_data : T228;
  assign T228 = T111 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_data;
  assign outer_write_acq_data = T229;
  assign T229 = T264 ? T250 : T230;
  assign T230 = T248 ? data_buffer_1 : data_buffer_0;
  assign T231 = T238 ? io_inner_acquire_bits_data : T232;
  assign T232 = T233 ? io_inner_acquire_bits_data : data_buffer_0;
  assign T233 = T237 & T234;
  assign T234 = T235[1'h0:1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = io_inner_acquire_bits_addr_beat;
  assign T237 = collect_iacq_data & io_inner_acquire_valid;
  assign T238 = T56 & T239;
  assign T239 = T240[1'h0:1'h0];
  assign T240 = 1'h1 << T241;
  assign T241 = 2'h0;
  assign T242 = T246 ? io_inner_acquire_bits_data : T243;
  assign T243 = T244 ? io_inner_acquire_bits_data : data_buffer_1;
  assign T244 = T237 & T245;
  assign T245 = T235[1'h1:1'h1];
  assign T246 = T56 & T247;
  assign T247 = T240[1'h1:1'h1];
  assign T248 = T249[1'h0:1'h0];
  assign T249 = oacq_data_cnt;
  assign oacq_data_cnt = T108 ? R104 : 2'h0;
  assign T250 = T263 ? data_buffer_3 : data_buffer_2;
  assign T251 = T255 ? io_inner_acquire_bits_data : T252;
  assign T252 = T253 ? io_inner_acquire_bits_data : data_buffer_2;
  assign T253 = T237 & T254;
  assign T254 = T235[2'h2:2'h2];
  assign T255 = T56 & T256;
  assign T256 = T240[2'h2:2'h2];
  assign T257 = T261 ? io_inner_acquire_bits_data : T258;
  assign T258 = T259 ? io_inner_acquire_bits_data : data_buffer_3;
  assign T259 = T237 & T260;
  assign T260 = T235[2'h3:2'h3];
  assign T261 = T56 & T262;
  assign T262 = T240[2'h3:2'h3];
  assign T263 = T249[1'h0:1'h0];
  assign T264 = T249[1'h1:1'h1];
  assign outer_read_data = 4'h0;
  assign io_outer_acquire_bits_addr_beat = T265;
  assign T265 = T121 ? outer_read_addr_beat : T266;
  assign T266 = T118 ? outer_write_acq_addr_beat : T267;
  assign T267 = T111 ? outer_write_rel_addr_beat : outer_read_addr_beat;
  assign outer_write_rel_addr_beat = io_inner_release_bits_addr_beat;
  assign outer_write_acq_addr_beat = oacq_data_cnt;
  assign outer_read_addr_beat = 2'h0;
  assign io_outer_acquire_bits_client_xact_id = T268;
  assign T268 = T121 ? outer_read_client_xact_id : T269;
  assign T269 = T118 ? outer_write_acq_client_xact_id : T270;
  assign T270 = T111 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h2;
  assign outer_write_acq_client_xact_id = 3'h2;
  assign outer_read_client_xact_id = 3'h2;
  assign io_outer_acquire_bits_addr_block = T271;
  assign T271 = T121 ? outer_read_addr_block : T272;
  assign T272 = T118 ? outer_write_acq_addr_block : T273;
  assign T273 = T111 ? outer_write_rel_addr_block : outer_read_addr_block;
  assign outer_write_rel_addr_block = xact_addr_block;
  assign outer_write_acq_addr_block = xact_addr_block;
  assign outer_read_addr_block = xact_addr_block;
  assign io_outer_acquire_valid = T274;
  assign T274 = T121 ? T301 : T275;
  assign T275 = T118 ? T276 : T111;
  assign T276 = T298 | T277;
  assign T277 = T282 & T278;
  assign T278 = T279 - 1'h1;
  assign T279 = 1'h1 << T280;
  assign T280 = T281 + 2'h1;
  assign T281 = oacq_data_cnt - oacq_data_cnt;
  assign T282 = iacq_data_valid >> oacq_data_cnt;
  assign T382 = reset ? 4'h0 : T283;
  assign T283 = T56 ? T291 : T284;
  assign T284 = T237 ? T285 : iacq_data_valid;
  assign T285 = T289 | T286;
  assign T286 = T383 & T287;
  assign T287 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T383 = T288 ? 4'hf : 4'h0;
  assign T288 = 1'h1;
  assign T289 = iacq_data_valid & T290;
  assign T290 = ~ T287;
  assign T291 = T292 << io_inner_acquire_bits_addr_beat;
  assign T292 = io_inner_acquire_bits_is_builtin_type & T293;
  assign T293 = T295 | T294;
  assign T294 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T295 = T297 | T296;
  assign T296 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T297 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T298 = T300 | T299;
  assign T299 = collect_iacq_data ^ 1'h1;
  assign T300 = pending_ognt_ack ^ 1'h1;
  assign T301 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T302;
  assign T302 = T99 ? T303 : 1'h0;
  assign T303 = T304 | io_outer_acquire_ready;
  assign T304 = T305 ^ 1'h1;
  assign T305 = T307 | T306;
  assign T306 = 3'h2 == io_inner_release_bits_r_type;
  assign T307 = T309 | T308;
  assign T308 = 3'h1 == io_inner_release_bits_r_type;
  assign T309 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T310;
  assign T310 = T384;
  assign T384 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T317;
  assign T317 = T318;
  assign T318 = xact_is_builtin_type ? T323 : T319;
  assign T319 = T322 ? 2'h1 : T320;
  assign T320 = T321 ? 2'h0 : 2'h2;
  assign T321 = xact_a_type == 3'h1;
  assign T322 = xact_a_type == 3'h0;
  assign T323 = T332 ? 2'h2 : T324;
  assign T324 = T331 ? 2'h0 : T325;
  assign T325 = T330 ? 2'h2 : T326;
  assign T326 = T329 ? 2'h0 : T327;
  assign T327 = T328 ? 2'h0 : 2'h2;
  assign T328 = xact_a_type == 3'h4;
  assign T329 = xact_a_type == 3'h2;
  assign T330 = xact_a_type == 3'h0;
  assign T331 = xact_a_type == 3'h3;
  assign T332 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T333;
  assign T333 = xact_addr_block;
  assign io_inner_probe_valid = T334;
  assign T334 = T99 ? T335 : 1'h0;
  assign T335 = pending_probes != 1'h0;
  assign T385 = T386[1'h0:1'h0];
  assign T386 = reset ? 4'h0 : T311;
  assign T311 = T316 ? T388 : T312;
  assign T312 = T88 ? mask_incoherent : T387;
  assign T387 = {3'h0, pending_probes};
  assign T388 = {2'h0, T313};
  assign T313 = T389 & T314;
  assign T314 = ~ T315;
  assign T315 = 1'h1 << 1'h0;
  assign T389 = {1'h0, pending_probes};
  assign T316 = T99 & io_inner_probe_ready;
  assign io_inner_finish_ready = T147;
  assign io_inner_grant_bits_client_id = T336;
  assign T336 = xact_client_id;
  assign io_inner_grant_bits_g_type = T337;
  assign T337 = T390;
  assign T390 = {1'h0, T338};
  assign T338 = xact_is_builtin_type ? T341 : T391;
  assign T391 = {1'h0, T339};
  assign T339 = T340 ? 2'h0 : 2'h1;
  assign T340 = xact_a_type == 3'h0;
  assign T341 = T352 ? 3'h4 : T342;
  assign T342 = T351 ? 3'h5 : T343;
  assign T343 = T350 ? 3'h3 : T344;
  assign T344 = T349 ? 3'h3 : T345;
  assign T345 = T348 ? 3'h4 : T346;
  assign T346 = T347 ? 3'h1 : 3'h3;
  assign T347 = xact_a_type == 3'h5;
  assign T348 = xact_a_type == 3'h4;
  assign T349 = xact_a_type == 3'h3;
  assign T350 = xact_a_type == 3'h2;
  assign T351 = xact_a_type == 3'h1;
  assign T352 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T353;
  assign T353 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T354;
  assign T354 = 3'h2;
  assign io_inner_grant_bits_client_xact_id = T355;
  assign T355 = xact_client_xact_id;
  assign io_inner_grant_bits_data = T356;
  assign T356 = 4'h0;
  assign io_inner_grant_bits_addr_beat = T357;
  assign T357 = 2'h0;
  assign io_inner_grant_valid = T358;
  assign T358 = T145 ? 1'h1 : T359;
  assign T359 = T139 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T360;
  assign T360 = T57 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics, subblock Gets/Puts, or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T172 <= 1'b1;
  if(!T173 && T172 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T148 <= 1'b1;
  if(!T149 && T148 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T146) begin
      state <= 3'h0;
    end else if(T144) begin
      state <= T140;
    end else if(T126) begin
      state <= T122;
    end else if(T119) begin
      state <= 3'h5;
    end else if(T117) begin
      state <= T116;
    end else if(T114) begin
      state <= T112;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T16;
    end
    if(T56) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T56) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T367;
    if(reset) begin
      R104 <= 2'h0;
    end else if(T107) begin
      R104 <= T106;
    end
    if(reset) begin
      R130 <= 2'h0;
    end else if(T133) begin
      R130 <= T132;
    end
    if(T56) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T56) begin
      collect_iacq_data <= T169;
    end else if(T159) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R163 <= 2'h0;
    end else if(T166) begin
      R163 <= T165;
    end
    if(T56) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T56) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T117) begin
      pending_ognt_ack <= 1'h1;
    end else if(T100) begin
      pending_ognt_ack <= 1'h1;
    end else if(T212) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T238) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T233) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T246) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T244) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T255) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T253) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T261) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T259) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T56) begin
      iacq_data_valid <= T291;
    end else if(T237) begin
      iacq_data_valid <= T285;
    end
    pending_probes <= T385;
  end
endmodule

module BroadcastAcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [3:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [9:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [3:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[9:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [2:0] state;
  wire[2:0] T361;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire pending_outer_read_;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T362;
  wire[2:0] T22;
  wire[2:0] T363;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire pending_outer_write_;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[3:0] mask_incoherent;
  wire[3:0] T364;
  wire T48;
  wire T49;
  wire[3:0] mask_self;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T365;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T366;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire pending_outer_read;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire pending_outer_write;
  wire T66;
  wire T67;
  reg [2:0] xact_a_type;
  wire[2:0] T68;
  wire T69;
  wire T70;
  wire T71;
  reg  xact_is_builtin_type;
  wire T72;
  wire T73;
  wire T74;
  reg  release_count;
  wire T367;
  wire[2:0] T368;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T369;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T370;
  wire T83;
  wire[2:0] T371;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T372;
  wire T87;
  wire T88;
  wire[2:0] T373;
  wire T89;
  wire[2:0] T374;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire oacq_data_done;
  wire T101;
  wire T102;
  wire T103;
  reg [1:0] R104;
  wire[1:0] T375;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire ignt_data_done;
  wire T127;
  wire T128;
  wire T129;
  reg [1:0] R130;
  wire[1:0] T376;
  wire[1:0] T131;
  wire[1:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[2:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  reg[0:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  xact_client_xact_id;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  reg  collect_iacq_data;
  wire T377;
  wire T157;
  wire T158;
  wire T159;
  wire iacq_data_done;
  wire T160;
  wire T161;
  wire T162;
  reg [1:0] R163;
  wire[1:0] T378;
  wire[1:0] T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  reg[0:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg [1:0] xact_client_id;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg [25:0] xact_addr_block;
  wire[25:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg  pending_ognt_ack;
  wire T379;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[9:0] T213;
  wire[9:0] T214;
  wire[9:0] T215;
  wire[9:0] outer_write_rel_union;
  wire[9:0] T380;
  wire[1:0] T216;
  wire T217;
  wire[9:0] outer_write_acq_union;
  wire[9:0] T381;
  wire[1:0] T218;
  wire T219;
  wire[9:0] outer_read_union;
  wire[2:0] T220;
  wire[2:0] T221;
  wire[2:0] T222;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[2:0] outer_read_a_type;
  wire T223;
  wire T224;
  wire T225;
  wire outer_write_rel_is_builtin_type;
  wire outer_write_acq_is_builtin_type;
  wire outer_read_is_builtin_type;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T229;
  wire[3:0] T230;
  reg [3:0] data_buffer_0;
  wire[3:0] T231;
  wire[3:0] T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire[3:0] T240;
  wire[1:0] T241;
  reg [3:0] data_buffer_1;
  wire[3:0] T242;
  wire[3:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T250;
  reg [3:0] data_buffer_2;
  wire[3:0] T251;
  wire[3:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  reg [3:0] data_buffer_3;
  wire[3:0] T257;
  wire[3:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] outer_read_data;
  wire[1:0] T265;
  wire[1:0] T266;
  wire[1:0] T267;
  wire[1:0] outer_write_rel_addr_beat;
  wire[1:0] outer_write_acq_addr_beat;
  wire[1:0] outer_read_addr_beat;
  wire[2:0] T268;
  wire[2:0] T269;
  wire[2:0] T270;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[25:0] T271;
  wire[25:0] T272;
  wire[25:0] T273;
  wire[25:0] outer_write_rel_addr_block;
  wire[25:0] outer_write_acq_addr_block;
  wire[25:0] outer_read_addr_block;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[1:0] T280;
  wire[1:0] T281;
  wire T282;
  reg [3:0] iacq_data_valid;
  wire[3:0] T382;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[3:0] T286;
  wire[3:0] T287;
  wire[3:0] T383;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire[1:0] T310;
  wire[1:0] T384;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire[25:0] T333;
  wire T334;
  wire T335;
  reg  pending_probes;
  wire T385;
  wire[3:0] T386;
  wire[3:0] T311;
  wire[3:0] T312;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire[1:0] T389;
  wire T316;
  wire[1:0] T336;
  wire[3:0] T337;
  wire[3:0] T390;
  wire[2:0] T338;
  wire[2:0] T391;
  wire[1:0] T339;
  wire T340;
  wire[2:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[2:0] T354;
  wire T355;
  wire[3:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R104 = {1{$random}};
    R130 = {1{$random}};
    T148 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R163 = {1{$random}};
    T172 = 1'b0;
    xact_client_id = {1{$random}};
    T182 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    data_buffer_0 = {1{$random}};
    data_buffer_1 = {1{$random}};
    data_buffer_2 = {1{$random}};
    data_buffer_3 = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T7 & T6;
  assign T6 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T7 = state == 3'h0;
  assign T361 = reset ? 3'h0 : T8;
  assign T8 = T146 ? 3'h0 : T9;
  assign T9 = T144 ? T140 : T10;
  assign T10 = T126 ? T122 : T11;
  assign T11 = T119 ? 3'h5 : T12;
  assign T12 = T117 ? T116 : T13;
  assign T13 = T114 ? T112 : T14;
  assign T14 = T73 ? T58 : T15;
  assign T15 = T56 ? T16 : state;
  assign T16 = T47 ? 3'h1 : T17;
  assign T17 = pending_outer_write_ ? 3'h3 : T18;
  assign T18 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T41 ? T38 : T19;
  assign T19 = T37 | T20;
  assign T20 = 4'h1 == T21;
  assign T21 = T362;
  assign T362 = {1'h0, T22};
  assign T22 = io_inner_acquire_bits_is_builtin_type ? T25 : T363;
  assign T363 = {1'h0, T23};
  assign T23 = T24 ? 2'h0 : 2'h1;
  assign T24 = io_inner_acquire_bits_a_type == 3'h0;
  assign T25 = T36 ? 3'h4 : T26;
  assign T26 = T35 ? 3'h5 : T27;
  assign T27 = T34 ? 3'h3 : T28;
  assign T28 = T33 ? 3'h3 : T29;
  assign T29 = T32 ? 3'h4 : T30;
  assign T30 = T31 ? 3'h1 : 3'h3;
  assign T31 = io_inner_acquire_bits_a_type == 3'h5;
  assign T32 = io_inner_acquire_bits_a_type == 3'h4;
  assign T33 = io_inner_acquire_bits_a_type == 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h2;
  assign T35 = io_inner_acquire_bits_a_type == 3'h1;
  assign T36 = io_inner_acquire_bits_a_type == 3'h0;
  assign T37 = 4'h0 == T21;
  assign T38 = T40 | T39;
  assign T39 = 4'h4 == T21;
  assign T40 = 4'h5 == T21;
  assign T41 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T42;
  assign T42 = T44 | T43;
  assign T43 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T46 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T47 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T364;
  assign T364 = {3'h0, T48};
  assign T48 = ~ T49;
  assign T49 = io_incoherent_0;
  assign mask_self = T53 | T50;
  assign T50 = T365 & T51;
  assign T51 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T365 = T52 ? 4'hf : 4'h0;
  assign T52 = 1'h0;
  assign T53 = T366 & T54;
  assign T54 = ~ T51;
  assign T366 = {3'h0, T55};
  assign T55 = 1'h1;
  assign T56 = T57 & io_inner_acquire_valid;
  assign T57 = 3'h0 == state;
  assign T58 = pending_outer_write ? 3'h3 : T59;
  assign T59 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T63 : T60;
  assign T60 = T62 | T61;
  assign T61 = 4'h1 == io_inner_grant_bits_g_type;
  assign T62 = 4'h0 == io_inner_grant_bits_g_type;
  assign T63 = T65 | T64;
  assign T64 = 4'h4 == io_inner_grant_bits_g_type;
  assign T65 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T66;
  assign T66 = T69 | T67;
  assign T67 = 3'h4 == xact_a_type;
  assign T68 = T56 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T69 = T71 | T70;
  assign T70 = 3'h3 == xact_a_type;
  assign T71 = 3'h2 == xact_a_type;
  assign T72 = T56 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T73 = T100 & T74;
  assign T74 = release_count == 1'h1;
  assign T367 = T368[1'h0:1'h0];
  assign T368 = reset ? 3'h0 : T75;
  assign T75 = T91 ? T374 : T76;
  assign T76 = T100 ? T373 : T77;
  assign T77 = T88 ? T78 : T369;
  assign T369 = {2'h0, release_count};
  assign T78 = T371 + T79;
  assign T79 = {1'h0, T80};
  assign T80 = T370 + T81;
  assign T81 = {1'h0, T82};
  assign T82 = mask_incoherent[2'h3:2'h3];
  assign T370 = {1'h0, T83};
  assign T83 = mask_incoherent[2'h2:2'h2];
  assign T371 = {1'h0, T84};
  assign T84 = T372 + T85;
  assign T85 = {1'h0, T86};
  assign T86 = mask_incoherent[1'h1:1'h1];
  assign T372 = {1'h0, T87};
  assign T87 = mask_incoherent[1'h0:1'h0];
  assign T88 = T56 & T47;
  assign T373 = {2'h0, T89};
  assign T89 = release_count - 1'h1;
  assign T374 = {2'h0, T90};
  assign T90 = release_count - 1'h1;
  assign T91 = T98 & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T95 | T94;
  assign T94 = 3'h2 == io_inner_release_bits_r_type;
  assign T95 = T97 | T96;
  assign T96 = 3'h1 == io_inner_release_bits_r_type;
  assign T97 = 3'h0 == io_inner_release_bits_r_type;
  assign T98 = T99 & io_inner_release_valid;
  assign T99 = 3'h1 == state;
  assign T100 = T110 & oacq_data_done;
  assign oacq_data_done = T108 ? T102 : T101;
  assign T101 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T102 = T107 & T103;
  assign T103 = R104 == 2'h3;
  assign T375 = reset ? 2'h0 : T105;
  assign T105 = T107 ? T106 : R104;
  assign T106 = R104 + 2'h1;
  assign T107 = T101 & T108;
  assign T108 = io_outer_acquire_bits_is_builtin_type & T109;
  assign T109 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T110 = T111 & io_outer_acquire_ready;
  assign T111 = T98 & T93;
  assign T112 = pending_outer_write ? 3'h3 : T113;
  assign T113 = pending_outer_read ? 3'h2 : 3'h4;
  assign T114 = T91 & T115;
  assign T115 = release_count == 1'h1;
  assign T116 = pending_outer_read ? 3'h2 : 3'h5;
  assign T117 = T118 & oacq_data_done;
  assign T118 = 3'h3 == state;
  assign T119 = T121 & T120;
  assign T120 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T121 = 3'h2 == state;
  assign T122 = T123 ? 3'h6 : 3'h0;
  assign T123 = T124 ^ 1'h1;
  assign T124 = io_inner_grant_bits_is_builtin_type & T125;
  assign T125 = io_inner_grant_bits_g_type == 4'h0;
  assign T126 = T139 & ignt_data_done;
  assign ignt_data_done = T134 ? T128 : T127;
  assign T127 = io_inner_grant_ready & io_inner_grant_valid;
  assign T128 = T133 & T129;
  assign T129 = R130 == 2'h3;
  assign T376 = reset ? 2'h0 : T131;
  assign T131 = T133 ? T132 : R130;
  assign T132 = R130 + 2'h1;
  assign T133 = T127 & T134;
  assign T134 = io_inner_grant_bits_is_builtin_type ? T138 : T135;
  assign T135 = T137 | T136;
  assign T136 = 4'h1 == io_inner_grant_bits_g_type;
  assign T137 = 4'h0 == io_inner_grant_bits_g_type;
  assign T138 = 4'h5 == io_inner_grant_bits_g_type;
  assign T139 = 3'h5 == state;
  assign T140 = T141 ? 3'h6 : 3'h0;
  assign T141 = T142 ^ 1'h1;
  assign T142 = io_inner_grant_bits_is_builtin_type & T143;
  assign T143 = io_inner_grant_bits_g_type == 4'h0;
  assign T144 = T145 & io_inner_grant_ready;
  assign T145 = 3'h4 == state;
  assign T146 = T147 & io_inner_finish_valid;
  assign T147 = 3'h6 == state;
  assign T149 = T150 | reset;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T154 & T152;
  assign T152 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T153 = T56 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T154 = T156 & T155;
  assign T155 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T156 = T171 & collect_iacq_data;
  assign T377 = reset ? 1'h0 : T157;
  assign T157 = T56 ? T169 : T158;
  assign T158 = T159 ? 1'h0 : collect_iacq_data;
  assign T159 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T167 ? T161 : T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T166 & T162;
  assign T162 = R163 == 2'h3;
  assign T378 = reset ? 2'h0 : T164;
  assign T164 = T166 ? T165 : R163;
  assign T165 = R163 + 2'h1;
  assign T166 = T160 & T167;
  assign T167 = io_inner_acquire_bits_is_builtin_type & T168;
  assign T168 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T169 = io_inner_acquire_bits_is_builtin_type & T170;
  assign T170 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T171 = state != 3'h0;
  assign T173 = T174 | reset;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T178 & T176;
  assign T176 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T177 = T56 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T178 = T180 & T179;
  assign T179 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T180 = T181 & collect_iacq_data;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T193 & T186;
  assign T186 = T188 | T187;
  assign T187 = 3'h5 == xact_a_type;
  assign T188 = T190 | T189;
  assign T189 = 3'h4 == xact_a_type;
  assign T190 = T192 | T191;
  assign T191 = 3'h2 == xact_a_type;
  assign T192 = 3'h0 == xact_a_type;
  assign T193 = T194 & xact_is_builtin_type;
  assign T194 = state != 3'h0;
  assign io_has_release_match = T195;
  assign T195 = T197 & T196;
  assign T196 = state == 3'h1;
  assign T197 = T199 & T198;
  assign T198 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T199 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T200 = T56 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T201;
  assign T201 = T202 & collect_iacq_data;
  assign T202 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T203;
  assign T203 = T205 & T204;
  assign T204 = collect_iacq_data ^ 1'h1;
  assign T205 = T207 & T206;
  assign T206 = state != 3'h0;
  assign T207 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T208;
  assign T208 = T139 ? io_inner_grant_ready : pending_ognt_ack;
  assign T379 = reset ? 1'h0 : T209;
  assign T209 = T117 ? 1'h1 : T210;
  assign T210 = T100 ? 1'h1 : T211;
  assign T211 = T212 ? 1'h0 : pending_ognt_ack;
  assign T212 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_union = T213;
  assign T213 = T121 ? outer_read_union : T214;
  assign T214 = T118 ? outer_write_acq_union : T215;
  assign T215 = T111 ? outer_write_rel_union : outer_read_union;
  assign outer_write_rel_union = T380;
  assign T380 = {8'h0, T216};
  assign T216 = {T217, 1'h1};
  assign T217 = 1'h1;
  assign outer_write_acq_union = T381;
  assign T381 = {8'h0, T218};
  assign T218 = {T219, 1'h1};
  assign T219 = 1'h1;
  assign outer_read_union = 10'h1c1;
  assign io_outer_acquire_bits_a_type = T220;
  assign T220 = T121 ? outer_read_a_type : T221;
  assign T221 = T118 ? outer_write_acq_a_type : T222;
  assign T222 = T111 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign outer_read_a_type = 3'h1;
  assign io_outer_acquire_bits_is_builtin_type = T223;
  assign T223 = T121 ? outer_read_is_builtin_type : T224;
  assign T224 = T118 ? outer_write_acq_is_builtin_type : T225;
  assign T225 = T111 ? outer_write_rel_is_builtin_type : outer_read_is_builtin_type;
  assign outer_write_rel_is_builtin_type = 1'h1;
  assign outer_write_acq_is_builtin_type = 1'h1;
  assign outer_read_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_data = T226;
  assign T226 = T121 ? outer_read_data : T227;
  assign T227 = T118 ? outer_write_acq_data : T228;
  assign T228 = T111 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_data;
  assign outer_write_acq_data = T229;
  assign T229 = T264 ? T250 : T230;
  assign T230 = T248 ? data_buffer_1 : data_buffer_0;
  assign T231 = T238 ? io_inner_acquire_bits_data : T232;
  assign T232 = T233 ? io_inner_acquire_bits_data : data_buffer_0;
  assign T233 = T237 & T234;
  assign T234 = T235[1'h0:1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = io_inner_acquire_bits_addr_beat;
  assign T237 = collect_iacq_data & io_inner_acquire_valid;
  assign T238 = T56 & T239;
  assign T239 = T240[1'h0:1'h0];
  assign T240 = 1'h1 << T241;
  assign T241 = 2'h0;
  assign T242 = T246 ? io_inner_acquire_bits_data : T243;
  assign T243 = T244 ? io_inner_acquire_bits_data : data_buffer_1;
  assign T244 = T237 & T245;
  assign T245 = T235[1'h1:1'h1];
  assign T246 = T56 & T247;
  assign T247 = T240[1'h1:1'h1];
  assign T248 = T249[1'h0:1'h0];
  assign T249 = oacq_data_cnt;
  assign oacq_data_cnt = T108 ? R104 : 2'h0;
  assign T250 = T263 ? data_buffer_3 : data_buffer_2;
  assign T251 = T255 ? io_inner_acquire_bits_data : T252;
  assign T252 = T253 ? io_inner_acquire_bits_data : data_buffer_2;
  assign T253 = T237 & T254;
  assign T254 = T235[2'h2:2'h2];
  assign T255 = T56 & T256;
  assign T256 = T240[2'h2:2'h2];
  assign T257 = T261 ? io_inner_acquire_bits_data : T258;
  assign T258 = T259 ? io_inner_acquire_bits_data : data_buffer_3;
  assign T259 = T237 & T260;
  assign T260 = T235[2'h3:2'h3];
  assign T261 = T56 & T262;
  assign T262 = T240[2'h3:2'h3];
  assign T263 = T249[1'h0:1'h0];
  assign T264 = T249[1'h1:1'h1];
  assign outer_read_data = 4'h0;
  assign io_outer_acquire_bits_addr_beat = T265;
  assign T265 = T121 ? outer_read_addr_beat : T266;
  assign T266 = T118 ? outer_write_acq_addr_beat : T267;
  assign T267 = T111 ? outer_write_rel_addr_beat : outer_read_addr_beat;
  assign outer_write_rel_addr_beat = io_inner_release_bits_addr_beat;
  assign outer_write_acq_addr_beat = oacq_data_cnt;
  assign outer_read_addr_beat = 2'h0;
  assign io_outer_acquire_bits_client_xact_id = T268;
  assign T268 = T121 ? outer_read_client_xact_id : T269;
  assign T269 = T118 ? outer_write_acq_client_xact_id : T270;
  assign T270 = T111 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h3;
  assign outer_write_acq_client_xact_id = 3'h3;
  assign outer_read_client_xact_id = 3'h3;
  assign io_outer_acquire_bits_addr_block = T271;
  assign T271 = T121 ? outer_read_addr_block : T272;
  assign T272 = T118 ? outer_write_acq_addr_block : T273;
  assign T273 = T111 ? outer_write_rel_addr_block : outer_read_addr_block;
  assign outer_write_rel_addr_block = xact_addr_block;
  assign outer_write_acq_addr_block = xact_addr_block;
  assign outer_read_addr_block = xact_addr_block;
  assign io_outer_acquire_valid = T274;
  assign T274 = T121 ? T301 : T275;
  assign T275 = T118 ? T276 : T111;
  assign T276 = T298 | T277;
  assign T277 = T282 & T278;
  assign T278 = T279 - 1'h1;
  assign T279 = 1'h1 << T280;
  assign T280 = T281 + 2'h1;
  assign T281 = oacq_data_cnt - oacq_data_cnt;
  assign T282 = iacq_data_valid >> oacq_data_cnt;
  assign T382 = reset ? 4'h0 : T283;
  assign T283 = T56 ? T291 : T284;
  assign T284 = T237 ? T285 : iacq_data_valid;
  assign T285 = T289 | T286;
  assign T286 = T383 & T287;
  assign T287 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T383 = T288 ? 4'hf : 4'h0;
  assign T288 = 1'h1;
  assign T289 = iacq_data_valid & T290;
  assign T290 = ~ T287;
  assign T291 = T292 << io_inner_acquire_bits_addr_beat;
  assign T292 = io_inner_acquire_bits_is_builtin_type & T293;
  assign T293 = T295 | T294;
  assign T294 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T295 = T297 | T296;
  assign T296 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T297 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T298 = T300 | T299;
  assign T299 = collect_iacq_data ^ 1'h1;
  assign T300 = pending_ognt_ack ^ 1'h1;
  assign T301 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T302;
  assign T302 = T99 ? T303 : 1'h0;
  assign T303 = T304 | io_outer_acquire_ready;
  assign T304 = T305 ^ 1'h1;
  assign T305 = T307 | T306;
  assign T306 = 3'h2 == io_inner_release_bits_r_type;
  assign T307 = T309 | T308;
  assign T308 = 3'h1 == io_inner_release_bits_r_type;
  assign T309 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T310;
  assign T310 = T384;
  assign T384 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T317;
  assign T317 = T318;
  assign T318 = xact_is_builtin_type ? T323 : T319;
  assign T319 = T322 ? 2'h1 : T320;
  assign T320 = T321 ? 2'h0 : 2'h2;
  assign T321 = xact_a_type == 3'h1;
  assign T322 = xact_a_type == 3'h0;
  assign T323 = T332 ? 2'h2 : T324;
  assign T324 = T331 ? 2'h0 : T325;
  assign T325 = T330 ? 2'h2 : T326;
  assign T326 = T329 ? 2'h0 : T327;
  assign T327 = T328 ? 2'h0 : 2'h2;
  assign T328 = xact_a_type == 3'h4;
  assign T329 = xact_a_type == 3'h2;
  assign T330 = xact_a_type == 3'h0;
  assign T331 = xact_a_type == 3'h3;
  assign T332 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T333;
  assign T333 = xact_addr_block;
  assign io_inner_probe_valid = T334;
  assign T334 = T99 ? T335 : 1'h0;
  assign T335 = pending_probes != 1'h0;
  assign T385 = T386[1'h0:1'h0];
  assign T386 = reset ? 4'h0 : T311;
  assign T311 = T316 ? T388 : T312;
  assign T312 = T88 ? mask_incoherent : T387;
  assign T387 = {3'h0, pending_probes};
  assign T388 = {2'h0, T313};
  assign T313 = T389 & T314;
  assign T314 = ~ T315;
  assign T315 = 1'h1 << 1'h0;
  assign T389 = {1'h0, pending_probes};
  assign T316 = T99 & io_inner_probe_ready;
  assign io_inner_finish_ready = T147;
  assign io_inner_grant_bits_client_id = T336;
  assign T336 = xact_client_id;
  assign io_inner_grant_bits_g_type = T337;
  assign T337 = T390;
  assign T390 = {1'h0, T338};
  assign T338 = xact_is_builtin_type ? T341 : T391;
  assign T391 = {1'h0, T339};
  assign T339 = T340 ? 2'h0 : 2'h1;
  assign T340 = xact_a_type == 3'h0;
  assign T341 = T352 ? 3'h4 : T342;
  assign T342 = T351 ? 3'h5 : T343;
  assign T343 = T350 ? 3'h3 : T344;
  assign T344 = T349 ? 3'h3 : T345;
  assign T345 = T348 ? 3'h4 : T346;
  assign T346 = T347 ? 3'h1 : 3'h3;
  assign T347 = xact_a_type == 3'h5;
  assign T348 = xact_a_type == 3'h4;
  assign T349 = xact_a_type == 3'h3;
  assign T350 = xact_a_type == 3'h2;
  assign T351 = xact_a_type == 3'h1;
  assign T352 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T353;
  assign T353 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T354;
  assign T354 = 3'h3;
  assign io_inner_grant_bits_client_xact_id = T355;
  assign T355 = xact_client_xact_id;
  assign io_inner_grant_bits_data = T356;
  assign T356 = 4'h0;
  assign io_inner_grant_bits_addr_beat = T357;
  assign T357 = 2'h0;
  assign io_inner_grant_valid = T358;
  assign T358 = T145 ? 1'h1 : T359;
  assign T359 = T139 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T360;
  assign T360 = T57 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics, subblock Gets/Puts, or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T172 <= 1'b1;
  if(!T173 && T172 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T148 <= 1'b1;
  if(!T149 && T148 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T146) begin
      state <= 3'h0;
    end else if(T144) begin
      state <= T140;
    end else if(T126) begin
      state <= T122;
    end else if(T119) begin
      state <= 3'h5;
    end else if(T117) begin
      state <= T116;
    end else if(T114) begin
      state <= T112;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T16;
    end
    if(T56) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T56) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T367;
    if(reset) begin
      R104 <= 2'h0;
    end else if(T107) begin
      R104 <= T106;
    end
    if(reset) begin
      R130 <= 2'h0;
    end else if(T133) begin
      R130 <= T132;
    end
    if(T56) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T56) begin
      collect_iacq_data <= T169;
    end else if(T159) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R163 <= 2'h0;
    end else if(T166) begin
      R163 <= T165;
    end
    if(T56) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T56) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T117) begin
      pending_ognt_ack <= 1'h1;
    end else if(T100) begin
      pending_ognt_ack <= 1'h1;
    end else if(T212) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T238) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T233) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T246) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T244) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T255) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T253) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T261) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T259) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T56) begin
      iacq_data_valid <= T291;
    end else if(T237) begin
      iacq_data_valid <= T285;
    end
    pending_probes <= T385;
  end
endmodule

module BroadcastAcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [3:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [9:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[3:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [3:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[9:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [3:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg [2:0] state;
  wire[2:0] T361;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire pending_outer_read_;
  wire T19;
  wire T20;
  wire[3:0] T21;
  wire[3:0] T362;
  wire[2:0] T22;
  wire[2:0] T363;
  wire[1:0] T23;
  wire T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire pending_outer_write_;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[3:0] mask_incoherent;
  wire[3:0] T364;
  wire T48;
  wire T49;
  wire[3:0] mask_self;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T365;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T366;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire pending_outer_read;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire pending_outer_write;
  wire T66;
  wire T67;
  reg [2:0] xact_a_type;
  wire[2:0] T68;
  wire T69;
  wire T70;
  wire T71;
  reg  xact_is_builtin_type;
  wire T72;
  wire T73;
  wire T74;
  reg  release_count;
  wire T367;
  wire[2:0] T368;
  wire[2:0] T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T369;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T370;
  wire T83;
  wire[2:0] T371;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[1:0] T372;
  wire T87;
  wire T88;
  wire[2:0] T373;
  wire T89;
  wire[2:0] T374;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire oacq_data_done;
  wire T101;
  wire T102;
  wire T103;
  reg [1:0] R104;
  wire[1:0] T375;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[2:0] T112;
  wire[2:0] T113;
  wire T114;
  wire T115;
  wire[2:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire ignt_data_done;
  wire T127;
  wire T128;
  wire T129;
  reg [1:0] R130;
  wire[1:0] T376;
  wire[1:0] T131;
  wire[1:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[2:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  reg[0:0] T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg  xact_client_xact_id;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  reg  collect_iacq_data;
  wire T377;
  wire T157;
  wire T158;
  wire T159;
  wire iacq_data_done;
  wire T160;
  wire T161;
  wire T162;
  reg [1:0] R163;
  wire[1:0] T378;
  wire[1:0] T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  reg[0:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg [1:0] xact_client_id;
  wire[1:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg[0:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg [25:0] xact_addr_block;
  wire[25:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg  pending_ognt_ack;
  wire T379;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[9:0] T213;
  wire[9:0] T214;
  wire[9:0] T215;
  wire[9:0] outer_write_rel_union;
  wire[9:0] T380;
  wire[1:0] T216;
  wire T217;
  wire[9:0] outer_write_acq_union;
  wire[9:0] T381;
  wire[1:0] T218;
  wire T219;
  wire[9:0] outer_read_union;
  wire[2:0] T220;
  wire[2:0] T221;
  wire[2:0] T222;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[2:0] outer_read_a_type;
  wire T223;
  wire T224;
  wire T225;
  wire outer_write_rel_is_builtin_type;
  wire outer_write_acq_is_builtin_type;
  wire outer_read_is_builtin_type;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] outer_write_rel_data;
  wire[3:0] outer_write_acq_data;
  wire[3:0] T229;
  wire[3:0] T230;
  reg [3:0] data_buffer_0;
  wire[3:0] T231;
  wire[3:0] T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[1:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire[3:0] T240;
  wire[1:0] T241;
  reg [3:0] data_buffer_1;
  wire[3:0] T242;
  wire[3:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T250;
  reg [3:0] data_buffer_2;
  wire[3:0] T251;
  wire[3:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  reg [3:0] data_buffer_3;
  wire[3:0] T257;
  wire[3:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] outer_read_data;
  wire[1:0] T265;
  wire[1:0] T266;
  wire[1:0] T267;
  wire[1:0] outer_write_rel_addr_beat;
  wire[1:0] outer_write_acq_addr_beat;
  wire[1:0] outer_read_addr_beat;
  wire[2:0] T268;
  wire[2:0] T269;
  wire[2:0] T270;
  wire[2:0] outer_write_rel_client_xact_id;
  wire[2:0] outer_write_acq_client_xact_id;
  wire[2:0] outer_read_client_xact_id;
  wire[25:0] T271;
  wire[25:0] T272;
  wire[25:0] T273;
  wire[25:0] outer_write_rel_addr_block;
  wire[25:0] outer_write_acq_addr_block;
  wire[25:0] outer_read_addr_block;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[1:0] T280;
  wire[1:0] T281;
  wire T282;
  reg [3:0] iacq_data_valid;
  wire[3:0] T382;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[3:0] T286;
  wire[3:0] T287;
  wire[3:0] T383;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire[1:0] T310;
  wire[1:0] T384;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire[25:0] T333;
  wire T334;
  wire T335;
  reg  pending_probes;
  wire T385;
  wire[3:0] T386;
  wire[3:0] T311;
  wire[3:0] T312;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire[1:0] T389;
  wire T316;
  wire[1:0] T336;
  wire[3:0] T337;
  wire[3:0] T390;
  wire[2:0] T338;
  wire[2:0] T391;
  wire[1:0] T339;
  wire T340;
  wire[2:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire[2:0] T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire[2:0] T354;
  wire T355;
  wire[3:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R104 = {1{$random}};
    R130 = {1{$random}};
    T148 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R163 = {1{$random}};
    T172 = 1'b0;
    xact_client_id = {1{$random}};
    T182 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    data_buffer_0 = {1{$random}};
    data_buffer_1 = {1{$random}};
    data_buffer_2 = {1{$random}};
    data_buffer_3 = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T7 & T6;
  assign T6 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T7 = state == 3'h0;
  assign T361 = reset ? 3'h0 : T8;
  assign T8 = T146 ? 3'h0 : T9;
  assign T9 = T144 ? T140 : T10;
  assign T10 = T126 ? T122 : T11;
  assign T11 = T119 ? 3'h5 : T12;
  assign T12 = T117 ? T116 : T13;
  assign T13 = T114 ? T112 : T14;
  assign T14 = T73 ? T58 : T15;
  assign T15 = T56 ? T16 : state;
  assign T16 = T47 ? 3'h1 : T17;
  assign T17 = pending_outer_write_ ? 3'h3 : T18;
  assign T18 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T41 ? T38 : T19;
  assign T19 = T37 | T20;
  assign T20 = 4'h1 == T21;
  assign T21 = T362;
  assign T362 = {1'h0, T22};
  assign T22 = io_inner_acquire_bits_is_builtin_type ? T25 : T363;
  assign T363 = {1'h0, T23};
  assign T23 = T24 ? 2'h0 : 2'h1;
  assign T24 = io_inner_acquire_bits_a_type == 3'h0;
  assign T25 = T36 ? 3'h4 : T26;
  assign T26 = T35 ? 3'h5 : T27;
  assign T27 = T34 ? 3'h3 : T28;
  assign T28 = T33 ? 3'h3 : T29;
  assign T29 = T32 ? 3'h4 : T30;
  assign T30 = T31 ? 3'h1 : 3'h3;
  assign T31 = io_inner_acquire_bits_a_type == 3'h5;
  assign T32 = io_inner_acquire_bits_a_type == 3'h4;
  assign T33 = io_inner_acquire_bits_a_type == 3'h3;
  assign T34 = io_inner_acquire_bits_a_type == 3'h2;
  assign T35 = io_inner_acquire_bits_a_type == 3'h1;
  assign T36 = io_inner_acquire_bits_a_type == 3'h0;
  assign T37 = 4'h0 == T21;
  assign T38 = T40 | T39;
  assign T39 = 4'h4 == T21;
  assign T40 = 4'h5 == T21;
  assign T41 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T42;
  assign T42 = T44 | T43;
  assign T43 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T46 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T47 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T364;
  assign T364 = {3'h0, T48};
  assign T48 = ~ T49;
  assign T49 = io_incoherent_0;
  assign mask_self = T53 | T50;
  assign T50 = T365 & T51;
  assign T51 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T365 = T52 ? 4'hf : 4'h0;
  assign T52 = 1'h0;
  assign T53 = T366 & T54;
  assign T54 = ~ T51;
  assign T366 = {3'h0, T55};
  assign T55 = 1'h1;
  assign T56 = T57 & io_inner_acquire_valid;
  assign T57 = 3'h0 == state;
  assign T58 = pending_outer_write ? 3'h3 : T59;
  assign T59 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T63 : T60;
  assign T60 = T62 | T61;
  assign T61 = 4'h1 == io_inner_grant_bits_g_type;
  assign T62 = 4'h0 == io_inner_grant_bits_g_type;
  assign T63 = T65 | T64;
  assign T64 = 4'h4 == io_inner_grant_bits_g_type;
  assign T65 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T66;
  assign T66 = T69 | T67;
  assign T67 = 3'h4 == xact_a_type;
  assign T68 = T56 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T69 = T71 | T70;
  assign T70 = 3'h3 == xact_a_type;
  assign T71 = 3'h2 == xact_a_type;
  assign T72 = T56 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T73 = T100 & T74;
  assign T74 = release_count == 1'h1;
  assign T367 = T368[1'h0:1'h0];
  assign T368 = reset ? 3'h0 : T75;
  assign T75 = T91 ? T374 : T76;
  assign T76 = T100 ? T373 : T77;
  assign T77 = T88 ? T78 : T369;
  assign T369 = {2'h0, release_count};
  assign T78 = T371 + T79;
  assign T79 = {1'h0, T80};
  assign T80 = T370 + T81;
  assign T81 = {1'h0, T82};
  assign T82 = mask_incoherent[2'h3:2'h3];
  assign T370 = {1'h0, T83};
  assign T83 = mask_incoherent[2'h2:2'h2];
  assign T371 = {1'h0, T84};
  assign T84 = T372 + T85;
  assign T85 = {1'h0, T86};
  assign T86 = mask_incoherent[1'h1:1'h1];
  assign T372 = {1'h0, T87};
  assign T87 = mask_incoherent[1'h0:1'h0];
  assign T88 = T56 & T47;
  assign T373 = {2'h0, T89};
  assign T89 = release_count - 1'h1;
  assign T374 = {2'h0, T90};
  assign T90 = release_count - 1'h1;
  assign T91 = T98 & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T95 | T94;
  assign T94 = 3'h2 == io_inner_release_bits_r_type;
  assign T95 = T97 | T96;
  assign T96 = 3'h1 == io_inner_release_bits_r_type;
  assign T97 = 3'h0 == io_inner_release_bits_r_type;
  assign T98 = T99 & io_inner_release_valid;
  assign T99 = 3'h1 == state;
  assign T100 = T110 & oacq_data_done;
  assign oacq_data_done = T108 ? T102 : T101;
  assign T101 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T102 = T107 & T103;
  assign T103 = R104 == 2'h3;
  assign T375 = reset ? 2'h0 : T105;
  assign T105 = T107 ? T106 : R104;
  assign T106 = R104 + 2'h1;
  assign T107 = T101 & T108;
  assign T108 = io_outer_acquire_bits_is_builtin_type & T109;
  assign T109 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T110 = T111 & io_outer_acquire_ready;
  assign T111 = T98 & T93;
  assign T112 = pending_outer_write ? 3'h3 : T113;
  assign T113 = pending_outer_read ? 3'h2 : 3'h4;
  assign T114 = T91 & T115;
  assign T115 = release_count == 1'h1;
  assign T116 = pending_outer_read ? 3'h2 : 3'h5;
  assign T117 = T118 & oacq_data_done;
  assign T118 = 3'h3 == state;
  assign T119 = T121 & T120;
  assign T120 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T121 = 3'h2 == state;
  assign T122 = T123 ? 3'h6 : 3'h0;
  assign T123 = T124 ^ 1'h1;
  assign T124 = io_inner_grant_bits_is_builtin_type & T125;
  assign T125 = io_inner_grant_bits_g_type == 4'h0;
  assign T126 = T139 & ignt_data_done;
  assign ignt_data_done = T134 ? T128 : T127;
  assign T127 = io_inner_grant_ready & io_inner_grant_valid;
  assign T128 = T133 & T129;
  assign T129 = R130 == 2'h3;
  assign T376 = reset ? 2'h0 : T131;
  assign T131 = T133 ? T132 : R130;
  assign T132 = R130 + 2'h1;
  assign T133 = T127 & T134;
  assign T134 = io_inner_grant_bits_is_builtin_type ? T138 : T135;
  assign T135 = T137 | T136;
  assign T136 = 4'h1 == io_inner_grant_bits_g_type;
  assign T137 = 4'h0 == io_inner_grant_bits_g_type;
  assign T138 = 4'h5 == io_inner_grant_bits_g_type;
  assign T139 = 3'h5 == state;
  assign T140 = T141 ? 3'h6 : 3'h0;
  assign T141 = T142 ^ 1'h1;
  assign T142 = io_inner_grant_bits_is_builtin_type & T143;
  assign T143 = io_inner_grant_bits_g_type == 4'h0;
  assign T144 = T145 & io_inner_grant_ready;
  assign T145 = 3'h4 == state;
  assign T146 = T147 & io_inner_finish_valid;
  assign T147 = 3'h6 == state;
  assign T149 = T150 | reset;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T154 & T152;
  assign T152 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T153 = T56 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T154 = T156 & T155;
  assign T155 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T156 = T171 & collect_iacq_data;
  assign T377 = reset ? 1'h0 : T157;
  assign T157 = T56 ? T169 : T158;
  assign T158 = T159 ? 1'h0 : collect_iacq_data;
  assign T159 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T167 ? T161 : T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T166 & T162;
  assign T162 = R163 == 2'h3;
  assign T378 = reset ? 2'h0 : T164;
  assign T164 = T166 ? T165 : R163;
  assign T165 = R163 + 2'h1;
  assign T166 = T160 & T167;
  assign T167 = io_inner_acquire_bits_is_builtin_type & T168;
  assign T168 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T169 = io_inner_acquire_bits_is_builtin_type & T170;
  assign T170 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T171 = state != 3'h0;
  assign T173 = T174 | reset;
  assign T174 = T175 ^ 1'h1;
  assign T175 = T178 & T176;
  assign T176 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T177 = T56 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T178 = T180 & T179;
  assign T179 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T180 = T181 & collect_iacq_data;
  assign T181 = state != 3'h0;
  assign T183 = T184 | reset;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T193 & T186;
  assign T186 = T188 | T187;
  assign T187 = 3'h5 == xact_a_type;
  assign T188 = T190 | T189;
  assign T189 = 3'h4 == xact_a_type;
  assign T190 = T192 | T191;
  assign T191 = 3'h2 == xact_a_type;
  assign T192 = 3'h0 == xact_a_type;
  assign T193 = T194 & xact_is_builtin_type;
  assign T194 = state != 3'h0;
  assign io_has_release_match = T195;
  assign T195 = T197 & T196;
  assign T196 = state == 3'h1;
  assign T197 = T199 & T198;
  assign T198 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T199 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T200 = T56 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T201;
  assign T201 = T202 & collect_iacq_data;
  assign T202 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T203;
  assign T203 = T205 & T204;
  assign T204 = collect_iacq_data ^ 1'h1;
  assign T205 = T207 & T206;
  assign T206 = state != 3'h0;
  assign T207 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T208;
  assign T208 = T139 ? io_inner_grant_ready : pending_ognt_ack;
  assign T379 = reset ? 1'h0 : T209;
  assign T209 = T117 ? 1'h1 : T210;
  assign T210 = T100 ? 1'h1 : T211;
  assign T211 = T212 ? 1'h0 : pending_ognt_ack;
  assign T212 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_union = T213;
  assign T213 = T121 ? outer_read_union : T214;
  assign T214 = T118 ? outer_write_acq_union : T215;
  assign T215 = T111 ? outer_write_rel_union : outer_read_union;
  assign outer_write_rel_union = T380;
  assign T380 = {8'h0, T216};
  assign T216 = {T217, 1'h1};
  assign T217 = 1'h1;
  assign outer_write_acq_union = T381;
  assign T381 = {8'h0, T218};
  assign T218 = {T219, 1'h1};
  assign T219 = 1'h1;
  assign outer_read_union = 10'h1c1;
  assign io_outer_acquire_bits_a_type = T220;
  assign T220 = T121 ? outer_read_a_type : T221;
  assign T221 = T118 ? outer_write_acq_a_type : T222;
  assign T222 = T111 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign outer_read_a_type = 3'h1;
  assign io_outer_acquire_bits_is_builtin_type = T223;
  assign T223 = T121 ? outer_read_is_builtin_type : T224;
  assign T224 = T118 ? outer_write_acq_is_builtin_type : T225;
  assign T225 = T111 ? outer_write_rel_is_builtin_type : outer_read_is_builtin_type;
  assign outer_write_rel_is_builtin_type = 1'h1;
  assign outer_write_acq_is_builtin_type = 1'h1;
  assign outer_read_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_data = T226;
  assign T226 = T121 ? outer_read_data : T227;
  assign T227 = T118 ? outer_write_acq_data : T228;
  assign T228 = T111 ? outer_write_rel_data : outer_read_data;
  assign outer_write_rel_data = io_inner_release_bits_data;
  assign outer_write_acq_data = T229;
  assign T229 = T264 ? T250 : T230;
  assign T230 = T248 ? data_buffer_1 : data_buffer_0;
  assign T231 = T238 ? io_inner_acquire_bits_data : T232;
  assign T232 = T233 ? io_inner_acquire_bits_data : data_buffer_0;
  assign T233 = T237 & T234;
  assign T234 = T235[1'h0:1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = io_inner_acquire_bits_addr_beat;
  assign T237 = collect_iacq_data & io_inner_acquire_valid;
  assign T238 = T56 & T239;
  assign T239 = T240[1'h0:1'h0];
  assign T240 = 1'h1 << T241;
  assign T241 = 2'h0;
  assign T242 = T246 ? io_inner_acquire_bits_data : T243;
  assign T243 = T244 ? io_inner_acquire_bits_data : data_buffer_1;
  assign T244 = T237 & T245;
  assign T245 = T235[1'h1:1'h1];
  assign T246 = T56 & T247;
  assign T247 = T240[1'h1:1'h1];
  assign T248 = T249[1'h0:1'h0];
  assign T249 = oacq_data_cnt;
  assign oacq_data_cnt = T108 ? R104 : 2'h0;
  assign T250 = T263 ? data_buffer_3 : data_buffer_2;
  assign T251 = T255 ? io_inner_acquire_bits_data : T252;
  assign T252 = T253 ? io_inner_acquire_bits_data : data_buffer_2;
  assign T253 = T237 & T254;
  assign T254 = T235[2'h2:2'h2];
  assign T255 = T56 & T256;
  assign T256 = T240[2'h2:2'h2];
  assign T257 = T261 ? io_inner_acquire_bits_data : T258;
  assign T258 = T259 ? io_inner_acquire_bits_data : data_buffer_3;
  assign T259 = T237 & T260;
  assign T260 = T235[2'h3:2'h3];
  assign T261 = T56 & T262;
  assign T262 = T240[2'h3:2'h3];
  assign T263 = T249[1'h0:1'h0];
  assign T264 = T249[1'h1:1'h1];
  assign outer_read_data = 4'h0;
  assign io_outer_acquire_bits_addr_beat = T265;
  assign T265 = T121 ? outer_read_addr_beat : T266;
  assign T266 = T118 ? outer_write_acq_addr_beat : T267;
  assign T267 = T111 ? outer_write_rel_addr_beat : outer_read_addr_beat;
  assign outer_write_rel_addr_beat = io_inner_release_bits_addr_beat;
  assign outer_write_acq_addr_beat = oacq_data_cnt;
  assign outer_read_addr_beat = 2'h0;
  assign io_outer_acquire_bits_client_xact_id = T268;
  assign T268 = T121 ? outer_read_client_xact_id : T269;
  assign T269 = T118 ? outer_write_acq_client_xact_id : T270;
  assign T270 = T111 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_write_rel_client_xact_id = 3'h4;
  assign outer_write_acq_client_xact_id = 3'h4;
  assign outer_read_client_xact_id = 3'h4;
  assign io_outer_acquire_bits_addr_block = T271;
  assign T271 = T121 ? outer_read_addr_block : T272;
  assign T272 = T118 ? outer_write_acq_addr_block : T273;
  assign T273 = T111 ? outer_write_rel_addr_block : outer_read_addr_block;
  assign outer_write_rel_addr_block = xact_addr_block;
  assign outer_write_acq_addr_block = xact_addr_block;
  assign outer_read_addr_block = xact_addr_block;
  assign io_outer_acquire_valid = T274;
  assign T274 = T121 ? T301 : T275;
  assign T275 = T118 ? T276 : T111;
  assign T276 = T298 | T277;
  assign T277 = T282 & T278;
  assign T278 = T279 - 1'h1;
  assign T279 = 1'h1 << T280;
  assign T280 = T281 + 2'h1;
  assign T281 = oacq_data_cnt - oacq_data_cnt;
  assign T282 = iacq_data_valid >> oacq_data_cnt;
  assign T382 = reset ? 4'h0 : T283;
  assign T283 = T56 ? T291 : T284;
  assign T284 = T237 ? T285 : iacq_data_valid;
  assign T285 = T289 | T286;
  assign T286 = T383 & T287;
  assign T287 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T383 = T288 ? 4'hf : 4'h0;
  assign T288 = 1'h1;
  assign T289 = iacq_data_valid & T290;
  assign T290 = ~ T287;
  assign T291 = T292 << io_inner_acquire_bits_addr_beat;
  assign T292 = io_inner_acquire_bits_is_builtin_type & T293;
  assign T293 = T295 | T294;
  assign T294 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T295 = T297 | T296;
  assign T296 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T297 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T298 = T300 | T299;
  assign T299 = collect_iacq_data ^ 1'h1;
  assign T300 = pending_ognt_ack ^ 1'h1;
  assign T301 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T302;
  assign T302 = T99 ? T303 : 1'h0;
  assign T303 = T304 | io_outer_acquire_ready;
  assign T304 = T305 ^ 1'h1;
  assign T305 = T307 | T306;
  assign T306 = 3'h2 == io_inner_release_bits_r_type;
  assign T307 = T309 | T308;
  assign T308 = 3'h1 == io_inner_release_bits_r_type;
  assign T309 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T310;
  assign T310 = T384;
  assign T384 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T317;
  assign T317 = T318;
  assign T318 = xact_is_builtin_type ? T323 : T319;
  assign T319 = T322 ? 2'h1 : T320;
  assign T320 = T321 ? 2'h0 : 2'h2;
  assign T321 = xact_a_type == 3'h1;
  assign T322 = xact_a_type == 3'h0;
  assign T323 = T332 ? 2'h2 : T324;
  assign T324 = T331 ? 2'h0 : T325;
  assign T325 = T330 ? 2'h2 : T326;
  assign T326 = T329 ? 2'h0 : T327;
  assign T327 = T328 ? 2'h0 : 2'h2;
  assign T328 = xact_a_type == 3'h4;
  assign T329 = xact_a_type == 3'h2;
  assign T330 = xact_a_type == 3'h0;
  assign T331 = xact_a_type == 3'h3;
  assign T332 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T333;
  assign T333 = xact_addr_block;
  assign io_inner_probe_valid = T334;
  assign T334 = T99 ? T335 : 1'h0;
  assign T335 = pending_probes != 1'h0;
  assign T385 = T386[1'h0:1'h0];
  assign T386 = reset ? 4'h0 : T311;
  assign T311 = T316 ? T388 : T312;
  assign T312 = T88 ? mask_incoherent : T387;
  assign T387 = {3'h0, pending_probes};
  assign T388 = {2'h0, T313};
  assign T313 = T389 & T314;
  assign T314 = ~ T315;
  assign T315 = 1'h1 << 1'h0;
  assign T389 = {1'h0, pending_probes};
  assign T316 = T99 & io_inner_probe_ready;
  assign io_inner_finish_ready = T147;
  assign io_inner_grant_bits_client_id = T336;
  assign T336 = xact_client_id;
  assign io_inner_grant_bits_g_type = T337;
  assign T337 = T390;
  assign T390 = {1'h0, T338};
  assign T338 = xact_is_builtin_type ? T341 : T391;
  assign T391 = {1'h0, T339};
  assign T339 = T340 ? 2'h0 : 2'h1;
  assign T340 = xact_a_type == 3'h0;
  assign T341 = T352 ? 3'h4 : T342;
  assign T342 = T351 ? 3'h5 : T343;
  assign T343 = T350 ? 3'h3 : T344;
  assign T344 = T349 ? 3'h3 : T345;
  assign T345 = T348 ? 3'h4 : T346;
  assign T346 = T347 ? 3'h1 : 3'h3;
  assign T347 = xact_a_type == 3'h5;
  assign T348 = xact_a_type == 3'h4;
  assign T349 = xact_a_type == 3'h3;
  assign T350 = xact_a_type == 3'h2;
  assign T351 = xact_a_type == 3'h1;
  assign T352 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T353;
  assign T353 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T354;
  assign T354 = 3'h4;
  assign io_inner_grant_bits_client_xact_id = T355;
  assign T355 = xact_client_xact_id;
  assign io_inner_grant_bits_data = T356;
  assign T356 = 4'h0;
  assign io_inner_grant_bits_addr_beat = T357;
  assign T357 = 2'h0;
  assign io_inner_grant_valid = T358;
  assign T358 = T145 ? 1'h1 : T359;
  assign T359 = T139 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T360;
  assign T360 = T57 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T182 <= 1'b1;
  if(!T183 && T182 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics, subblock Gets/Puts, or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T172 <= 1'b1;
  if(!T173 && T172 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T148 <= 1'b1;
  if(!T149 && T148 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T146) begin
      state <= 3'h0;
    end else if(T144) begin
      state <= T140;
    end else if(T126) begin
      state <= T122;
    end else if(T119) begin
      state <= 3'h5;
    end else if(T117) begin
      state <= T116;
    end else if(T114) begin
      state <= T112;
    end else if(T73) begin
      state <= T58;
    end else if(T56) begin
      state <= T16;
    end
    if(T56) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T56) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T367;
    if(reset) begin
      R104 <= 2'h0;
    end else if(T107) begin
      R104 <= T106;
    end
    if(reset) begin
      R130 <= 2'h0;
    end else if(T133) begin
      R130 <= T132;
    end
    if(T56) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T56) begin
      collect_iacq_data <= T169;
    end else if(T159) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R163 <= 2'h0;
    end else if(T166) begin
      R163 <= T165;
    end
    if(T56) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T56) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T117) begin
      pending_ognt_ack <= 1'h1;
    end else if(T100) begin
      pending_ognt_ack <= 1'h1;
    end else if(T212) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T238) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T233) begin
      data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T246) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T244) begin
      data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T255) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T253) begin
      data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T261) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T259) begin
      data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T56) begin
      iacq_data_valid <= T291;
    end else if(T237) begin
      iacq_data_valid <= T285;
    end
    pending_probes <= T385;
  end
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_addr_beat,
    input [127:0] io_in_4_bits_data,
    input  io_in_4_bits_client_xact_id,
    input [2:0] io_in_4_bits_manager_xact_id,
    input  io_in_4_bits_is_builtin_type,
    input [3:0] io_in_4_bits_g_type,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_addr_beat,
    input [127:0] io_in_3_bits_data,
    input  io_in_3_bits_client_xact_id,
    input [2:0] io_in_3_bits_manager_xact_id,
    input  io_in_3_bits_is_builtin_type,
    input [3:0] io_in_3_bits_g_type,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_addr_beat,
    input [127:0] io_in_2_bits_data,
    input  io_in_2_bits_client_xact_id,
    input [2:0] io_in_2_bits_manager_xact_id,
    input  io_in_2_bits_is_builtin_type,
    input [3:0] io_in_2_bits_g_type,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [127:0] io_in_1_bits_data,
    input  io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [127:0] io_in_0_bits_data,
    input  io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output io_out_bits_client_xact_id,
    output[2:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T192;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T193;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  locked;
  wire T194;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] R41;
  wire[1:0] T195;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[2:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire[3:0] T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire T55;
  wire[3:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire T71;
  wire[2:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire[127:0] T84;
  wire[127:0] T85;
  wire[127:0] T86;
  wire T87;
  wire[127:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire[1:0] T92;
  wire[1:0] T93;
  wire[1:0] T94;
  wire T95;
  wire[1:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R41 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T192 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T193 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T35 & T30;
  assign T30 = io_out_bits_is_builtin_type ? T34 : T31;
  assign T31 = T33 | T32;
  assign T32 = 4'h1 == io_out_bits_g_type;
  assign T33 = 4'h0 == io_out_bits_g_type;
  assign T34 = 4'h5 == io_out_bits_g_type;
  assign T35 = io_out_ready & io_out_valid;
  assign T194 = reset ? 1'h0 : T36;
  assign T36 = T38 ? 1'h0 : T37;
  assign T37 = T27 ? 1'h1 : locked;
  assign T38 = T35 & T39;
  assign T39 = T40 == 2'h0;
  assign T40 = R41 + 2'h1;
  assign T195 = reset ? 2'h0 : T42;
  assign T42 = T29 ? T40 : R41;
  assign io_out_bits_client_id = T43;
  assign T43 = T51 ? io_in_4_bits_client_id : T44;
  assign T44 = T50 ? T48 : T45;
  assign T45 = T46 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T46 = T47[1'h0:1'h0];
  assign T47 = chosen;
  assign T48 = T49 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T49 = T47[1'h0:1'h0];
  assign T50 = T47[1'h1:1'h1];
  assign T51 = T47[2'h2:2'h2];
  assign io_out_bits_g_type = T52;
  assign T52 = T59 ? io_in_4_bits_g_type : T53;
  assign T53 = T58 ? T56 : T54;
  assign T54 = T55 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign T55 = T47[1'h0:1'h0];
  assign T56 = T57 ? io_in_3_bits_g_type : io_in_2_bits_g_type;
  assign T57 = T47[1'h0:1'h0];
  assign T58 = T47[1'h1:1'h1];
  assign T59 = T47[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T60;
  assign T60 = T67 ? io_in_4_bits_is_builtin_type : T61;
  assign T61 = T66 ? T64 : T62;
  assign T62 = T63 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T63 = T47[1'h0:1'h0];
  assign T64 = T65 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T65 = T47[1'h0:1'h0];
  assign T66 = T47[1'h1:1'h1];
  assign T67 = T47[2'h2:2'h2];
  assign io_out_bits_manager_xact_id = T68;
  assign T68 = T75 ? io_in_4_bits_manager_xact_id : T69;
  assign T69 = T74 ? T72 : T70;
  assign T70 = T71 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign T71 = T47[1'h0:1'h0];
  assign T72 = T73 ? io_in_3_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign T73 = T47[1'h0:1'h0];
  assign T74 = T47[1'h1:1'h1];
  assign T75 = T47[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T76;
  assign T76 = T83 ? io_in_4_bits_client_xact_id : T77;
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T79 = T47[1'h0:1'h0];
  assign T80 = T81 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T81 = T47[1'h0:1'h0];
  assign T82 = T47[1'h1:1'h1];
  assign T83 = T47[2'h2:2'h2];
  assign io_out_bits_data = T84;
  assign T84 = T91 ? io_in_4_bits_data : T85;
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T87 = T47[1'h0:1'h0];
  assign T88 = T89 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T89 = T47[1'h0:1'h0];
  assign T90 = T47[1'h1:1'h1];
  assign T91 = T47[2'h2:2'h2];
  assign io_out_bits_addr_beat = T92;
  assign T92 = T99 ? io_in_4_bits_addr_beat : T93;
  assign T93 = T98 ? T96 : T94;
  assign T94 = T95 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T95 = T47[1'h0:1'h0];
  assign T96 = T97 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T97 = T47[1'h0:1'h0];
  assign T98 = T47[1'h1:1'h1];
  assign T99 = T47[2'h2:2'h2];
  assign io_out_valid = T100;
  assign T100 = T107 ? io_in_4_valid : T101;
  assign T101 = T106 ? T104 : T102;
  assign T102 = T103 ? io_in_1_valid : io_in_0_valid;
  assign T103 = T47[1'h0:1'h0];
  assign T104 = T105 ? io_in_3_valid : io_in_2_valid;
  assign T105 = T47[1'h0:1'h0];
  assign T106 = T47[1'h1:1'h1];
  assign T107 = T47[2'h2:2'h2];
  assign io_in_0_ready = T108;
  assign T108 = T109 & io_out_ready;
  assign T109 = locked ? T127 : T110;
  assign T110 = T126 | T111;
  assign T111 = T112 ^ 1'h1;
  assign T112 = T115 | T113;
  assign T113 = io_in_4_valid & T114;
  assign T114 = last_grant < 3'h4;
  assign T115 = T118 | T116;
  assign T116 = io_in_3_valid & T117;
  assign T117 = last_grant < 3'h3;
  assign T118 = T121 | T119;
  assign T119 = io_in_2_valid & T120;
  assign T120 = last_grant < 3'h2;
  assign T121 = T124 | T122;
  assign T122 = io_in_1_valid & T123;
  assign T123 = last_grant < 3'h1;
  assign T124 = io_in_0_valid & T125;
  assign T125 = last_grant < 3'h0;
  assign T126 = last_grant < 3'h0;
  assign T127 = lockIdx == 3'h0;
  assign io_in_1_ready = T128;
  assign T128 = T129 & io_out_ready;
  assign T129 = locked ? T140 : T130;
  assign T130 = T137 | T131;
  assign T131 = T132 ^ 1'h1;
  assign T132 = T133 | io_in_0_valid;
  assign T133 = T134 | T113;
  assign T134 = T135 | T116;
  assign T135 = T136 | T119;
  assign T136 = T124 | T122;
  assign T137 = T139 & T138;
  assign T138 = last_grant < 3'h1;
  assign T139 = T124 ^ 1'h1;
  assign T140 = lockIdx == 3'h1;
  assign io_in_2_ready = T141;
  assign T141 = T142 & io_out_ready;
  assign T142 = locked ? T155 : T143;
  assign T143 = T151 | T144;
  assign T144 = T145 ^ 1'h1;
  assign T145 = T146 | io_in_1_valid;
  assign T146 = T147 | io_in_0_valid;
  assign T147 = T148 | T113;
  assign T148 = T149 | T116;
  assign T149 = T150 | T119;
  assign T150 = T124 | T122;
  assign T151 = T153 & T152;
  assign T152 = last_grant < 3'h2;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T124 | T122;
  assign T155 = lockIdx == 3'h2;
  assign io_in_3_ready = T156;
  assign T156 = T157 & io_out_ready;
  assign T157 = locked ? T172 : T158;
  assign T158 = T167 | T159;
  assign T159 = T160 ^ 1'h1;
  assign T160 = T161 | io_in_2_valid;
  assign T161 = T162 | io_in_1_valid;
  assign T162 = T163 | io_in_0_valid;
  assign T163 = T164 | T113;
  assign T164 = T165 | T116;
  assign T165 = T166 | T119;
  assign T166 = T124 | T122;
  assign T167 = T169 & T168;
  assign T168 = last_grant < 3'h3;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T171 | T119;
  assign T171 = T124 | T122;
  assign T172 = lockIdx == 3'h3;
  assign io_in_4_ready = T173;
  assign T173 = T174 & io_out_ready;
  assign T174 = locked ? T191 : T175;
  assign T175 = T185 | T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T178 | io_in_3_valid;
  assign T178 = T179 | io_in_2_valid;
  assign T179 = T180 | io_in_1_valid;
  assign T180 = T181 | io_in_0_valid;
  assign T181 = T182 | T113;
  assign T182 = T183 | T116;
  assign T183 = T184 | T119;
  assign T184 = T124 | T122;
  assign T185 = T187 & T186;
  assign T186 = last_grant < 3'h4;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T189 | T116;
  assign T189 = T190 | T119;
  assign T190 = T124 | T122;
  assign T191 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T38) begin
      locked <= 1'h0;
    end else if(T27) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R41 <= 2'h0;
    end else if(T29) begin
      R41 <= T40;
    end
  end
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [1:0] io_in_4_bits_p_type,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [1:0] io_in_3_bits_p_type,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_p_type,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_p_type,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_p_type,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_p_type,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T141;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T142;
  reg  locked;
  wire T143;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  reg [1:0] R22;
  wire[1:0] T144;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[25:0] T41;
  wire[25:0] T42;
  wire[25:0] T43;
  wire T44;
  wire[25:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R22 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T141 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T142 = reset ? 3'h4 : lockIdx;
  assign T143 = reset ? 1'h0 : T18;
  assign T18 = T19 ? 1'h0 : locked;
  assign T19 = T23 & T20;
  assign T20 = T21 == 2'h0;
  assign T21 = R22 + 2'h1;
  assign T144 = reset ? 2'h0 : R22;
  assign T23 = io_out_ready & io_out_valid;
  assign io_out_bits_client_id = T24;
  assign T24 = T32 ? io_in_4_bits_client_id : T25;
  assign T25 = T31 ? T29 : T26;
  assign T26 = T27 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T27 = T28[1'h0:1'h0];
  assign T28 = chosen;
  assign T29 = T30 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T30 = T28[1'h0:1'h0];
  assign T31 = T28[1'h1:1'h1];
  assign T32 = T28[2'h2:2'h2];
  assign io_out_bits_p_type = T33;
  assign T33 = T40 ? io_in_4_bits_p_type : T34;
  assign T34 = T39 ? T37 : T35;
  assign T35 = T36 ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign T36 = T28[1'h0:1'h0];
  assign T37 = T38 ? io_in_3_bits_p_type : io_in_2_bits_p_type;
  assign T38 = T28[1'h0:1'h0];
  assign T39 = T28[1'h1:1'h1];
  assign T40 = T28[2'h2:2'h2];
  assign io_out_bits_addr_block = T41;
  assign T41 = T48 ? io_in_4_bits_addr_block : T42;
  assign T42 = T47 ? T45 : T43;
  assign T43 = T44 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T44 = T28[1'h0:1'h0];
  assign T45 = T46 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T46 = T28[1'h0:1'h0];
  assign T47 = T28[1'h1:1'h1];
  assign T48 = T28[2'h2:2'h2];
  assign io_out_valid = T49;
  assign T49 = T56 ? io_in_4_valid : T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52 ? io_in_1_valid : io_in_0_valid;
  assign T52 = T28[1'h0:1'h0];
  assign T53 = T54 ? io_in_3_valid : io_in_2_valid;
  assign T54 = T28[1'h0:1'h0];
  assign T55 = T28[1'h1:1'h1];
  assign T56 = T28[2'h2:2'h2];
  assign io_in_0_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = locked ? T76 : T59;
  assign T59 = T75 | T60;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T64 | T62;
  assign T62 = io_in_4_valid & T63;
  assign T63 = last_grant < 3'h4;
  assign T64 = T67 | T65;
  assign T65 = io_in_3_valid & T66;
  assign T66 = last_grant < 3'h3;
  assign T67 = T70 | T68;
  assign T68 = io_in_2_valid & T69;
  assign T69 = last_grant < 3'h2;
  assign T70 = T73 | T71;
  assign T71 = io_in_1_valid & T72;
  assign T72 = last_grant < 3'h1;
  assign T73 = io_in_0_valid & T74;
  assign T74 = last_grant < 3'h0;
  assign T75 = last_grant < 3'h0;
  assign T76 = lockIdx == 3'h0;
  assign io_in_1_ready = T77;
  assign T77 = T78 & io_out_ready;
  assign T78 = locked ? T89 : T79;
  assign T79 = T86 | T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T82 | io_in_0_valid;
  assign T82 = T83 | T62;
  assign T83 = T84 | T65;
  assign T84 = T85 | T68;
  assign T85 = T73 | T71;
  assign T86 = T88 & T87;
  assign T87 = last_grant < 3'h1;
  assign T88 = T73 ^ 1'h1;
  assign T89 = lockIdx == 3'h1;
  assign io_in_2_ready = T90;
  assign T90 = T91 & io_out_ready;
  assign T91 = locked ? T104 : T92;
  assign T92 = T100 | T93;
  assign T93 = T94 ^ 1'h1;
  assign T94 = T95 | io_in_1_valid;
  assign T95 = T96 | io_in_0_valid;
  assign T96 = T97 | T62;
  assign T97 = T98 | T65;
  assign T98 = T99 | T68;
  assign T99 = T73 | T71;
  assign T100 = T102 & T101;
  assign T101 = last_grant < 3'h2;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T73 | T71;
  assign T104 = lockIdx == 3'h2;
  assign io_in_3_ready = T105;
  assign T105 = T106 & io_out_ready;
  assign T106 = locked ? T121 : T107;
  assign T107 = T116 | T108;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T110 | io_in_2_valid;
  assign T110 = T111 | io_in_1_valid;
  assign T111 = T112 | io_in_0_valid;
  assign T112 = T113 | T62;
  assign T113 = T114 | T65;
  assign T114 = T115 | T68;
  assign T115 = T73 | T71;
  assign T116 = T118 & T117;
  assign T117 = last_grant < 3'h3;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | T68;
  assign T120 = T73 | T71;
  assign T121 = lockIdx == 3'h3;
  assign io_in_4_ready = T122;
  assign T122 = T123 & io_out_ready;
  assign T123 = locked ? T140 : T124;
  assign T124 = T134 | T125;
  assign T125 = T126 ^ 1'h1;
  assign T126 = T127 | io_in_3_valid;
  assign T127 = T128 | io_in_2_valid;
  assign T128 = T129 | io_in_1_valid;
  assign T129 = T130 | io_in_0_valid;
  assign T130 = T131 | T62;
  assign T131 = T132 | T65;
  assign T132 = T133 | T68;
  assign T133 = T73 | T71;
  assign T134 = T136 & T135;
  assign T135 = last_grant < 3'h4;
  assign T136 = T137 ^ 1'h1;
  assign T137 = T138 | T65;
  assign T138 = T139 | T68;
  assign T139 = T73 | T71;
  assign T140 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T19) begin
      locked <= 1'h0;
    end
    if(reset) begin
      R22 <= 2'h0;
    end
  end
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [2:0] io_in_4_bits_client_xact_id,
    input [1:0] io_in_4_bits_addr_beat,
    input [3:0] io_in_4_bits_data,
    input  io_in_4_bits_is_builtin_type,
    input [2:0] io_in_4_bits_a_type,
    input [9:0] io_in_4_bits_union,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [2:0] io_in_3_bits_client_xact_id,
    input [1:0] io_in_3_bits_addr_beat,
    input [3:0] io_in_3_bits_data,
    input  io_in_3_bits_is_builtin_type,
    input [2:0] io_in_3_bits_a_type,
    input [9:0] io_in_3_bits_union,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [2:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input [3:0] io_in_2_bits_data,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [9:0] io_in_2_bits_union,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [2:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input [3:0] io_in_1_bits_data,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [9:0] io_in_1_bits_union,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [2:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input [3:0] io_in_0_bits_data,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [9:0] io_in_0_bits_union,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[2:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output[3:0] io_out_bits_data,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[9:0] io_out_bits_union,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T189;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T190;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  locked;
  wire T191;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  reg [1:0] R38;
  wire[1:0] T192;
  wire[1:0] T39;
  wire[9:0] T40;
  wire[9:0] T41;
  wire[9:0] T42;
  wire T43;
  wire[2:0] T44;
  wire[9:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire[2:0] T51;
  wire T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[3:0] T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire[3:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[25:0] T89;
  wire[25:0] T90;
  wire[25:0] T91;
  wire T92;
  wire[25:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R38 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T189 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T190 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T32 & T30;
  assign T30 = io_out_bits_is_builtin_type & T31;
  assign T31 = 3'h3 == io_out_bits_a_type;
  assign T32 = io_out_ready & io_out_valid;
  assign T191 = reset ? 1'h0 : T33;
  assign T33 = T35 ? 1'h0 : T34;
  assign T34 = T27 ? 1'h1 : locked;
  assign T35 = T32 & T36;
  assign T36 = T37 == 2'h0;
  assign T37 = R38 + 2'h1;
  assign T192 = reset ? 2'h0 : T39;
  assign T39 = T29 ? T37 : R38;
  assign io_out_bits_union = T40;
  assign T40 = T48 ? io_in_4_bits_union : T41;
  assign T41 = T47 ? T45 : T42;
  assign T42 = T43 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = chosen;
  assign T45 = T46 ? io_in_3_bits_union : io_in_2_bits_union;
  assign T46 = T44[1'h0:1'h0];
  assign T47 = T44[1'h1:1'h1];
  assign T48 = T44[2'h2:2'h2];
  assign io_out_bits_a_type = T49;
  assign T49 = T56 ? io_in_4_bits_a_type : T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T52 = T44[1'h0:1'h0];
  assign T53 = T54 ? io_in_3_bits_a_type : io_in_2_bits_a_type;
  assign T54 = T44[1'h0:1'h0];
  assign T55 = T44[1'h1:1'h1];
  assign T56 = T44[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T57;
  assign T57 = T64 ? io_in_4_bits_is_builtin_type : T58;
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T60 = T44[1'h0:1'h0];
  assign T61 = T62 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T62 = T44[1'h0:1'h0];
  assign T63 = T44[1'h1:1'h1];
  assign T64 = T44[2'h2:2'h2];
  assign io_out_bits_data = T65;
  assign T65 = T72 ? io_in_4_bits_data : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T68 = T44[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T70 = T44[1'h0:1'h0];
  assign T71 = T44[1'h1:1'h1];
  assign T72 = T44[2'h2:2'h2];
  assign io_out_bits_addr_beat = T73;
  assign T73 = T80 ? io_in_4_bits_addr_beat : T74;
  assign T74 = T79 ? T77 : T75;
  assign T75 = T76 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T76 = T44[1'h0:1'h0];
  assign T77 = T78 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T78 = T44[1'h0:1'h0];
  assign T79 = T44[1'h1:1'h1];
  assign T80 = T44[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T81;
  assign T81 = T88 ? io_in_4_bits_client_xact_id : T82;
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T84 = T44[1'h0:1'h0];
  assign T85 = T86 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T86 = T44[1'h0:1'h0];
  assign T87 = T44[1'h1:1'h1];
  assign T88 = T44[2'h2:2'h2];
  assign io_out_bits_addr_block = T89;
  assign T89 = T96 ? io_in_4_bits_addr_block : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T92 = T44[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T94 = T44[1'h0:1'h0];
  assign T95 = T44[1'h1:1'h1];
  assign T96 = T44[2'h2:2'h2];
  assign io_out_valid = T97;
  assign T97 = T104 ? io_in_4_valid : T98;
  assign T98 = T103 ? T101 : T99;
  assign T99 = T100 ? io_in_1_valid : io_in_0_valid;
  assign T100 = T44[1'h0:1'h0];
  assign T101 = T102 ? io_in_3_valid : io_in_2_valid;
  assign T102 = T44[1'h0:1'h0];
  assign T103 = T44[1'h1:1'h1];
  assign T104 = T44[2'h2:2'h2];
  assign io_in_0_ready = T105;
  assign T105 = T106 & io_out_ready;
  assign T106 = locked ? T124 : T107;
  assign T107 = T123 | T108;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T112 | T110;
  assign T110 = io_in_4_valid & T111;
  assign T111 = last_grant < 3'h4;
  assign T112 = T115 | T113;
  assign T113 = io_in_3_valid & T114;
  assign T114 = last_grant < 3'h3;
  assign T115 = T118 | T116;
  assign T116 = io_in_2_valid & T117;
  assign T117 = last_grant < 3'h2;
  assign T118 = T121 | T119;
  assign T119 = io_in_1_valid & T120;
  assign T120 = last_grant < 3'h1;
  assign T121 = io_in_0_valid & T122;
  assign T122 = last_grant < 3'h0;
  assign T123 = last_grant < 3'h0;
  assign T124 = lockIdx == 3'h0;
  assign io_in_1_ready = T125;
  assign T125 = T126 & io_out_ready;
  assign T126 = locked ? T137 : T127;
  assign T127 = T134 | T128;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | io_in_0_valid;
  assign T130 = T131 | T110;
  assign T131 = T132 | T113;
  assign T132 = T133 | T116;
  assign T133 = T121 | T119;
  assign T134 = T136 & T135;
  assign T135 = last_grant < 3'h1;
  assign T136 = T121 ^ 1'h1;
  assign T137 = lockIdx == 3'h1;
  assign io_in_2_ready = T138;
  assign T138 = T139 & io_out_ready;
  assign T139 = locked ? T152 : T140;
  assign T140 = T148 | T141;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T143 | io_in_1_valid;
  assign T143 = T144 | io_in_0_valid;
  assign T144 = T145 | T110;
  assign T145 = T146 | T113;
  assign T146 = T147 | T116;
  assign T147 = T121 | T119;
  assign T148 = T150 & T149;
  assign T149 = last_grant < 3'h2;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T121 | T119;
  assign T152 = lockIdx == 3'h2;
  assign io_in_3_ready = T153;
  assign T153 = T154 & io_out_ready;
  assign T154 = locked ? T169 : T155;
  assign T155 = T164 | T156;
  assign T156 = T157 ^ 1'h1;
  assign T157 = T158 | io_in_2_valid;
  assign T158 = T159 | io_in_1_valid;
  assign T159 = T160 | io_in_0_valid;
  assign T160 = T161 | T110;
  assign T161 = T162 | T113;
  assign T162 = T163 | T116;
  assign T163 = T121 | T119;
  assign T164 = T166 & T165;
  assign T165 = last_grant < 3'h3;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | T116;
  assign T168 = T121 | T119;
  assign T169 = lockIdx == 3'h3;
  assign io_in_4_ready = T170;
  assign T170 = T171 & io_out_ready;
  assign T171 = locked ? T188 : T172;
  assign T172 = T182 | T173;
  assign T173 = T174 ^ 1'h1;
  assign T174 = T175 | io_in_3_valid;
  assign T175 = T176 | io_in_2_valid;
  assign T176 = T177 | io_in_1_valid;
  assign T177 = T178 | io_in_0_valid;
  assign T178 = T179 | T110;
  assign T179 = T180 | T113;
  assign T180 = T181 | T116;
  assign T181 = T121 | T119;
  assign T182 = T184 & T183;
  assign T183 = last_grant < 3'h4;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T186 | T113;
  assign T186 = T187 | T116;
  assign T187 = T121 | T119;
  assign T188 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T35) begin
      locked <= 1'h0;
    end else if(T27) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R38 <= 2'h0;
    end else if(T29) begin
      R38 <= T37;
    end
  end
endmodule

module ClientUncachedTileLinkIOArbiter(input clk, input reset,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [25:0] io_in_4_acquire_bits_addr_block,
    input [2:0] io_in_4_acquire_bits_client_xact_id,
    input [1:0] io_in_4_acquire_bits_addr_beat,
    input [3:0] io_in_4_acquire_bits_data,
    input  io_in_4_acquire_bits_is_builtin_type,
    input [2:0] io_in_4_acquire_bits_a_type,
    input [9:0] io_in_4_acquire_bits_union,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_addr_beat,
    output[3:0] io_in_4_grant_bits_data,
    output[2:0] io_in_4_grant_bits_client_xact_id,
    output io_in_4_grant_bits_manager_xact_id,
    output io_in_4_grant_bits_is_builtin_type,
    output[3:0] io_in_4_grant_bits_g_type,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [25:0] io_in_3_acquire_bits_addr_block,
    input [2:0] io_in_3_acquire_bits_client_xact_id,
    input [1:0] io_in_3_acquire_bits_addr_beat,
    input [3:0] io_in_3_acquire_bits_data,
    input  io_in_3_acquire_bits_is_builtin_type,
    input [2:0] io_in_3_acquire_bits_a_type,
    input [9:0] io_in_3_acquire_bits_union,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_addr_beat,
    output[3:0] io_in_3_grant_bits_data,
    output[2:0] io_in_3_grant_bits_client_xact_id,
    output io_in_3_grant_bits_manager_xact_id,
    output io_in_3_grant_bits_is_builtin_type,
    output[3:0] io_in_3_grant_bits_g_type,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [25:0] io_in_2_acquire_bits_addr_block,
    input [2:0] io_in_2_acquire_bits_client_xact_id,
    input [1:0] io_in_2_acquire_bits_addr_beat,
    input [3:0] io_in_2_acquire_bits_data,
    input  io_in_2_acquire_bits_is_builtin_type,
    input [2:0] io_in_2_acquire_bits_a_type,
    input [9:0] io_in_2_acquire_bits_union,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_addr_beat,
    output[3:0] io_in_2_grant_bits_data,
    output[2:0] io_in_2_grant_bits_client_xact_id,
    output io_in_2_grant_bits_manager_xact_id,
    output io_in_2_grant_bits_is_builtin_type,
    output[3:0] io_in_2_grant_bits_g_type,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [25:0] io_in_1_acquire_bits_addr_block,
    input [2:0] io_in_1_acquire_bits_client_xact_id,
    input [1:0] io_in_1_acquire_bits_addr_beat,
    input [3:0] io_in_1_acquire_bits_data,
    input  io_in_1_acquire_bits_is_builtin_type,
    input [2:0] io_in_1_acquire_bits_a_type,
    input [9:0] io_in_1_acquire_bits_union,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_addr_beat,
    output[3:0] io_in_1_grant_bits_data,
    output[2:0] io_in_1_grant_bits_client_xact_id,
    output io_in_1_grant_bits_manager_xact_id,
    output io_in_1_grant_bits_is_builtin_type,
    output[3:0] io_in_1_grant_bits_g_type,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [25:0] io_in_0_acquire_bits_addr_block,
    input [2:0] io_in_0_acquire_bits_client_xact_id,
    input [1:0] io_in_0_acquire_bits_addr_beat,
    input [3:0] io_in_0_acquire_bits_data,
    input  io_in_0_acquire_bits_is_builtin_type,
    input [2:0] io_in_0_acquire_bits_a_type,
    input [9:0] io_in_0_acquire_bits_union,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_addr_beat,
    output[3:0] io_in_0_grant_bits_data,
    output[2:0] io_in_0_grant_bits_client_xact_id,
    output io_in_0_grant_bits_manager_xact_id,
    output io_in_0_grant_bits_is_builtin_type,
    output[3:0] io_in_0_grant_bits_g_type,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output[3:0] io_out_acquire_bits_data,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[9:0] io_out_acquire_bits_union,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [3:0] io_out_grant_bits_data,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type
);

  wire[2:0] T30;
  wire[5:0] T0;
  wire[2:0] T31;
  wire[5:0] T1;
  wire[2:0] T32;
  wire[5:0] T2;
  wire[2:0] T33;
  wire[5:0] T3;
  wire[2:0] T34;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T21;
  wire T23;
  wire T25;
  wire T27;
  wire T29;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[25:0] LockingRRArbiter_io_out_bits_addr_block;
  wire[2:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_addr_beat;
  wire[3:0] LockingRRArbiter_io_out_bits_data;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_a_type;
  wire[9:0] LockingRRArbiter_io_out_bits_union;


  assign T30 = T0[2'h2:1'h0];
  assign T0 = {io_in_0_acquire_bits_client_xact_id, 3'h0};
  assign T31 = T1[2'h2:1'h0];
  assign T1 = {io_in_1_acquire_bits_client_xact_id, 3'h1};
  assign T32 = T2[2'h2:1'h0];
  assign T2 = {io_in_2_acquire_bits_client_xact_id, 3'h2};
  assign T33 = T3[2'h2:1'h0];
  assign T3 = {io_in_3_acquire_bits_client_xact_id, 3'h3};
  assign T34 = T4[2'h2:1'h0];
  assign T4 = {io_in_4_acquire_bits_client_xact_id, 3'h4};
  assign io_out_grant_ready = T5;
  assign T5 = T18 ? io_in_4_grant_ready : T6;
  assign T6 = T16 ? io_in_3_grant_ready : T7;
  assign T7 = T14 ? io_in_2_grant_ready : T8;
  assign T8 = T12 ? io_in_1_grant_ready : T9;
  assign T9 = T10 ? io_in_0_grant_ready : 1'h0;
  assign T10 = T11 == 3'h0;
  assign T11 = io_out_grant_bits_client_xact_id;
  assign T12 = T13 == 3'h1;
  assign T13 = io_out_grant_bits_client_xact_id;
  assign T14 = T15 == 3'h2;
  assign T15 = io_out_grant_bits_client_xact_id;
  assign T16 = T17 == 3'h3;
  assign T17 = io_out_grant_bits_client_xact_id;
  assign T18 = T19 == 3'h4;
  assign T19 = io_out_grant_bits_client_xact_id;
  assign io_out_acquire_bits_union = LockingRRArbiter_io_out_bits_union;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_data = LockingRRArbiter_io_out_bits_data;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_io_out_bits_addr_block;
  assign io_out_acquire_valid = LockingRRArbiter_io_out_valid;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_client_xact_id = 3'h0;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_valid = T21;
  assign T21 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_io_in_0_ready;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_client_xact_id = 3'h0;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_valid = T23;
  assign T23 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_io_in_1_ready;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_client_xact_id = 3'h0;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_valid = T25;
  assign T25 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = LockingRRArbiter_io_in_2_ready;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_client_xact_id = 3'h0;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_valid = T27;
  assign T27 = T16 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = LockingRRArbiter_io_in_3_ready;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_client_xact_id = 3'h0;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_valid = T29;
  assign T29 = T18 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = LockingRRArbiter_io_in_4_ready;
  LockingRRArbiter_4 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_addr_block( io_in_4_acquire_bits_addr_block ),
       .io_in_4_bits_client_xact_id( T34 ),
       .io_in_4_bits_addr_beat( io_in_4_acquire_bits_addr_beat ),
       .io_in_4_bits_data( io_in_4_acquire_bits_data ),
       .io_in_4_bits_is_builtin_type( io_in_4_acquire_bits_is_builtin_type ),
       .io_in_4_bits_a_type( io_in_4_acquire_bits_a_type ),
       .io_in_4_bits_union( io_in_4_acquire_bits_union ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_addr_block( io_in_3_acquire_bits_addr_block ),
       .io_in_3_bits_client_xact_id( T33 ),
       .io_in_3_bits_addr_beat( io_in_3_acquire_bits_addr_beat ),
       .io_in_3_bits_data( io_in_3_acquire_bits_data ),
       .io_in_3_bits_is_builtin_type( io_in_3_acquire_bits_is_builtin_type ),
       .io_in_3_bits_a_type( io_in_3_acquire_bits_a_type ),
       .io_in_3_bits_union( io_in_3_acquire_bits_union ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_addr_block( io_in_2_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( T32 ),
       .io_in_2_bits_addr_beat( io_in_2_acquire_bits_addr_beat ),
       .io_in_2_bits_data( io_in_2_acquire_bits_data ),
       .io_in_2_bits_is_builtin_type( io_in_2_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( io_in_2_acquire_bits_a_type ),
       .io_in_2_bits_union( io_in_2_acquire_bits_union ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_addr_block( io_in_1_acquire_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T31 ),
       .io_in_1_bits_addr_beat( io_in_1_acquire_bits_addr_beat ),
       .io_in_1_bits_data( io_in_1_acquire_bits_data ),
       .io_in_1_bits_is_builtin_type( io_in_1_acquire_bits_is_builtin_type ),
       .io_in_1_bits_a_type( io_in_1_acquire_bits_a_type ),
       .io_in_1_bits_union( io_in_1_acquire_bits_union ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_addr_block( io_in_0_acquire_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T30 ),
       .io_in_0_bits_addr_beat( io_in_0_acquire_bits_addr_beat ),
       .io_in_0_bits_data( io_in_0_acquire_bits_data ),
       .io_in_0_bits_is_builtin_type( io_in_0_acquire_bits_is_builtin_type ),
       .io_in_0_bits_a_type( io_in_0_acquire_bits_a_type ),
       .io_in_0_bits_union( io_in_0_acquire_bits_union ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( LockingRRArbiter_io_out_bits_addr_beat ),
       .io_out_bits_data( LockingRRArbiter_io_out_bits_data ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( LockingRRArbiter_io_out_bits_a_type ),
       .io_out_bits_union( LockingRRArbiter_io_out_bits_union )
       //.io_chosen(  )
  );
endmodule

module L2BroadcastHub(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input  io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input [127:0] io_inner_acquire_bits_data,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[127:0] io_inner_grant_bits_data,
    output io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [25:0] io_inner_release_bits_addr_block,
    input  io_inner_release_bits_client_xact_id,
    input [1:0] io_inner_release_bits_addr_beat,
    input [127:0] io_inner_release_bits_data,
    input [2:0] io_inner_release_bits_r_type,
    input  io_inner_release_bits_voluntary,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [127:0] io_outer_grant_bits_data,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[4:0] releaseMatches;
  wire[4:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[3:0] T228;
  wire[127:0] T229;
  wire[127:0] T230;
  wire[127:0] T231;
  wire[127:0] T232;
  wire[127:0] T233;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  reg [1:0] rel_data_cnt;
  wire[1:0] T234;
  wire[1:0] T14;
  wire[1:0] T15;
  wire vwbdq_enq;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T235;
  wire[2:0] T236;
  wire[2:0] T237;
  wire[2:0] T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T25;
  wire T26;
  wire[9:0] T243;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T244;
  wire[1:0] T245;
  wire[1:0] T246;
  wire T247;
  wire[3:0] T31;
  reg [3:0] sdq_val;
  wire[3:0] T248;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[3:0] T249;
  wire sdq_enq;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T250;
  wire free_sdq;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[3:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T251;
  wire T252;
  wire T70;
  wire T71;
  wire[2:0] acquire_idx;
  wire[2:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire[2:0] T256;
  wire T257;
  wire[4:0] acquireReadys;
  wire[4:0] T73;
  wire[2:0] T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire T258;
  wire T259;
  wire T260;
  wire[2:0] T261;
  wire[2:0] T262;
  wire[2:0] T263;
  wire[2:0] T264;
  wire T265;
  wire[4:0] acquireMatches;
  wire[4:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T266;
  wire T267;
  wire T268;
  wire T82;
  wire T83;
  wire T84;
  wire block_acquires;
  wire T85;
  wire sdq_rdy;
  wire T86;
  wire T87;
  wire[4:0] acquireConflicts;
  wire[4:0] T88;
  wire[2:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[9:0] T269;
  wire[3:0] T100;
  wire[3:0] T101;
  wire[1:0] T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[9:0] T270;
  wire[3:0] T116;
  wire[3:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[9:0] T271;
  wire[3:0] T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[3:0] T140;
  wire[3:0] T141;
  wire[1:0] T142;
  wire[1:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[9:0] T272;
  wire[3:0] T148;
  wire[3:0] T149;
  wire[1:0] T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire[16:0] T156;
  wire T157;
  wire[15:0] T158;
  wire[15:0] T273;
  wire T159;
  wire[127:0] T160;
  wire[127:0] T161;
  wire[127:0] T162;
  wire[127:0] T163;
  reg [127:0] vwbdq_0;
  wire[127:0] T164;
  wire T165;
  wire T166;
  wire[3:0] T167;
  wire[1:0] T168;
  reg [127:0] vwbdq_1;
  wire[127:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] T173;
  wire[127:0] T174;
  reg [127:0] vwbdq_2;
  wire[127:0] T175;
  wire T176;
  wire T177;
  reg [127:0] vwbdq_3;
  wire[127:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[127:0] T184;
  wire[127:0] T185;
  reg [127:0] sdq_0;
  wire[127:0] T186;
  wire T187;
  wire T188;
  wire[3:0] T189;
  wire[1:0] T190;
  reg [127:0] sdq_1;
  wire[127:0] T191;
  wire T192;
  wire T193;
  wire T194;
  wire[1:0] T195;
  wire[127:0] T196;
  reg [127:0] sdq_2;
  wire[127:0] T197;
  wire T198;
  wire T199;
  reg [127:0] sdq_3;
  wire[127:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire[2:0] T209;
  wire[2:0] T210;
  wire T211;
  wire[4:0] releaseReadys;
  wire[4:0] T212;
  wire[2:0] T213;
  wire[1:0] T214;
  wire[1:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[2:0] T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_probe_valid;
  wire BroadcastVoluntaryReleaseTracker_io_inner_release_ready;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type;
  wire[9:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union;
  wire BroadcastVoluntaryReleaseTracker_io_outer_grant_ready;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_match;
  wire BroadcastVoluntaryReleaseTracker_io_has_release_match;
  wire BroadcastAcquireTracker_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_data;
  wire BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_g_type;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_finish_ready;
  wire BroadcastAcquireTracker_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_release_ready;
  wire BroadcastAcquireTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_a_type;
  wire[9:0] BroadcastAcquireTracker_io_outer_acquire_bits_union;
  wire BroadcastAcquireTracker_io_outer_grant_ready;
  wire BroadcastAcquireTracker_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_io_has_acquire_match;
  wire BroadcastAcquireTracker_io_has_release_match;
  wire BroadcastAcquireTracker_1_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_1_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_data;
  wire BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_g_type;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_finish_ready;
  wire BroadcastAcquireTracker_1_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_release_ready;
  wire BroadcastAcquireTracker_1_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type;
  wire[9:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_union;
  wire BroadcastAcquireTracker_1_io_outer_grant_ready;
  wire BroadcastAcquireTracker_1_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_1_io_has_acquire_match;
  wire BroadcastAcquireTracker_1_io_has_release_match;
  wire BroadcastAcquireTracker_2_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_2_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_data;
  wire BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_g_type;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_finish_ready;
  wire BroadcastAcquireTracker_2_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_release_ready;
  wire BroadcastAcquireTracker_2_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type;
  wire[9:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_union;
  wire BroadcastAcquireTracker_2_io_outer_grant_ready;
  wire BroadcastAcquireTracker_2_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_2_io_has_acquire_match;
  wire BroadcastAcquireTracker_2_io_has_release_match;
  wire BroadcastAcquireTracker_3_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_3_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_data;
  wire BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_g_type;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_finish_ready;
  wire BroadcastAcquireTracker_3_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_release_ready;
  wire BroadcastAcquireTracker_3_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type;
  wire[9:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_union;
  wire BroadcastAcquireTracker_3_io_outer_grant_ready;
  wire BroadcastAcquireTracker_3_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_3_io_has_acquire_match;
  wire BroadcastAcquireTracker_3_io_has_release_match;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire LockingRRArbiter_io_out_bits_client_xact_id;
  wire[2:0] LockingRRArbiter_io_out_bits_manager_xact_id;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[3:0] LockingRRArbiter_io_out_bits_g_type;
  wire[1:0] LockingRRArbiter_io_out_bits_client_id;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[25:0] LockingRRArbiter_1_io_out_bits_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_p_type;
  wire[1:0] LockingRRArbiter_1_io_out_bits_client_id;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_4_grant_bits_data;
  wire[2:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_3_grant_bits_data;
  wire[2:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_2_grant_bits_data;
  wire[2:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_1_grant_bits_data;
  wire[2:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire[3:0] outer_arb_io_in_0_grant_bits_data;
  wire[2:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire outer_arb_io_out_acquire_valid;
  wire[25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire[2:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire[1:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire[3:0] outer_arb_io_out_acquire_bits_data;
  wire outer_arb_io_out_acquire_bits_is_builtin_type;
  wire[2:0] outer_arb_io_out_acquire_bits_a_type;
  wire[9:0] outer_arb_io_out_acquire_bits_union;
  wire outer_arb_io_out_grant_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    rel_data_cnt = {1{$random}};
    sdq_val = {1{$random}};
    vwbdq_0 = {4{$random}};
    vwbdq_1 = {4{$random}};
    vwbdq_2 = {4{$random}};
    vwbdq_3 = {4{$random}};
    sdq_0 = {4{$random}};
    sdq_1 = {4{$random}};
    sdq_2 = {4{$random}};
    sdq_3 = {4{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_inner_release_valid & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = releaseMatches != 5'h0;
  assign releaseMatches = T6;
  assign T6 = {T9, T7};
  assign T7 = {BroadcastAcquireTracker_1_io_has_release_match, T8};
  assign T8 = {BroadcastAcquireTracker_io_has_release_match, BroadcastVoluntaryReleaseTracker_io_has_release_match};
  assign T9 = {BroadcastAcquireTracker_3_io_has_release_match, BroadcastAcquireTracker_2_io_has_release_match};
  assign T228 = io_outer_grant_bits_data[2'h3:1'h0];
  assign T229 = {124'h0, BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data};
  assign T230 = {124'h0, BroadcastAcquireTracker_io_inner_grant_bits_data};
  assign T231 = {124'h0, BroadcastAcquireTracker_1_io_inner_grant_bits_data};
  assign T232 = {124'h0, BroadcastAcquireTracker_2_io_inner_grant_bits_data};
  assign T233 = {124'h0, BroadcastAcquireTracker_3_io_inner_grant_bits_data};
  assign T10 = T11;
  assign T11 = {T13, T12};
  assign T12 = 2'h2;
  assign T13 = rel_data_cnt;
  assign T234 = reset ? 2'h0 : T14;
  assign T14 = vwbdq_enq ? T15 : rel_data_cnt;
  assign T15 = rel_data_cnt + 2'h1;
  assign vwbdq_enq = T21 & T16;
  assign T16 = T18 | T17;
  assign T17 = 3'h2 == io_inner_release_bits_r_type;
  assign T18 = T20 | T19;
  assign T19 = 3'h1 == io_inner_release_bits_r_type;
  assign T20 = 3'h0 == io_inner_release_bits_r_type;
  assign T21 = T22 & io_inner_release_bits_voluntary;
  assign T22 = io_inner_release_ready & io_inner_release_valid;
  assign T23 = io_inner_release_valid & T24;
  assign T24 = T235 == 3'h4;
  assign T235 = T242 ? 1'h0 : T236;
  assign T236 = T241 ? 1'h1 : T237;
  assign T237 = T240 ? 2'h2 : T238;
  assign T238 = T239 ? 2'h3 : 3'h4;
  assign T239 = releaseMatches[2'h3:2'h3];
  assign T240 = releaseMatches[2'h2:2'h2];
  assign T241 = releaseMatches[1'h1:1'h1];
  assign T242 = releaseMatches[1'h0:1'h0];
  assign T25 = io_inner_finish_valid & T26;
  assign T26 = io_inner_finish_bits_manager_xact_id == 3'h4;
  assign T243 = io_inner_acquire_bits_union[4'h9:1'h0];
  assign T27 = T28;
  assign T28 = {T30, T29};
  assign T29 = 2'h0;
  assign T30 = T244;
  assign T244 = T252 ? 1'h0 : T245;
  assign T245 = T251 ? 1'h1 : T246;
  assign T246 = T247 ? 2'h2 : 2'h3;
  assign T247 = T31[2'h2:2'h2];
  assign T31 = ~ sdq_val;
  assign T248 = reset ? 4'h0 : T32;
  assign T32 = T69 ? T33 : sdq_val;
  assign T33 = T53 | T34;
  assign T34 = T43 & T35;
  assign T35 = 4'h0 - T249;
  assign T249 = {3'h0, sdq_enq};
  assign sdq_enq = T42 & T36;
  assign T36 = io_inner_acquire_bits_is_builtin_type & T37;
  assign T37 = T39 | T38;
  assign T38 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T39 = T41 | T40;
  assign T40 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T41 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T42 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T43 = T52 ? 4'h1 : T44;
  assign T44 = T51 ? 4'h2 : T45;
  assign T45 = T50 ? 4'h4 : T46;
  assign T46 = T47 ? 4'h8 : 4'h0;
  assign T47 = T48[2'h3:2'h3];
  assign T48 = ~ T49;
  assign T49 = sdq_val[2'h3:1'h0];
  assign T50 = T48[2'h2:2'h2];
  assign T51 = T48[1'h1:1'h1];
  assign T52 = T48[1'h0:1'h0];
  assign T53 = sdq_val & T54;
  assign T54 = ~ T55;
  assign T55 = T67 & T56;
  assign T56 = 4'h0 - T250;
  assign T250 = {3'h0, free_sdq};
  assign free_sdq = T59 & T57;
  assign T57 = T58 == 2'h0;
  assign T58 = outer_arb_io_out_acquire_bits_data[1'h1:1'h0];
  assign T59 = T66 & T60;
  assign T60 = io_outer_acquire_bits_is_builtin_type & T61;
  assign T61 = T63 | T62;
  assign T62 = 3'h4 == io_outer_acquire_bits_a_type;
  assign T63 = T65 | T64;
  assign T64 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T65 = 3'h2 == io_outer_acquire_bits_a_type;
  assign T66 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T67 = 1'h1 << T68;
  assign T68 = outer_arb_io_out_acquire_bits_data[2'h3:2'h2];
  assign T69 = io_outer_acquire_valid | sdq_enq;
  assign T251 = T31[1'h1:1'h1];
  assign T252 = T31[1'h0:1'h0];
  assign T70 = T83 & T71;
  assign T71 = acquire_idx == 3'h4;
  assign acquire_idx = T82 ? T261 : T253;
  assign T253 = T260 ? 1'h0 : T254;
  assign T254 = T259 ? 1'h1 : T255;
  assign T255 = T258 ? 2'h2 : T256;
  assign T256 = T257 ? 2'h3 : 3'h4;
  assign T257 = acquireReadys[2'h3:2'h3];
  assign acquireReadys = T73;
  assign T73 = {T76, T74};
  assign T74 = {BroadcastAcquireTracker_1_io_inner_acquire_ready, T75};
  assign T75 = {BroadcastAcquireTracker_io_inner_acquire_ready, BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready};
  assign T76 = {BroadcastAcquireTracker_3_io_inner_acquire_ready, BroadcastAcquireTracker_2_io_inner_acquire_ready};
  assign T258 = acquireReadys[2'h2:2'h2];
  assign T259 = acquireReadys[1'h1:1'h1];
  assign T260 = acquireReadys[1'h0:1'h0];
  assign T261 = T268 ? 1'h0 : T262;
  assign T262 = T267 ? 1'h1 : T263;
  assign T263 = T266 ? 2'h2 : T264;
  assign T264 = T265 ? 2'h3 : 3'h4;
  assign T265 = acquireMatches[2'h3:2'h3];
  assign acquireMatches = T78;
  assign T78 = {T81, T79};
  assign T79 = {BroadcastAcquireTracker_1_io_has_acquire_match, T80};
  assign T80 = {BroadcastAcquireTracker_io_has_acquire_match, BroadcastVoluntaryReleaseTracker_io_has_acquire_match};
  assign T81 = {BroadcastAcquireTracker_3_io_has_acquire_match, BroadcastAcquireTracker_2_io_has_acquire_match};
  assign T266 = acquireMatches[2'h2:2'h2];
  assign T267 = acquireMatches[1'h1:1'h1];
  assign T268 = acquireMatches[1'h0:1'h0];
  assign T82 = acquireMatches != 5'h0;
  assign T83 = io_inner_acquire_valid & T84;
  assign T84 = block_acquires ^ 1'h1;
  assign block_acquires = T87 | T85;
  assign T85 = sdq_rdy ^ 1'h1;
  assign sdq_rdy = T86 ^ 1'h1;
  assign T86 = sdq_val == 4'hf;
  assign T87 = acquireConflicts != 5'h0;
  assign acquireConflicts = T88;
  assign T88 = {T91, T89};
  assign T89 = {BroadcastAcquireTracker_1_io_has_acquire_conflict, T90};
  assign T90 = {BroadcastAcquireTracker_io_has_acquire_conflict, BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict};
  assign T91 = {BroadcastAcquireTracker_3_io_has_acquire_conflict, BroadcastAcquireTracker_2_io_has_acquire_conflict};
  assign T92 = T93;
  assign T93 = {T95, T94};
  assign T94 = 2'h2;
  assign T95 = rel_data_cnt;
  assign T96 = io_inner_release_valid & T97;
  assign T97 = T235 == 3'h3;
  assign T98 = io_inner_finish_valid & T99;
  assign T99 = io_inner_finish_bits_manager_xact_id == 3'h3;
  assign T269 = io_inner_acquire_bits_union[4'h9:1'h0];
  assign T100 = T101;
  assign T101 = {T103, T102};
  assign T102 = 2'h0;
  assign T103 = T244;
  assign T104 = T106 & T105;
  assign T105 = acquire_idx == 3'h3;
  assign T106 = io_inner_acquire_valid & T107;
  assign T107 = block_acquires ^ 1'h1;
  assign T108 = T109;
  assign T109 = {T111, T110};
  assign T110 = 2'h2;
  assign T111 = rel_data_cnt;
  assign T112 = io_inner_release_valid & T113;
  assign T113 = T235 == 3'h2;
  assign T114 = io_inner_finish_valid & T115;
  assign T115 = io_inner_finish_bits_manager_xact_id == 3'h2;
  assign T270 = io_inner_acquire_bits_union[4'h9:1'h0];
  assign T116 = T117;
  assign T117 = {T119, T118};
  assign T118 = 2'h0;
  assign T119 = T244;
  assign T120 = T122 & T121;
  assign T121 = acquire_idx == 3'h2;
  assign T122 = io_inner_acquire_valid & T123;
  assign T123 = block_acquires ^ 1'h1;
  assign T124 = T125;
  assign T125 = {T127, T126};
  assign T126 = 2'h2;
  assign T127 = rel_data_cnt;
  assign T128 = io_inner_release_valid & T129;
  assign T129 = T235 == 3'h1;
  assign T130 = io_inner_finish_valid & T131;
  assign T131 = io_inner_finish_bits_manager_xact_id == 3'h1;
  assign T271 = io_inner_acquire_bits_union[4'h9:1'h0];
  assign T132 = T133;
  assign T133 = {T135, T134};
  assign T134 = 2'h0;
  assign T135 = T244;
  assign T136 = T138 & T137;
  assign T137 = acquire_idx == 3'h1;
  assign T138 = io_inner_acquire_valid & T139;
  assign T139 = block_acquires ^ 1'h1;
  assign T140 = T141;
  assign T141 = {T143, T142};
  assign T142 = 2'h1;
  assign T143 = rel_data_cnt;
  assign T144 = io_inner_release_valid & T145;
  assign T145 = T235 == 3'h0;
  assign T146 = io_inner_finish_valid & T147;
  assign T147 = io_inner_finish_bits_manager_xact_id == 3'h0;
  assign T272 = io_inner_acquire_bits_union[4'h9:1'h0];
  assign T148 = T149;
  assign T149 = {T151, T150};
  assign T150 = 2'h0;
  assign T151 = T244;
  assign T152 = T154 & T153;
  assign T153 = acquire_idx == 3'h0;
  assign T154 = io_inner_acquire_valid & T155;
  assign T155 = block_acquires ^ 1'h1;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_union = T156;
  assign T156 = {T158, T157};
  assign T157 = outer_arb_io_out_acquire_bits_union[1'h0:1'h0];
  assign T158 = 16'h0 - T273;
  assign T273 = {15'h0, T159};
  assign T159 = outer_arb_io_out_acquire_bits_union[1'h1:1'h1];
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_data = T160;
  assign T160 = T205 ? T184 : T161;
  assign T161 = T183 ? T162 : io_inner_release_bits_data;
  assign T162 = T182 ? T174 : T163;
  assign T163 = T172 ? vwbdq_1 : vwbdq_0;
  assign T164 = T165 ? io_inner_release_bits_data : vwbdq_0;
  assign T165 = vwbdq_enq & T166;
  assign T166 = T167[1'h0:1'h0];
  assign T167 = 1'h1 << T168;
  assign T168 = rel_data_cnt;
  assign T169 = T170 ? io_inner_release_bits_data : vwbdq_1;
  assign T170 = vwbdq_enq & T171;
  assign T171 = T167[1'h1:1'h1];
  assign T172 = T173[1'h0:1'h0];
  assign T173 = T68;
  assign T174 = T181 ? vwbdq_3 : vwbdq_2;
  assign T175 = T176 ? io_inner_release_bits_data : vwbdq_2;
  assign T176 = vwbdq_enq & T177;
  assign T177 = T167[2'h2:2'h2];
  assign T178 = T179 ? io_inner_release_bits_data : vwbdq_3;
  assign T179 = vwbdq_enq & T180;
  assign T180 = T167[2'h3:2'h3];
  assign T181 = T173[1'h0:1'h0];
  assign T182 = T173[1'h1:1'h1];
  assign T183 = T58 == 2'h1;
  assign T184 = T204 ? T196 : T185;
  assign T185 = T194 ? sdq_1 : sdq_0;
  assign T186 = T187 ? io_inner_acquire_bits_data : sdq_0;
  assign T187 = sdq_enq & T188;
  assign T188 = T189[1'h0:1'h0];
  assign T189 = 1'h1 << T190;
  assign T190 = T244;
  assign T191 = T192 ? io_inner_acquire_bits_data : sdq_1;
  assign T192 = sdq_enq & T193;
  assign T193 = T189[1'h1:1'h1];
  assign T194 = T195[1'h0:1'h0];
  assign T195 = T68;
  assign T196 = T203 ? sdq_3 : sdq_2;
  assign T197 = T198 ? io_inner_acquire_bits_data : sdq_2;
  assign T198 = sdq_enq & T199;
  assign T199 = T189[2'h2:2'h2];
  assign T200 = T201 ? io_inner_acquire_bits_data : sdq_3;
  assign T201 = sdq_enq & T202;
  assign T202 = T189[2'h3:2'h3];
  assign T203 = T195[1'h0:1'h0];
  assign T204 = T195[1'h1:1'h1];
  assign T205 = T58 == 2'h0;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T206;
  assign T206 = T211 & T207;
  assign T207 = T208 - 1'h1;
  assign T208 = 1'h1 << T209;
  assign T209 = T210 + 3'h1;
  assign T210 = T235 - T235;
  assign T211 = releaseReadys >> T235;
  assign releaseReadys = T212;
  assign T212 = {T215, T213};
  assign T213 = {BroadcastAcquireTracker_1_io_inner_release_ready, T214};
  assign T214 = {BroadcastAcquireTracker_io_inner_release_ready, BroadcastVoluntaryReleaseTracker_io_inner_release_ready};
  assign T215 = {BroadcastAcquireTracker_3_io_inner_release_ready, BroadcastAcquireTracker_2_io_inner_release_ready};
  assign io_inner_probe_bits_client_id = LockingRRArbiter_1_io_out_bits_client_id;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_1_io_out_bits_p_type;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_1_io_out_bits_addr_block;
  assign io_inner_probe_valid = LockingRRArbiter_1_io_out_valid;
  assign io_inner_finish_ready = T216;
  assign T216 = T224 ? BroadcastAcquireTracker_3_io_inner_finish_ready : T217;
  assign T217 = T223 ? T221 : T218;
  assign T218 = T219 ? BroadcastAcquireTracker_io_inner_finish_ready : BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  assign T219 = T220[1'h0:1'h0];
  assign T220 = io_inner_finish_bits_manager_xact_id;
  assign T221 = T222 ? BroadcastAcquireTracker_2_io_inner_finish_ready : BroadcastAcquireTracker_1_io_inner_finish_ready;
  assign T222 = T220[1'h0:1'h0];
  assign T223 = T220[1'h1:1'h1];
  assign T224 = T220[2'h2:2'h2];
  assign io_inner_grant_bits_client_id = LockingRRArbiter_io_out_bits_client_id;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_io_out_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = LockingRRArbiter_io_out_valid;
  assign io_inner_acquire_ready = T225;
  assign T225 = T227 & T226;
  assign T226 = block_acquires ^ 1'h1;
  assign T227 = acquireReadys != 5'h0;
  BroadcastVoluntaryReleaseTracker BroadcastVoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T152 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( T148 ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( T272 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_0_ready ),
       .io_inner_grant_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastVoluntaryReleaseTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T146 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_inner_probe_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_addr_block(  )
       //.io_inner_probe_bits_p_type(  )
       //.io_inner_probe_bits_client_id(  )
       .io_inner_release_ready( BroadcastVoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T144 ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_data( T140 ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_has_acquire_conflict( BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastVoluntaryReleaseTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastVoluntaryReleaseTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_0 BroadcastAcquireTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T136 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( T132 ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( T271 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_1_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T130 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_io_inner_release_ready ),
       .io_inner_release_valid( T128 ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_data( T124 ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_1 BroadcastAcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T120 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( T116 ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( T270 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_2_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_1_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_1_io_inner_finish_ready ),
       .io_inner_finish_valid( T114 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T112 ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_data( T108 ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_1_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_1_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_1_io_has_release_match )
  );
  BroadcastAcquireTracker_2 BroadcastAcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T104 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( T100 ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( T269 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_3_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_2_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_2_io_inner_finish_ready ),
       .io_inner_finish_valid( T98 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T96 ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_data( T92 ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_2_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_2_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_2_io_has_release_match )
  );
  BroadcastAcquireTracker_3 BroadcastAcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T70 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( T27 ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( T243 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_4_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_3_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_3_io_inner_finish_ready ),
       .io_inner_finish_valid( T25 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T23 ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_data( T10 ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_3_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_3_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_3_io_has_release_match )
  );
  LockingRRArbiter_2 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_in_4_bits_data( T233 ),
       .io_in_4_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_in_4_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_in_4_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_in_4_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_in_3_bits_data( T232 ),
       .io_in_3_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_in_3_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_in_3_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_in_3_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_in_2_bits_data( T231 ),
       .io_in_2_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_in_2_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_in_2_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_in_2_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_in_1_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_in_1_bits_data( T230 ),
       .io_in_1_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_1_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_1_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_1_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_in_0_bits_data( T229 ),
       .io_in_0_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_0_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_0_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_0_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_in_0_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       //.io_out_bits_data(  )
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( LockingRRArbiter_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( LockingRRArbiter_io_out_bits_g_type ),
       .io_out_bits_client_id( LockingRRArbiter_io_out_bits_client_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_in_4_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_in_3_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_in_2_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_in_1_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_in_1_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_addr_block(  )
       //.io_in_0_bits_p_type(  )
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_1_io_out_bits_addr_block ),
       .io_out_bits_p_type( LockingRRArbiter_1_io_out_bits_p_type ),
       .io_out_bits_client_id( LockingRRArbiter_1_io_out_bits_client_id )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign LockingRRArbiter_1.io_in_0_bits_addr_block = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_p_type = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  ClientUncachedTileLinkIOArbiter outer_arb(.clk(clk), .reset(reset),
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_in_4_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_in_4_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_in_4_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_in_4_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_in_4_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_in_4_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_in_4_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_in_4_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_in_4_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_in_4_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_in_4_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_in_4_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_in_3_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_in_3_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_in_3_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_in_3_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_in_3_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_in_3_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_in_3_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_in_3_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_in_3_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_in_3_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_in_3_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_in_3_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_in_2_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_in_2_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_in_2_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_in_2_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_in_2_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_in_2_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_in_2_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_in_2_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_in_2_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_in_2_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_in_2_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_in_2_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_in_1_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_1_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_1_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_in_1_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_1_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_in_1_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_in_1_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_in_1_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_in_1_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_in_1_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_in_1_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_in_1_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_in_0_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_0_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_0_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_in_0_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_0_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_in_0_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_in_0_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_in_0_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_in_0_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_in_0_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_in_0_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_in_0_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( outer_arb_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( outer_arb_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( outer_arb_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_data( outer_arb_io_out_acquire_bits_data ),
       .io_out_acquire_bits_is_builtin_type( outer_arb_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( outer_arb_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( outer_arb_io_out_acquire_bits_union ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_addr_beat( io_outer_grant_bits_addr_beat ),
       .io_out_grant_bits_data( T228 ),
       .io_out_grant_bits_client_xact_id( io_outer_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( io_outer_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( io_outer_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( io_outer_grant_bits_g_type )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Non-voluntary release should always have a Tracker waiting for it.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      rel_data_cnt <= 2'h0;
    end else if(vwbdq_enq) begin
      rel_data_cnt <= T15;
    end
    if(reset) begin
      sdq_val <= 4'h0;
    end else if(T69) begin
      sdq_val <= T33;
    end
    if(T165) begin
      vwbdq_0 <= io_inner_release_bits_data;
    end
    if(T170) begin
      vwbdq_1 <= io_inner_release_bits_data;
    end
    if(T176) begin
      vwbdq_2 <= io_inner_release_bits_data;
    end
    if(T179) begin
      vwbdq_3 <= io_inner_release_bits_data;
    end
    if(T187) begin
      sdq_0 <= io_inner_acquire_bits_data;
    end
    if(T192) begin
      sdq_1 <= io_inner_acquire_bits_data;
    end
    if(T198) begin
      sdq_2 <= io_inner_acquire_bits_data;
    end
    if(T201) begin
      sdq_3 <= io_inner_acquire_bits_data;
    end
  end
endmodule

module FinishQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_fin_manager_xact_id,
    input  io_enq_bits_dst,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_fin_manager_xact_id,
    output io_deq_bits_dst,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  reg [1:0] ram [1:0];
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_dst = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_fin_manager_xact_id, io_enq_bits_dst};
  assign io_deq_bits_fin_manager_xact_id = T15;
  assign T15 = T11[1'h1:1'h1];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module FinishUnit_3(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input  io_grant_bits_header_src,
    input  io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [127:0] io_grant_bits_payload_data,
    input [2:0] io_grant_bits_payload_client_xact_id,
    input  io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[127:0] io_refill_bits_data,
    output[2:0] io_refill_bits_client_xact_id,
    output io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    input  io_finish_ready,
    output io_finish_valid,
    output io_finish_bits_header_src,
    output io_finish_bits_header_dst,
    output io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T29;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T18 & T2;
  assign T2 = T14 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T29 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T13 : T12;
  assign T12 = 4'h0 == io_grant_bits_payload_g_type;
  assign T13 = 4'h5 == io_grant_bits_payload_g_type;
  assign T14 = T15 ^ 1'h1;
  assign T15 = io_grant_bits_payload_is_builtin_type ? T17 : T16;
  assign T16 = 4'h0 == io_grant_bits_payload_g_type;
  assign T17 = 4'h5 == io_grant_bits_payload_g_type;
  assign T18 = T22 & T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = io_grant_bits_payload_is_builtin_type & T21;
  assign T21 = io_grant_bits_payload_g_type == 4'h0;
  assign T22 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 1'h0;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = io_grant_valid;
  assign io_grant_ready = T23;
  assign T23 = T24 & io_refill_ready;
  assign T24 = FinishQueue_io_enq_ready | T25;
  assign T25 = T26 ^ 1'h1;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_grant_bits_payload_is_builtin_type & T28;
  assign T28 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue_1 FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_3(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [2:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[127:0] io_client_grant_bits_data,
    output[2:0] io_client_grant_bits_client_xact_id,
    output io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [25:0] io_client_release_bits_addr_block,
    input [2:0] io_client_release_bits_client_xact_id,
    input [1:0] io_client_release_bits_addr_beat,
    input [127:0] io_client_release_bits_data,
    input [2:0] io_client_release_bits_r_type,
    input  io_client_release_bits_voluntary,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output io_network_acquire_bits_header_src,
    output io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[2:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input  io_network_grant_bits_header_src,
    input  io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [127:0] io_network_grant_bits_payload_data,
    input [2:0] io_network_grant_bits_payload_client_xact_id,
    input  io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output io_network_finish_bits_header_src,
    output io_network_finish_bits_header_dst,
    output io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input  io_network_probe_bits_header_src,
    input  io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output io_network_release_bits_header_src,
    output io_network_release_bits_header_dst,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[2:0] io_network_release_bits_payload_client_xact_id,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[127:0] io_network_release_bits_payload_data,
    output[2:0] io_network_release_bits_payload_r_type,
    output io_network_release_bits_payload_voluntary
);

  wire rel_with_header_bits_payload_voluntary;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire[127:0] rel_with_header_bits_payload_data;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[2:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire rel_with_header_bits_header_dst;
  wire rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[2:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire acq_with_header_bits_header_dst;
  wire acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[127:0] finisher_io_refill_bits_data;
  wire[2:0] finisher_io_refill_bits_client_xact_id;
  wire finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire finisher_io_finish_valid;
  wire finisher_io_finish_bits_header_src;
  wire finisher_io_finish_bits_header_dst;
  wire finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 1'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 1'h0;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 1'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 1'h0;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_3 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module TileLinkEnqueuer(
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input  io_client_acquire_bits_header_src,
    input  io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [2:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output io_client_grant_bits_header_src,
    output io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[127:0] io_client_grant_bits_payload_data,
    output[2:0] io_client_grant_bits_payload_client_xact_id,
    output io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input  io_client_finish_bits_header_src,
    input  io_client_finish_bits_header_dst,
    input  io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output io_client_probe_bits_header_src,
    output io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input  io_client_release_bits_header_src,
    input  io_client_release_bits_header_dst,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [2:0] io_client_release_bits_payload_client_xact_id,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [127:0] io_client_release_bits_payload_data,
    input [2:0] io_client_release_bits_payload_r_type,
    input  io_client_release_bits_payload_voluntary,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output io_manager_acquire_bits_header_src,
    output io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[2:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input  io_manager_grant_bits_header_src,
    input  io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [127:0] io_manager_grant_bits_payload_data,
    input [2:0] io_manager_grant_bits_payload_client_xact_id,
    input  io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output io_manager_finish_bits_header_src,
    output io_manager_finish_bits_header_dst,
    output io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input  io_manager_probe_bits_header_src,
    input  io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output io_manager_release_bits_header_src,
    output io_manager_release_bits_header_dst,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[2:0] io_manager_release_bits_payload_client_xact_id,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[127:0] io_manager_release_bits_payload_data,
    output[2:0] io_manager_release_bits_payload_r_type,
    output io_manager_release_bits_payload_voluntary
);



  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_acquire_ready = io_manager_acquire_ready;
endmodule

module ManagerTileLinkNetworkPort_1(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output[2:0] io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output[127:0] io_manager_acquire_bits_data,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [127:0] io_manager_grant_bits_data,
    input [2:0] io_manager_grant_bits_client_xact_id,
    input  io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input  io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input  io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[25:0] io_manager_release_bits_addr_block,
    output[2:0] io_manager_release_bits_client_xact_id,
    output[1:0] io_manager_release_bits_addr_beat,
    output[127:0] io_manager_release_bits_data,
    output[2:0] io_manager_release_bits_r_type,
    output io_manager_release_bits_voluntary,
    output io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input  io_network_acquire_bits_header_src,
    input  io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input [2:0] io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output io_network_grant_bits_header_src,
    output io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[127:0] io_network_grant_bits_payload_data,
    output[2:0] io_network_grant_bits_payload_client_xact_id,
    output io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input  io_network_finish_bits_header_src,
    input  io_network_finish_bits_header_dst,
    input  io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output io_network_probe_bits_header_src,
    output io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input  io_network_release_bits_header_src,
    input  io_network_release_bits_header_dst,
    input [25:0] io_network_release_bits_payload_addr_block,
    input [2:0] io_network_release_bits_payload_client_xact_id,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [127:0] io_network_release_bits_payload_data,
    input [2:0] io_network_release_bits_payload_r_type,
    input  io_network_release_bits_payload_voluntary
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[3:0] T7;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[127:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] T18;
  wire[127:0] T19;
  wire[1:0] T20;
  wire[2:0] T21;
  wire[25:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[16:0] T28;
  wire[2:0] T29;
  wire T30;
  wire[127:0] T31;
  wire[1:0] T32;
  wire[2:0] T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = io_manager_probe_bits_client_id;
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 1'h0;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_g_type = T7;
  assign T7 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T8;
  assign T8 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T9;
  assign T9 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T10;
  assign T10 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_data = T11;
  assign T11 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = io_manager_grant_bits_client_id;
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 1'h0;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src;
  assign io_manager_release_bits_voluntary = T17;
  assign T17 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_r_type = T18;
  assign T18 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_data = T19;
  assign T19 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_addr_beat = T20;
  assign T20 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_bits_client_xact_id = T21;
  assign T21 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T22;
  assign T22 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src;
  assign io_manager_acquire_bits_union = T28;
  assign T28 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T29;
  assign T29 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T30;
  assign T30 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_data = T31;
  assign T31 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module RocketChipTileLinkArbiter_1(input clk, input reset,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [25:0] io_clients_0_acquire_bits_addr_block,
    input [2:0] io_clients_0_acquire_bits_client_xact_id,
    input [1:0] io_clients_0_acquire_bits_addr_beat,
    input [127:0] io_clients_0_acquire_bits_data,
    input  io_clients_0_acquire_bits_is_builtin_type,
    input [2:0] io_clients_0_acquire_bits_a_type,
    input [16:0] io_clients_0_acquire_bits_union,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_addr_beat,
    output[127:0] io_clients_0_grant_bits_data,
    output[2:0] io_clients_0_grant_bits_client_xact_id,
    output io_clients_0_grant_bits_manager_xact_id,
    output io_clients_0_grant_bits_is_builtin_type,
    output[3:0] io_clients_0_grant_bits_g_type,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[25:0] io_clients_0_probe_bits_addr_block,
    output[1:0] io_clients_0_probe_bits_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [25:0] io_clients_0_release_bits_addr_block,
    input [2:0] io_clients_0_release_bits_client_xact_id,
    input [1:0] io_clients_0_release_bits_addr_beat,
    input [127:0] io_clients_0_release_bits_data,
    input [2:0] io_clients_0_release_bits_r_type,
    input  io_clients_0_release_bits_voluntary,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[25:0] io_managers_0_acquire_bits_addr_block,
    output[2:0] io_managers_0_acquire_bits_client_xact_id,
    output[1:0] io_managers_0_acquire_bits_addr_beat,
    output[127:0] io_managers_0_acquire_bits_data,
    output io_managers_0_acquire_bits_is_builtin_type,
    output[2:0] io_managers_0_acquire_bits_a_type,
    output[16:0] io_managers_0_acquire_bits_union,
    output io_managers_0_acquire_bits_client_id,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_addr_beat,
    input [127:0] io_managers_0_grant_bits_data,
    input [2:0] io_managers_0_grant_bits_client_xact_id,
    input  io_managers_0_grant_bits_manager_xact_id,
    input  io_managers_0_grant_bits_is_builtin_type,
    input [3:0] io_managers_0_grant_bits_g_type,
    input  io_managers_0_grant_bits_client_id,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output io_managers_0_finish_bits_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [25:0] io_managers_0_probe_bits_addr_block,
    input [1:0] io_managers_0_probe_bits_p_type,
    input  io_managers_0_probe_bits_client_id,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[25:0] io_managers_0_release_bits_addr_block,
    output[2:0] io_managers_0_release_bits_client_xact_id,
    output[1:0] io_managers_0_release_bits_addr_beat,
    output[127:0] io_managers_0_release_bits_data,
    output[2:0] io_managers_0_release_bits_r_type,
    output io_managers_0_release_bits_voluntary,
    output io_managers_0_release_bits_client_id
);

  wire TileLinkEnqueuer_io_client_acquire_ready;
  wire TileLinkEnqueuer_io_client_grant_valid;
  wire TileLinkEnqueuer_io_client_grant_bits_header_src;
  wire TileLinkEnqueuer_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_client_grant_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_io_client_finish_ready;
  wire TileLinkEnqueuer_io_client_probe_valid;
  wire TileLinkEnqueuer_io_client_probe_bits_header_src;
  wire TileLinkEnqueuer_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_io_client_release_ready;
  wire TileLinkEnqueuer_io_manager_acquire_valid;
  wire TileLinkEnqueuer_io_manager_acquire_bits_header_src;
  wire TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_io_manager_grant_ready;
  wire TileLinkEnqueuer_io_manager_finish_valid;
  wire TileLinkEnqueuer_io_manager_finish_bits_header_src;
  wire TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  wire TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_manager_probe_ready;
  wire TileLinkEnqueuer_io_manager_release_valid;
  wire TileLinkEnqueuer_io_manager_release_bits_header_src;
  wire TileLinkEnqueuer_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_io_manager_finish_valid;
  wire ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_io_manager_release_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_io_network_grant_valid;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_header_src;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat;
  wire[127:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type;
  wire ManagerTileLinkNetworkPort_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_io_network_probe_valid;
  wire ManagerTileLinkNetworkPort_io_network_probe_bits_header_src;
  wire ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_io_network_release_ready;
  wire TileLinkEnqueuer_1_io_client_acquire_ready;
  wire TileLinkEnqueuer_1_io_client_grant_valid;
  wire TileLinkEnqueuer_1_io_client_grant_bits_header_src;
  wire TileLinkEnqueuer_1_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type;
  wire TileLinkEnqueuer_1_io_client_finish_ready;
  wire TileLinkEnqueuer_1_io_client_probe_valid;
  wire TileLinkEnqueuer_1_io_client_probe_bits_header_src;
  wire TileLinkEnqueuer_1_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_1_io_client_release_ready;
  wire TileLinkEnqueuer_1_io_manager_acquire_valid;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_header_src;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  wire TileLinkEnqueuer_1_io_manager_grant_ready;
  wire TileLinkEnqueuer_1_io_manager_finish_valid;
  wire TileLinkEnqueuer_1_io_manager_finish_bits_header_src;
  wire TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  wire TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_manager_probe_ready;
  wire TileLinkEnqueuer_1_io_manager_release_valid;
  wire TileLinkEnqueuer_1_io_manager_release_bits_header_src;
  wire TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  wire[127:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  wire ClientTileLinkNetworkPort_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_client_grant_bits_data;
  wire[2:0] ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  wire ClientTileLinkNetworkPort_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_io_client_release_ready;
  wire ClientTileLinkNetworkPort_io_network_acquire_valid;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_header_src;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union;
  wire ClientTileLinkNetworkPort_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_io_network_finish_valid;
  wire ClientTileLinkNetworkPort_io_network_finish_bits_header_src;
  wire ClientTileLinkNetworkPort_io_network_finish_bits_header_dst;
  wire ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_io_network_release_valid;
  wire ClientTileLinkNetworkPort_io_network_release_bits_header_src;
  wire ClientTileLinkNetworkPort_io_network_release_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat;
  wire[127:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_data;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary;


  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_io_manager_release_valid;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_io_manager_probe_ready;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_io_manager_finish_valid;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_io_manager_grant_ready;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  assign io_clients_0_release_ready = ClientTileLinkNetworkPort_io_client_release_ready;
  assign io_clients_0_probe_bits_p_type = ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  assign io_clients_0_probe_bits_addr_block = ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  assign io_clients_0_probe_valid = ClientTileLinkNetworkPort_io_client_probe_valid;
  assign io_clients_0_grant_bits_g_type = ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  assign io_clients_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  assign io_clients_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  assign io_clients_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  assign io_clients_0_grant_bits_data = ClientTileLinkNetworkPort_io_client_grant_bits_data;
  assign io_clients_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  assign io_clients_0_grant_valid = ClientTileLinkNetworkPort_io_client_grant_valid;
  assign io_clients_0_acquire_ready = ClientTileLinkNetworkPort_io_client_acquire_ready;
  ClientTileLinkNetworkPort_3 ClientTileLinkNetworkPort(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_0_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_0_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_0_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_0_acquire_bits_addr_beat ),
       .io_client_acquire_bits_data( io_clients_0_acquire_bits_data ),
       .io_client_acquire_bits_is_builtin_type( io_clients_0_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_0_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_0_acquire_bits_union ),
       .io_client_grant_ready( io_clients_0_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_io_client_grant_bits_data ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_io_client_grant_bits_g_type ),
       .io_client_probe_ready( io_clients_0_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_io_client_release_ready ),
       .io_client_release_valid( io_clients_0_release_valid ),
       .io_client_release_bits_addr_block( io_clients_0_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_0_release_bits_client_xact_id ),
       .io_client_release_bits_addr_beat( io_clients_0_release_bits_addr_beat ),
       .io_client_release_bits_data( io_clients_0_release_bits_data ),
       .io_client_release_bits_r_type( io_clients_0_release_bits_r_type ),
       .io_client_release_bits_voluntary( io_clients_0_release_bits_voluntary ),
       .io_network_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_network_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer TileLinkEnqueuer(
       .io_client_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_manager_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_manager_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_manager_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_manager_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary )
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort(
       .io_manager_acquire_ready( io_managers_0_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_0_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_0_grant_bits_addr_beat ),
       .io_manager_grant_bits_data( io_managers_0_grant_bits_data ),
       .io_manager_grant_bits_client_xact_id( io_managers_0_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_0_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_0_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_0_grant_bits_g_type ),
       .io_manager_grant_bits_client_id( io_managers_0_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_0_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_0_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_0_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_0_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_0_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_0_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_io_manager_release_valid ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_io_manager_release_bits_data ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_io_manager_release_bits_r_type ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_network_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary )
  );
  TileLinkEnqueuer TileLinkEnqueuer_1(
       .io_client_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_client_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_client_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_client_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_client_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_client_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_client_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_client_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_client_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_client_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_client_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_client_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_client_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_manager_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary )
  );
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [127:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input  io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [127:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input  io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output[2:0] io_out_bits_client_xact_id,
    output io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output io_out_bits_client_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire[2:0] T5;
  wire[127:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_client_id = T0;
  assign T0 = T1 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T1 = chosen;
  assign io_out_bits_g_type = T2;
  assign T2 = T1 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign io_out_bits_is_builtin_type = T3;
  assign T3 = T1 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = T4;
  assign T4 = T1 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_data = T6;
  assign T6 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module MemIOTileLinkIOConverter(input clk, input reset,
    output io_tl_acquire_ready,
    input  io_tl_acquire_valid,
    input [25:0] io_tl_acquire_bits_addr_block,
    input [2:0] io_tl_acquire_bits_client_xact_id,
    input [1:0] io_tl_acquire_bits_addr_beat,
    input [127:0] io_tl_acquire_bits_data,
    input  io_tl_acquire_bits_is_builtin_type,
    input [2:0] io_tl_acquire_bits_a_type,
    input [16:0] io_tl_acquire_bits_union,
    input  io_tl_acquire_bits_client_id,
    input  io_tl_grant_ready,
    output io_tl_grant_valid,
    output[1:0] io_tl_grant_bits_addr_beat,
    output[127:0] io_tl_grant_bits_data,
    output[2:0] io_tl_grant_bits_client_xact_id,
    output io_tl_grant_bits_manager_xact_id,
    output io_tl_grant_bits_is_builtin_type,
    output[3:0] io_tl_grant_bits_g_type,
    output io_tl_grant_bits_client_id,
    output io_tl_finish_ready,
    input  io_tl_finish_valid,
    input  io_tl_finish_bits_manager_xact_id,
    input  io_tl_probe_ready,
    output io_tl_probe_valid,
    //output[25:0] io_tl_probe_bits_addr_block
    //output[1:0] io_tl_probe_bits_p_type
    //output io_tl_probe_bits_client_id
    output io_tl_release_ready,
    input  io_tl_release_valid,
    input [25:0] io_tl_release_bits_addr_block,
    input [2:0] io_tl_release_bits_client_xact_id,
    input [1:0] io_tl_release_bits_addr_beat,
    input [127:0] io_tl_release_bits_data,
    input [2:0] io_tl_release_bits_r_type,
    input  io_tl_release_bits_voluntary,
    input  io_tl_release_bits_client_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[5:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [5:0] io_mem_resp_bits_tag
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire[3:0] T119;
  wire[2:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[2:0] T8;
  wire[2:0] T120;
  wire[4:0] T9;
  wire[127:0] T10;
  wire[1:0] T11;
  reg [1:0] tl_cnt_in;
  wire[1:0] T121;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg [5:0] tag_out;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[5:0] T122;
  wire[4:0] T23;
  wire[3:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg  active_out;
  wire T123;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  make_grant_ack;
  wire T124;
  wire T37;
  wire T38;
  wire T39;
  wire acq_has_data;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  reg  tl_done_out;
  wire T125;
  wire T48;
  wire T49;
  wire tl_wrap_out;
  wire T50;
  reg [1:0] tl_cnt_out;
  wire[1:0] T126;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire rel_has_data;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  reg  has_data;
  wire T127;
  wire T66;
  wire T67;
  reg  cmd_sent_out;
  wire T128;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[5:0] T129;
  wire[4:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire[3:0] T77;
  wire[3:0] T130;
  wire[2:0] T78;
  reg  data_from_rel;
  wire T131;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T132;
  wire[4:0] T84;
  wire[127:0] T85;
  wire[1:0] T86;
  wire[127:0] T87;
  wire[127:0] T88;
  wire[127:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire[5:0] T105;
  wire[5:0] T106;
  wire[5:0] T133;
  wire[5:0] T134;
  wire[25:0] T107;
  wire[25:0] T108;
  reg [25:0] addr_out;
  wire[25:0] T109;
  wire[25:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire gnt_arb_io_in_1_ready;
  wire gnt_arb_io_in_0_ready;
  wire gnt_arb_io_out_valid;
  wire[1:0] gnt_arb_io_out_bits_addr_beat;
  wire[127:0] gnt_arb_io_out_bits_data;
  wire[2:0] gnt_arb_io_out_bits_client_xact_id;
  wire gnt_arb_io_out_bits_manager_xact_id;
  wire gnt_arb_io_out_bits_is_builtin_type;
  wire[3:0] gnt_arb_io_out_bits_g_type;
  wire gnt_arb_io_out_bits_client_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    tl_cnt_in = {1{$random}};
    tag_out = {1{$random}};
    active_out = {1{$random}};
    make_grant_ack = {1{$random}};
    tl_done_out = {1{$random}};
    tl_cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    data_from_rel = {1{$random}};
    addr_out = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_tl_probe_bits_client_id = {1{$random}};
//  assign io_tl_probe_bits_p_type = {1{$random}};
//  assign io_tl_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T1;
  assign T1 = io_mem_resp_bits_tag[3'h4:3'h4];
  assign T2 = T119;
  assign T119 = {1'h0, T3};
  assign T3 = T4 ? 3'h5 : 3'h0;
  assign T4 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign T5 = T6;
  assign T6 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign T7 = 1'h0;
  assign T8 = T120;
  assign T120 = T9[2'h2:1'h0];
  assign T9 = io_mem_resp_bits_tag >> 1'h1;
  assign T10 = io_mem_resp_bits_data;
  assign T11 = tl_cnt_in;
  assign T121 = reset ? 2'h0 : T12;
  assign T12 = T14 ? T13 : tl_cnt_in;
  assign T13 = tl_cnt_in + 2'h1;
  assign T14 = T18 & T15;
  assign T15 = io_tl_grant_bits_is_builtin_type ? T17 : T16;
  assign T16 = 4'h0 == io_tl_grant_bits_g_type;
  assign T17 = 4'h5 == io_tl_grant_bits_g_type;
  assign T18 = io_tl_grant_ready & io_tl_grant_valid;
  assign T19 = T20;
  assign T20 = tag_out[3'h4:3'h4];
  assign T21 = T74 ? T129 : T22;
  assign T22 = T25 ? T122 : tag_out;
  assign T122 = {1'h0, T23};
  assign T23 = {io_tl_release_bits_client_id, T24};
  assign T24 = {io_tl_release_bits_client_xact_id, io_tl_release_bits_voluntary};
  assign T25 = T26 & io_tl_release_valid;
  assign T26 = T29 & T27;
  assign T27 = io_mem_req_data_ready & T28;
  assign T28 = io_tl_release_valid | io_tl_acquire_valid;
  assign T29 = active_out ^ 1'h1;
  assign T123 = reset ? 1'h0 : T30;
  assign T30 = T34 ? 1'h0 : T31;
  assign T31 = T26 ? T32 : active_out;
  assign T32 = T33 | io_mem_req_data_valid;
  assign T33 = io_mem_req_cmd_ready ^ 1'h1;
  assign T34 = active_out & T35;
  assign T35 = T63 & T36;
  assign T36 = make_grant_ack ^ 1'h1;
  assign T124 = reset ? 1'h0 : T37;
  assign T37 = T45 ? 1'h0 : T38;
  assign T38 = T74 ? acq_has_data : T39;
  assign T39 = T25 ? 1'h1 : make_grant_ack;
  assign acq_has_data = io_tl_acquire_bits_is_builtin_type & T40;
  assign T40 = T42 | T41;
  assign T41 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T42 = T44 | T43;
  assign T43 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T44 = 3'h2 == io_tl_acquire_bits_a_type;
  assign T45 = T46 & gnt_arb_io_in_1_ready;
  assign T46 = active_out & T47;
  assign T47 = tl_done_out & make_grant_ack;
  assign T125 = reset ? 1'h0 : T48;
  assign T48 = T62 ? 1'h1 : T49;
  assign T49 = T26 ? tl_wrap_out : tl_done_out;
  assign tl_wrap_out = T53 & T50;
  assign T50 = tl_cnt_out == 2'h3;
  assign T126 = reset ? 2'h0 : T51;
  assign T51 = T53 ? T52 : tl_cnt_out;
  assign T52 = tl_cnt_out + 2'h1;
  assign T53 = T60 | T54;
  assign T54 = T59 & rel_has_data;
  assign rel_has_data = T56 | T55;
  assign T55 = 3'h2 == io_tl_release_bits_r_type;
  assign T56 = T58 | T57;
  assign T57 = 3'h1 == io_tl_release_bits_r_type;
  assign T58 = 3'h0 == io_tl_release_bits_r_type;
  assign T59 = io_tl_release_ready & io_tl_release_valid;
  assign T60 = T61 & acq_has_data;
  assign T61 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T62 = active_out & tl_wrap_out;
  assign T63 = cmd_sent_out & T64;
  assign T64 = T65 | tl_done_out;
  assign T65 = has_data ^ 1'h1;
  assign T127 = reset ? 1'h0 : T66;
  assign T66 = T74 ? acq_has_data : T67;
  assign T67 = T25 ? rel_has_data : has_data;
  assign T128 = reset ? 1'h0 : T68;
  assign T68 = active_out ? T70 : T69;
  assign T69 = T26 ? io_mem_req_cmd_ready : cmd_sent_out;
  assign T70 = cmd_sent_out | T71;
  assign T71 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign T129 = {1'h0, T72};
  assign T72 = {io_tl_acquire_bits_client_id, T73};
  assign T73 = {io_tl_acquire_bits_client_xact_id, io_tl_acquire_bits_is_builtin_type};
  assign T74 = T26 & T75;
  assign T75 = T76 & io_tl_acquire_valid;
  assign T76 = io_tl_release_valid ^ 1'h1;
  assign T77 = T130;
  assign T130 = {1'h0, T78};
  assign T78 = data_from_rel ? 3'h0 : 3'h3;
  assign T131 = reset ? 1'h0 : T79;
  assign T79 = T74 ? 1'h0 : T80;
  assign T80 = T25 ? 1'h1 : data_from_rel;
  assign T81 = 1'h1;
  assign T82 = 1'h0;
  assign T83 = T132;
  assign T132 = T84[2'h2:1'h0];
  assign T84 = tag_out >> 1'h1;
  assign T85 = 128'h0;
  assign T86 = 2'h0;
  assign io_mem_resp_ready = gnt_arb_io_in_0_ready;
  assign io_mem_req_data_bits_data = T87;
  assign T87 = T74 ? io_tl_acquire_bits_data : T88;
  assign T88 = T25 ? io_tl_release_bits_data : T89;
  assign T89 = data_from_rel ? io_tl_release_bits_data : io_tl_acquire_bits_data;
  assign io_mem_req_data_valid = T90;
  assign T90 = T100 ? io_tl_acquire_valid : T91;
  assign T91 = T96 ? io_tl_release_valid : T92;
  assign T92 = T29 ? T93 : 1'h0;
  assign T93 = T95 | T94;
  assign T94 = io_tl_acquire_valid & acq_has_data;
  assign T95 = io_tl_release_valid & rel_has_data;
  assign T96 = T97 & data_from_rel;
  assign T97 = active_out & T98;
  assign T98 = has_data & T99;
  assign T99 = tl_done_out ^ 1'h1;
  assign T100 = T97 & T101;
  assign T101 = data_from_rel ^ 1'h1;
  assign io_mem_req_cmd_bits_rw = T102;
  assign T102 = T74 ? acq_has_data : T103;
  assign T103 = T74 ? acq_has_data : T104;
  assign T104 = T25 ? rel_has_data : has_data;
  assign io_mem_req_cmd_bits_tag = T105;
  assign T105 = T74 ? T134 : T106;
  assign T106 = T25 ? T133 : tag_out;
  assign T133 = {1'h0, T23};
  assign T134 = {1'h0, T72};
  assign io_mem_req_cmd_bits_addr = T107;
  assign T107 = T74 ? io_tl_acquire_bits_addr_block : T108;
  assign T108 = T25 ? io_tl_release_bits_addr_block : addr_out;
  assign T109 = T74 ? io_tl_acquire_bits_addr_block : T110;
  assign T110 = T25 ? io_tl_release_bits_addr_block : addr_out;
  assign io_mem_req_cmd_valid = T111;
  assign T111 = active_out ? T112 : T26;
  assign T112 = cmd_sent_out ^ 1'h1;
  assign io_tl_release_ready = T113;
  assign T113 = T96 ? io_mem_req_data_ready : T114;
  assign T114 = T29 ? io_mem_req_data_ready : 1'h0;
  assign io_tl_probe_valid = 1'h0;
  assign io_tl_finish_ready = 1'h1;
  assign io_tl_grant_bits_client_id = gnt_arb_io_out_bits_client_id;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_acquire_ready = T115;
  assign T115 = T100 ? io_mem_req_data_ready : T116;
  assign T116 = T29 ? T117 : 1'h0;
  assign T117 = io_mem_req_data_ready & T118;
  assign T118 = io_tl_release_valid ^ 1'h1;
  Arbiter_8 gnt_arb(
       .io_in_1_ready( gnt_arb_io_in_1_ready ),
       .io_in_1_valid( T46 ),
       .io_in_1_bits_addr_beat( T86 ),
       .io_in_1_bits_data( T85 ),
       .io_in_1_bits_client_xact_id( T83 ),
       .io_in_1_bits_manager_xact_id( T82 ),
       .io_in_1_bits_is_builtin_type( T81 ),
       .io_in_1_bits_g_type( T77 ),
       .io_in_1_bits_client_id( T19 ),
       .io_in_0_ready( gnt_arb_io_in_0_ready ),
       .io_in_0_valid( io_mem_resp_valid ),
       .io_in_0_bits_addr_beat( T11 ),
       .io_in_0_bits_data( T10 ),
       .io_in_0_bits_client_xact_id( T8 ),
       .io_in_0_bits_manager_xact_id( T7 ),
       .io_in_0_bits_is_builtin_type( T5 ),
       .io_in_0_bits_g_type( T2 ),
       .io_in_0_bits_client_id( T0 ),
       .io_out_ready( io_tl_grant_ready ),
       .io_out_valid( gnt_arb_io_out_valid ),
       .io_out_bits_addr_beat( gnt_arb_io_out_bits_addr_beat ),
       .io_out_bits_data( gnt_arb_io_out_bits_data ),
       .io_out_bits_client_xact_id( gnt_arb_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( gnt_arb_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( gnt_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( gnt_arb_io_out_bits_g_type ),
       .io_out_bits_client_id( gnt_arb_io_out_bits_client_id )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_in <= 2'h0;
    end else if(T14) begin
      tl_cnt_in <= T13;
    end
    if(T74) begin
      tag_out <= T129;
    end else if(T25) begin
      tag_out <= T122;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T34) begin
      active_out <= 1'h0;
    end else if(T26) begin
      active_out <= T32;
    end
    if(reset) begin
      make_grant_ack <= 1'h0;
    end else if(T45) begin
      make_grant_ack <= 1'h0;
    end else if(T74) begin
      make_grant_ack <= acq_has_data;
    end else if(T25) begin
      make_grant_ack <= 1'h1;
    end
    if(reset) begin
      tl_done_out <= 1'h0;
    end else if(T62) begin
      tl_done_out <= 1'h1;
    end else if(T26) begin
      tl_done_out <= tl_wrap_out;
    end
    if(reset) begin
      tl_cnt_out <= 2'h0;
    end else if(T53) begin
      tl_cnt_out <= T52;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T74) begin
      has_data <= acq_has_data;
    end else if(T25) begin
      has_data <= rel_has_data;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(active_out) begin
      cmd_sent_out <= T70;
    end else if(T26) begin
      cmd_sent_out <= io_mem_req_cmd_ready;
    end
    if(reset) begin
      data_from_rel <= 1'h0;
    end else if(T74) begin
      data_from_rel <= 1'h0;
    end else if(T25) begin
      data_from_rel <= 1'h1;
    end
    if(T74) begin
      addr_out <= io_tl_acquire_bits_addr_block;
    end else if(T25) begin
      addr_out <= io_tl_release_bits_addr_block;
    end
  end
endmodule

module HellaFlowQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
    //output[4:0] io_count
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[127:0] T2;
  wire ren;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire atLeastTwo;
  wire T30;
  wire[4:0] T31;
  reg [4:0] deq_ptr;
  wire[4:0] T37;
  wire[4:0] T18;
  wire[4:0] T19;
  wire[4:0] T20;
  wire T21;
  wire do_deq;
  wire T22;
  wire do_flow;
  wire T10;
  wire T23;
  reg [4:0] enq_ptr;
  wire[4:0] T38;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire T15;
  wire do_enq;
  wire T9;
  wire T11;
  wire full;
  reg  maybe_full;
  wire T39;
  wire T32;
  wire T33;
  wire ptr_match;
  wire[4:0] raddr;
  wire[4:0] T24;
  wire[4:0] T25;
  wire deq_done;
  wire[127:0] T4;
  wire[127:0] T5;
  wire T6;
  wire T7;
  wire[4:0] T8;
  reg [4:0] R16;
  wire[4:0] T17;
  wire empty;
  wire T34;
  wire T35;
  reg  ram_out_valid;
  wire T36;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    R16 = {1{$random}};
    ram_out_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_count = {1{$random}};
// synthesis translate_on
`endif
  assign io_deq_bits_data = T0;
  assign T0 = empty ? io_enq_bits_data : T1;
  assign T1 = T2[7'h7f:1'h0];
  assign ren = io_deq_ready & T26;
  assign T26 = atLeastTwo | T27;
  assign T27 = T29 & T28;
  assign T28 = empty ^ 1'h1;
  assign T29 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T30;
  assign T30 = 5'h2 <= T31;
  assign T31 = enq_ptr - deq_ptr;
  assign T37 = reset ? 5'h0 : T18;
  assign T18 = do_deq ? T19 : deq_ptr;
  assign T19 = T21 ? 5'h0 : T20;
  assign T20 = deq_ptr + 5'h1;
  assign T21 = deq_ptr == 5'h17;
  assign do_deq = T23 & T22;
  assign T22 = do_flow ^ 1'h1;
  assign do_flow = T10;
  assign T10 = empty & io_deq_ready;
  assign T23 = io_deq_ready & io_deq_valid;
  assign T38 = reset ? 5'h0 : T12;
  assign T12 = do_enq ? T13 : enq_ptr;
  assign T13 = T15 ? 5'h0 : T14;
  assign T14 = enq_ptr + 5'h1;
  assign T15 = enq_ptr == 5'h17;
  assign do_enq = T11 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T11 = io_enq_ready & io_enq_valid;
  assign full = ptr_match & maybe_full;
  assign T39 = reset ? 1'h0 : T32;
  assign T32 = T33 ? do_enq : maybe_full;
  assign T33 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign raddr = io_deq_valid ? T24 : deq_ptr;
  assign T24 = deq_done ? 5'h0 : T25;
  assign T25 = deq_ptr + 5'h1;
  assign deq_done = do_deq & T21;
  HellaFlowQueue_T3 T3 (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(T6),
    .W0I(T5),
    .R1A(raddr),
    .R1E(ren),
    .R1O(T2)
  );
  assign T5 = io_enq_bits_data;
  assign T6 = do_enq & T7;
  assign T7 = T8 < 5'h18;
  assign T8 = enq_ptr[3'h4:1'h0];
  assign T17 = ren ? raddr : R16;
  assign empty = ptr_match & T34;
  assign T34 = maybe_full ^ 1'h1;
  assign io_deq_valid = T35;
  assign T35 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 5'h0;
    end else if(do_deq) begin
      deq_ptr <= T19;
    end
    if(reset) begin
      enq_ptr <= 5'h0;
    end else if(do_enq) begin
      enq_ptr <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T33) begin
      maybe_full <= do_enq;
    end
    if(ren) begin
      R16 <= raddr;
    end
    ram_out_valid <= ren;
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output io_count
);

  wire T9;
  wire[1:0] T0;
  reg  full;
  wire T10;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[127:0] T4;
  reg [127:0] ram [0:0];
  wire[127:0] T5;
  wire T6;
  wire empty;
  wire T7;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T9;
  assign T9 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T10 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_data = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T7;
  assign T7 = T8 | io_deq_ready;
  assign T8 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= io_enq_bits_data;
  end
endmodule

module HellaQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
    //output[4:0] io_count
);

  wire fq_io_enq_ready;
  wire fq_io_deq_valid;
  wire[127:0] fq_io_deq_bits_data;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[127:0] Queue_io_deq_bits_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_count = {1{$random}};
// synthesis translate_on
`endif
  assign io_deq_bits_data = Queue_io_deq_bits_data;
  assign io_deq_valid = Queue_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue_0 fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_data( io_enq_bits_data ),
       .io_deq_ready( Queue_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_data( fq_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_12 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_data( fq_io_deq_bits_data ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
endmodule

module HellaFlowQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [5:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[5:0] io_deq_bits_tag
    //output[4:0] io_count
);

  wire[5:0] T0;
  wire[5:0] T1;
  wire[5:0] T2;
  wire ren;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire atLeastTwo;
  wire T30;
  wire[4:0] T31;
  reg [4:0] deq_ptr;
  wire[4:0] T37;
  wire[4:0] T18;
  wire[4:0] T19;
  wire[4:0] T20;
  wire T21;
  wire do_deq;
  wire T22;
  wire do_flow;
  wire T10;
  wire T23;
  reg [4:0] enq_ptr;
  wire[4:0] T38;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire T15;
  wire do_enq;
  wire T9;
  wire T11;
  wire full;
  reg  maybe_full;
  wire T39;
  wire T32;
  wire T33;
  wire ptr_match;
  wire[4:0] raddr;
  wire[4:0] T24;
  wire[4:0] T25;
  wire deq_done;
  wire[5:0] T4;
  wire[5:0] T5;
  wire T6;
  wire T7;
  wire[4:0] T8;
  reg [4:0] R16;
  wire[4:0] T17;
  wire empty;
  wire T34;
  wire T35;
  reg  ram_out_valid;
  wire T36;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    maybe_full = {1{$random}};
    R16 = {1{$random}};
    ram_out_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_count = {1{$random}};
// synthesis translate_on
`endif
  assign io_deq_bits_tag = T0;
  assign T0 = empty ? io_enq_bits_tag : T1;
  assign T1 = T2[3'h5:1'h0];
  assign ren = io_deq_ready & T26;
  assign T26 = atLeastTwo | T27;
  assign T27 = T29 & T28;
  assign T28 = empty ^ 1'h1;
  assign T29 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T30;
  assign T30 = 5'h2 <= T31;
  assign T31 = enq_ptr - deq_ptr;
  assign T37 = reset ? 5'h0 : T18;
  assign T18 = do_deq ? T19 : deq_ptr;
  assign T19 = T21 ? 5'h0 : T20;
  assign T20 = deq_ptr + 5'h1;
  assign T21 = deq_ptr == 5'h17;
  assign do_deq = T23 & T22;
  assign T22 = do_flow ^ 1'h1;
  assign do_flow = T10;
  assign T10 = empty & io_deq_ready;
  assign T23 = io_deq_ready & io_deq_valid;
  assign T38 = reset ? 5'h0 : T12;
  assign T12 = do_enq ? T13 : enq_ptr;
  assign T13 = T15 ? 5'h0 : T14;
  assign T14 = enq_ptr + 5'h1;
  assign T15 = enq_ptr == 5'h17;
  assign do_enq = T11 & T9;
  assign T9 = do_flow ^ 1'h1;
  assign T11 = io_enq_ready & io_enq_valid;
  assign full = ptr_match & maybe_full;
  assign T39 = reset ? 1'h0 : T32;
  assign T32 = T33 ? do_enq : maybe_full;
  assign T33 = do_enq != do_deq;
  assign ptr_match = enq_ptr == deq_ptr;
  assign raddr = io_deq_valid ? T24 : deq_ptr;
  assign T24 = deq_done ? 5'h0 : T25;
  assign T25 = deq_ptr + 5'h1;
  assign deq_done = do_deq & T21;
  HellaFlowQueue_T3_1 T3 (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(T6),
    .W0I(T5),
    .R1A(raddr),
    .R1E(ren),
    .R1O(T2)
  );
  assign T5 = io_enq_bits_tag;
  assign T6 = do_enq & T7;
  assign T7 = T8 < 5'h18;
  assign T8 = enq_ptr[3'h4:1'h0];
  assign T17 = ren ? raddr : R16;
  assign empty = ptr_match & T34;
  assign T34 = maybe_full ^ 1'h1;
  assign io_deq_valid = T35;
  assign T35 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      deq_ptr <= 5'h0;
    end else if(do_deq) begin
      deq_ptr <= T19;
    end
    if(reset) begin
      enq_ptr <= 5'h0;
    end else if(do_enq) begin
      enq_ptr <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T33) begin
      maybe_full <= do_enq;
    end
    if(ren) begin
      R16 <= raddr;
    end
    ram_out_valid <= ren;
  end
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [5:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[5:0] io_deq_bits_tag,
    output io_count
);

  wire T9;
  wire[1:0] T0;
  reg  full;
  wire T10;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[5:0] T3;
  wire[5:0] T4;
  reg [5:0] ram [0:0];
  wire[5:0] T5;
  wire T6;
  wire empty;
  wire T7;
  wire T8;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T9;
  assign T9 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T10 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_tag = T3;
  assign T3 = T4[3'h5:1'h0];
  assign T4 = ram[1'h0];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T7;
  assign T7 = T8 | io_deq_ready;
  assign T8 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= io_enq_bits_tag;
  end
endmodule

module HellaQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [5:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[5:0] io_deq_bits_tag
    //output[4:0] io_count
);

  wire fq_io_enq_ready;
  wire fq_io_deq_valid;
  wire[5:0] fq_io_deq_bits_tag;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[5:0] Queue_io_deq_bits_tag;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_count = {1{$random}};
// synthesis translate_on
`endif
  assign io_deq_bits_tag = Queue_io_deq_bits_tag;
  assign io_deq_valid = Queue_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue_1 fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_tag( io_enq_bits_tag ),
       .io_deq_ready( Queue_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_tag( fq_io_deq_bits_tag )
       //.io_count(  )
  );
  Queue_13 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_tag( fq_io_deq_bits_tag ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_tag( Queue_io_deq_bits_tag )
       //.io_count(  )
  );
endmodule

module MemPipeIOMemIOConverter(input clk, input reset,
    output io_cpu_req_cmd_ready,
    input  io_cpu_req_cmd_valid,
    input [25:0] io_cpu_req_cmd_bits_addr,
    input [5:0] io_cpu_req_cmd_bits_tag,
    input  io_cpu_req_cmd_bits_rw,
    output io_cpu_req_data_ready,
    input  io_cpu_req_data_valid,
    input [127:0] io_cpu_req_data_bits_data,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[127:0] io_cpu_resp_bits_data,
    output[5:0] io_cpu_resp_bits_tag,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[5:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [5:0] io_mem_resp_bits_tag
);

  wire T0;
  wire cmdq_mask;
  wire watermark;
  reg [4:0] count;
  wire[4:0] T20;
  wire[4:0] T1;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire T5;
  wire T6;
  wire dec;
  wire T7;
  wire T8;
  wire T9;
  wire inc;
  wire T10;
  wire T11;
  wire T12;
  wire[4:0] T13;
  wire T14;
  wire T15;
  wire[4:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire resp_data_q_io_deq_valid;
  wire[127:0] resp_data_q_io_deq_bits_data;
  wire resp_tag_q_io_deq_valid;
  wire[5:0] resp_tag_q_io_deq_bits_tag;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    count = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_mem_req_data_bits_data = io_cpu_req_data_bits_data;
  assign io_mem_req_data_valid = io_cpu_req_data_valid;
  assign io_mem_req_cmd_bits_rw = io_cpu_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = io_cpu_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = io_cpu_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = T0;
  assign T0 = io_cpu_req_cmd_valid & cmdq_mask;
  assign cmdq_mask = io_cpu_req_cmd_bits_rw | watermark;
  assign watermark = 5'h4 <= count;
  assign T20 = reset ? 5'h18 : T1;
  assign T1 = T17 ? T16 : T2;
  assign T2 = T14 ? T13 : T3;
  assign T3 = T5 ? T4 : count;
  assign T4 = count + 5'h1;
  assign T5 = inc & T6;
  assign T6 = dec ^ 1'h1;
  assign dec = T7;
  assign T7 = T9 & T8;
  assign T8 = io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T9 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign inc = T10;
  assign T10 = T12 & T11;
  assign T11 = io_cpu_resp_ready & resp_tag_q_io_deq_valid;
  assign T12 = io_cpu_resp_ready & resp_data_q_io_deq_valid;
  assign T13 = count - 5'h4;
  assign T14 = T15 & dec;
  assign T15 = inc ^ 1'h1;
  assign T16 = count - 5'h3;
  assign T17 = inc & dec;
  assign io_cpu_resp_bits_tag = resp_tag_q_io_deq_bits_tag;
  assign io_cpu_resp_bits_data = resp_data_q_io_deq_bits_data;
  assign io_cpu_resp_valid = T18;
  assign T18 = resp_data_q_io_deq_valid & resp_tag_q_io_deq_valid;
  assign io_cpu_req_data_ready = io_mem_req_data_ready;
  assign io_cpu_req_cmd_ready = T19;
  assign T19 = io_mem_req_cmd_ready & cmdq_mask;
  HellaQueue_0 resp_data_q(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_data_q_io_deq_valid ),
       .io_deq_bits_data( resp_data_q_io_deq_bits_data )
       //.io_count(  )
  );
  HellaQueue_1 resp_tag_q(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_tag_q_io_deq_valid ),
       .io_deq_bits_tag( resp_tag_q_io_deq_bits_tag )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      count <= 5'h18;
    end else if(T17) begin
      count <= T16;
    end else if(T14) begin
      count <= T13;
    end else if(T5) begin
      count <= T4;
    end
  end
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [5:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[5:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T22;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T23;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T24;
  wire T8;
  wire T9;
  wire T10;
  wire[32:0] T11;
  reg [32:0] ram [1:0];
  wire[32:0] T12;
  wire[32:0] T13;
  wire[32:0] T14;
  wire[6:0] T15;
  wire[5:0] T16;
  wire[25:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire T21;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T22 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T23 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T24 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_rw = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_addr, T15};
  assign T15 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T16;
  assign T16 = T11[3'h6:1'h1];
  assign io_deq_bits_addr = T17;
  assign T17 = T11[6'h20:3'h7];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = T21 | io_deq_ready;
  assign T21 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[2:0] io_count
);

  wire[2:0] T0;
  wire[1:0] ptr_diff;
  reg [1:0] R1;
  wire[1:0] T17;
  wire[1:0] T2;
  wire[1:0] T3;
  wire do_deq;
  reg [1:0] R4;
  wire[1:0] T18;
  wire[1:0] T5;
  wire[1:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T19;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[127:0] T11;
  reg [127:0] ram [3:0];
  wire[127:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire T16;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T17 = reset ? 2'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T18 = reset ? 2'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 2'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T19 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = T16 | io_deq_ready;
  assign T16 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 2'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 2'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_data;
  end
endmodule

module MemPipeIOTileLinkIOConverter(input clk, input reset,
    output io_tl_acquire_ready,
    input  io_tl_acquire_valid,
    input [25:0] io_tl_acquire_bits_addr_block,
    input [2:0] io_tl_acquire_bits_client_xact_id,
    input [1:0] io_tl_acquire_bits_addr_beat,
    input [127:0] io_tl_acquire_bits_data,
    input  io_tl_acquire_bits_is_builtin_type,
    input [2:0] io_tl_acquire_bits_a_type,
    input [16:0] io_tl_acquire_bits_union,
    input  io_tl_acquire_bits_client_id,
    input  io_tl_grant_ready,
    output io_tl_grant_valid,
    output[1:0] io_tl_grant_bits_addr_beat,
    output[127:0] io_tl_grant_bits_data,
    output[2:0] io_tl_grant_bits_client_xact_id,
    output io_tl_grant_bits_manager_xact_id,
    output io_tl_grant_bits_is_builtin_type,
    output[3:0] io_tl_grant_bits_g_type,
    output io_tl_grant_bits_client_id,
    output io_tl_finish_ready,
    input  io_tl_finish_valid,
    input  io_tl_finish_bits_manager_xact_id,
    input  io_tl_probe_ready,
    output io_tl_probe_valid,
    //output[25:0] io_tl_probe_bits_addr_block
    //output[1:0] io_tl_probe_bits_p_type
    //output io_tl_probe_bits_client_id
    output io_tl_release_ready,
    input  io_tl_release_valid,
    input [25:0] io_tl_release_bits_addr_block,
    input [2:0] io_tl_release_bits_client_xact_id,
    input [1:0] io_tl_release_bits_addr_beat,
    input [127:0] io_tl_release_bits_data,
    input [2:0] io_tl_release_bits_r_type,
    input  io_tl_release_bits_voluntary,
    input  io_tl_release_bits_client_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[5:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [5:0] io_mem_resp_bits_tag
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[25:0] Queue_io_deq_bits_addr;
  wire[5:0] Queue_io_deq_bits_tag;
  wire Queue_io_deq_bits_rw;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[127:0] Queue_1_io_deq_bits_data;
  wire a_io_tl_acquire_ready;
  wire a_io_tl_grant_valid;
  wire[1:0] a_io_tl_grant_bits_addr_beat;
  wire[127:0] a_io_tl_grant_bits_data;
  wire[2:0] a_io_tl_grant_bits_client_xact_id;
  wire a_io_tl_grant_bits_manager_xact_id;
  wire a_io_tl_grant_bits_is_builtin_type;
  wire[3:0] a_io_tl_grant_bits_g_type;
  wire a_io_tl_grant_bits_client_id;
  wire a_io_tl_finish_ready;
  wire a_io_tl_probe_valid;
  wire a_io_tl_release_ready;
  wire a_io_mem_req_cmd_valid;
  wire[25:0] a_io_mem_req_cmd_bits_addr;
  wire[5:0] a_io_mem_req_cmd_bits_tag;
  wire a_io_mem_req_cmd_bits_rw;
  wire a_io_mem_req_data_valid;
  wire[127:0] a_io_mem_req_data_bits_data;
  wire a_io_mem_resp_ready;
  wire b_io_cpu_req_cmd_ready;
  wire b_io_cpu_req_data_ready;
  wire b_io_cpu_resp_valid;
  wire[127:0] b_io_cpu_resp_bits_data;
  wire[5:0] b_io_cpu_resp_bits_tag;
  wire b_io_mem_req_cmd_valid;
  wire[25:0] b_io_mem_req_cmd_bits_addr;
  wire[5:0] b_io_mem_req_cmd_bits_tag;
  wire b_io_mem_req_cmd_bits_rw;
  wire b_io_mem_req_data_valid;
  wire[127:0] b_io_mem_req_data_bits_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_tl_probe_bits_client_id = {1{$random}};
//  assign io_tl_probe_bits_p_type = {1{$random}};
//  assign io_tl_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_req_data_bits_data = b_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = b_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = b_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = b_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = b_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = b_io_mem_req_cmd_valid;
  assign io_tl_release_ready = a_io_tl_release_ready;
  assign io_tl_probe_valid = a_io_tl_probe_valid;
  assign io_tl_finish_ready = a_io_tl_finish_ready;
  assign io_tl_grant_bits_client_id = a_io_tl_grant_bits_client_id;
  assign io_tl_grant_bits_g_type = a_io_tl_grant_bits_g_type;
  assign io_tl_grant_bits_is_builtin_type = a_io_tl_grant_bits_is_builtin_type;
  assign io_tl_grant_bits_manager_xact_id = a_io_tl_grant_bits_manager_xact_id;
  assign io_tl_grant_bits_client_xact_id = a_io_tl_grant_bits_client_xact_id;
  assign io_tl_grant_bits_data = a_io_tl_grant_bits_data;
  assign io_tl_grant_bits_addr_beat = a_io_tl_grant_bits_addr_beat;
  assign io_tl_grant_valid = a_io_tl_grant_valid;
  assign io_tl_acquire_ready = a_io_tl_acquire_ready;
  MemIOTileLinkIOConverter a(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( a_io_tl_acquire_ready ),
       .io_tl_acquire_valid( io_tl_acquire_valid ),
       .io_tl_acquire_bits_addr_block( io_tl_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( io_tl_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( io_tl_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_data( io_tl_acquire_bits_data ),
       .io_tl_acquire_bits_is_builtin_type( io_tl_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( io_tl_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( io_tl_acquire_bits_union ),
       .io_tl_acquire_bits_client_id( io_tl_acquire_bits_client_id ),
       .io_tl_grant_ready( io_tl_grant_ready ),
       .io_tl_grant_valid( a_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( a_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_data( a_io_tl_grant_bits_data ),
       .io_tl_grant_bits_client_xact_id( a_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( a_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( a_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( a_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_client_id( a_io_tl_grant_bits_client_id ),
       .io_tl_finish_ready( a_io_tl_finish_ready ),
       .io_tl_finish_valid( io_tl_finish_valid ),
       .io_tl_finish_bits_manager_xact_id( io_tl_finish_bits_manager_xact_id ),
       .io_tl_probe_ready( io_tl_probe_ready ),
       .io_tl_probe_valid( a_io_tl_probe_valid ),
       //.io_tl_probe_bits_addr_block(  )
       //.io_tl_probe_bits_p_type(  )
       //.io_tl_probe_bits_client_id(  )
       .io_tl_release_ready( a_io_tl_release_ready ),
       .io_tl_release_valid( io_tl_release_valid ),
       .io_tl_release_bits_addr_block( io_tl_release_bits_addr_block ),
       .io_tl_release_bits_client_xact_id( io_tl_release_bits_client_xact_id ),
       .io_tl_release_bits_addr_beat( io_tl_release_bits_addr_beat ),
       .io_tl_release_bits_data( io_tl_release_bits_data ),
       .io_tl_release_bits_r_type( io_tl_release_bits_r_type ),
       .io_tl_release_bits_voluntary( io_tl_release_bits_voluntary ),
       .io_tl_release_bits_client_id( io_tl_release_bits_client_id ),
       .io_mem_req_cmd_ready( Queue_io_enq_ready ),
       .io_mem_req_cmd_valid( a_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_1_io_enq_ready ),
       .io_mem_req_data_valid( a_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( a_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( a_io_mem_resp_ready ),
       .io_mem_resp_valid( b_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_tag( b_io_cpu_resp_bits_tag )
  );
  MemPipeIOMemIOConverter b(.clk(clk), .reset(reset),
       .io_cpu_req_cmd_ready( b_io_cpu_req_cmd_ready ),
       .io_cpu_req_cmd_valid( Queue_io_deq_valid ),
       .io_cpu_req_cmd_bits_addr( Queue_io_deq_bits_addr ),
       .io_cpu_req_cmd_bits_tag( Queue_io_deq_bits_tag ),
       .io_cpu_req_cmd_bits_rw( Queue_io_deq_bits_rw ),
       .io_cpu_req_data_ready( b_io_cpu_req_data_ready ),
       .io_cpu_req_data_valid( Queue_1_io_deq_valid ),
       .io_cpu_req_data_bits_data( Queue_1_io_deq_bits_data ),
       .io_cpu_resp_ready( a_io_mem_resp_ready ),
       .io_cpu_resp_valid( b_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( b_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_tag( b_io_cpu_resp_bits_tag ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( b_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( b_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( b_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( b_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( b_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( b_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_3 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( a_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( a_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( a_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( b_io_cpu_req_cmd_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_4 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( a_io_mem_req_data_valid ),
       .io_enq_bits_data( a_io_mem_req_data_bits_data ),
       .io_deq_ready( b_io_cpu_req_data_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_data( Queue_1_io_deq_bits_data )
       //.io_count(  )
  );
endmodule

module ClientTileLinkIOWrapper_1(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [2:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[127:0] io_in_grant_bits_data,
    output[2:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output[127:0] io_out_acquire_bits_data,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [127:0] io_out_grant_bits_data,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[25:0] io_out_release_bits_addr_block
    //output[2:0] io_out_release_bits_client_xact_id
    //output[1:0] io_out_release_bits_addr_beat
    //output[127:0] io_out_release_bits_data
    //output[2:0] io_out_release_bits_r_type
    //output io_out_release_bits_voluntary
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input  io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    output io_tiles_cached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input  io_tiles_cached_0_release_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [127:0] io_tiles_cached_0_release_bits_data,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input  io_tiles_cached_0_release_bits_voluntary,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input  io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_tiles_uncached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output io_htif_uncached_acquire_ready,
    input  io_htif_uncached_acquire_valid,
    input [25:0] io_htif_uncached_acquire_bits_addr_block,
    input  io_htif_uncached_acquire_bits_client_xact_id,
    input [1:0] io_htif_uncached_acquire_bits_addr_beat,
    input [127:0] io_htif_uncached_acquire_bits_data,
    input  io_htif_uncached_acquire_bits_is_builtin_type,
    input [2:0] io_htif_uncached_acquire_bits_a_type,
    input [16:0] io_htif_uncached_acquire_bits_union,
    input  io_htif_uncached_grant_ready,
    output io_htif_uncached_grant_valid,
    output[1:0] io_htif_uncached_grant_bits_addr_beat,
    output[127:0] io_htif_uncached_grant_bits_data,
    output io_htif_uncached_grant_bits_client_xact_id,
    output[2:0] io_htif_uncached_grant_bits_manager_xact_id,
    output io_htif_uncached_grant_bits_is_builtin_type,
    output[3:0] io_htif_uncached_grant_bits_g_type,
    input  io_incoherent_0,
    input  io_mem_0_req_cmd_ready,
    output io_mem_0_req_cmd_valid,
    output[25:0] io_mem_0_req_cmd_bits_addr,
    output[5:0] io_mem_0_req_cmd_bits_tag,
    output io_mem_0_req_cmd_bits_rw,
    input  io_mem_0_req_data_ready,
    output io_mem_0_req_data_valid,
    output[127:0] io_mem_0_req_data_bits_data,
    output io_mem_0_resp_ready,
    input  io_mem_0_resp_valid,
    input [127:0] io_mem_0_resp_bits_data,
    input [5:0] io_mem_0_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire[5:0] T0;
  wire[127:0] T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[127:0] T6;
  wire T7;
  wire T8;
  wire[5:0] T9;
  wire[25:0] T10;
  wire T11;
  wire ClientTileLinkIOWrapper_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  wire ClientTileLinkIOWrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block;
  wire ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_io_out_acquire_bits_union;
  wire ClientTileLinkIOWrapper_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_io_out_release_valid;
  wire ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_1_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_union;
  wire ClientTileLinkIOWrapper_1_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_1_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_1_io_out_release_valid;
  wire ClientTileLinkIOWrapper_2_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_2_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_data;
  wire[2:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat;
  wire[127:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_union;
  wire ClientTileLinkIOWrapper_2_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_2_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_2_io_out_release_valid;
  wire L2BroadcastHub_io_inner_acquire_ready;
  wire L2BroadcastHub_io_inner_grant_valid;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_addr_beat;
  wire[127:0] L2BroadcastHub_io_inner_grant_bits_data;
  wire L2BroadcastHub_io_inner_grant_bits_client_xact_id;
  wire[2:0] L2BroadcastHub_io_inner_grant_bits_manager_xact_id;
  wire L2BroadcastHub_io_inner_grant_bits_is_builtin_type;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_g_type;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_id;
  wire L2BroadcastHub_io_inner_finish_ready;
  wire L2BroadcastHub_io_inner_probe_valid;
  wire[25:0] L2BroadcastHub_io_inner_probe_bits_addr_block;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_p_type;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_client_id;
  wire L2BroadcastHub_io_inner_release_ready;
  wire L2BroadcastHub_io_outer_acquire_valid;
  wire[25:0] L2BroadcastHub_io_outer_acquire_bits_addr_block;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_client_xact_id;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_addr_beat;
  wire[127:0] L2BroadcastHub_io_outer_acquire_bits_data;
  wire L2BroadcastHub_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_a_type;
  wire[16:0] L2BroadcastHub_io_outer_acquire_bits_union;
  wire L2BroadcastHub_io_outer_grant_ready;
  wire l1tol2net_io_clients_2_acquire_ready;
  wire l1tol2net_io_clients_2_grant_valid;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_addr_beat;
  wire[127:0] l1tol2net_io_clients_2_grant_bits_data;
  wire l1tol2net_io_clients_2_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_2_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_2_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_g_type;
  wire l1tol2net_io_clients_2_probe_valid;
  wire[25:0] l1tol2net_io_clients_2_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_2_probe_bits_p_type;
  wire l1tol2net_io_clients_2_release_ready;
  wire l1tol2net_io_clients_1_acquire_ready;
  wire l1tol2net_io_clients_1_grant_valid;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_addr_beat;
  wire[127:0] l1tol2net_io_clients_1_grant_bits_data;
  wire l1tol2net_io_clients_1_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_1_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_1_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_g_type;
  wire l1tol2net_io_clients_1_probe_valid;
  wire[25:0] l1tol2net_io_clients_1_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_1_probe_bits_p_type;
  wire l1tol2net_io_clients_1_release_ready;
  wire l1tol2net_io_clients_0_acquire_ready;
  wire l1tol2net_io_clients_0_grant_valid;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_addr_beat;
  wire[127:0] l1tol2net_io_clients_0_grant_bits_data;
  wire l1tol2net_io_clients_0_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_g_type;
  wire l1tol2net_io_clients_0_probe_valid;
  wire[25:0] l1tol2net_io_clients_0_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_0_probe_bits_p_type;
  wire l1tol2net_io_clients_0_release_ready;
  wire l1tol2net_io_managers_0_acquire_valid;
  wire[25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire[127:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire[2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire[16:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_id;
  wire l1tol2net_io_managers_0_grant_ready;
  wire l1tol2net_io_managers_0_finish_valid;
  wire[2:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire l1tol2net_io_managers_0_probe_ready;
  wire l1tol2net_io_managers_0_release_valid;
  wire[25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire[127:0] l1tol2net_io_managers_0_release_bits_data;
  wire[2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire l1tol2net_io_managers_0_release_bits_voluntary;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_id;
  wire RocketChipTileLinkArbiter_io_clients_0_acquire_ready;
  wire RocketChipTileLinkArbiter_io_clients_0_grant_valid;
  wire[1:0] RocketChipTileLinkArbiter_io_clients_0_grant_bits_addr_beat;
  wire[127:0] RocketChipTileLinkArbiter_io_clients_0_grant_bits_data;
  wire[2:0] RocketChipTileLinkArbiter_io_clients_0_grant_bits_client_xact_id;
  wire RocketChipTileLinkArbiter_io_clients_0_grant_bits_manager_xact_id;
  wire RocketChipTileLinkArbiter_io_clients_0_grant_bits_is_builtin_type;
  wire[3:0] RocketChipTileLinkArbiter_io_clients_0_grant_bits_g_type;
  wire RocketChipTileLinkArbiter_io_clients_0_probe_valid;
  wire[25:0] RocketChipTileLinkArbiter_io_clients_0_probe_bits_addr_block;
  wire[1:0] RocketChipTileLinkArbiter_io_clients_0_probe_bits_p_type;
  wire RocketChipTileLinkArbiter_io_clients_0_release_ready;
  wire RocketChipTileLinkArbiter_io_managers_0_acquire_valid;
  wire[25:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_block;
  wire[2:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_xact_id;
  wire[1:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_beat;
  wire[127:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_data;
  wire RocketChipTileLinkArbiter_io_managers_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_a_type;
  wire[16:0] RocketChipTileLinkArbiter_io_managers_0_acquire_bits_union;
  wire RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_id;
  wire RocketChipTileLinkArbiter_io_managers_0_grant_ready;
  wire RocketChipTileLinkArbiter_io_managers_0_finish_valid;
  wire RocketChipTileLinkArbiter_io_managers_0_finish_bits_manager_xact_id;
  wire RocketChipTileLinkArbiter_io_managers_0_probe_ready;
  wire RocketChipTileLinkArbiter_io_managers_0_release_valid;
  wire[25:0] RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_block;
  wire[2:0] RocketChipTileLinkArbiter_io_managers_0_release_bits_client_xact_id;
  wire[1:0] RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_beat;
  wire[127:0] RocketChipTileLinkArbiter_io_managers_0_release_bits_data;
  wire[2:0] RocketChipTileLinkArbiter_io_managers_0_release_bits_r_type;
  wire RocketChipTileLinkArbiter_io_managers_0_release_bits_voluntary;
  wire RocketChipTileLinkArbiter_io_managers_0_release_bits_client_id;
  wire MemPipeIOTileLinkIOConverter_io_tl_acquire_ready;
  wire MemPipeIOTileLinkIOConverter_io_tl_grant_valid;
  wire[1:0] MemPipeIOTileLinkIOConverter_io_tl_grant_bits_addr_beat;
  wire[127:0] MemPipeIOTileLinkIOConverter_io_tl_grant_bits_data;
  wire[2:0] MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id;
  wire MemPipeIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id;
  wire MemPipeIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type;
  wire[3:0] MemPipeIOTileLinkIOConverter_io_tl_grant_bits_g_type;
  wire MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_id;
  wire MemPipeIOTileLinkIOConverter_io_tl_finish_ready;
  wire MemPipeIOTileLinkIOConverter_io_tl_probe_valid;
  wire MemPipeIOTileLinkIOConverter_io_tl_release_ready;
  wire MemPipeIOTileLinkIOConverter_io_mem_req_cmd_valid;
  wire[25:0] MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_addr;
  wire[5:0] MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_tag;
  wire MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_rw;
  wire MemPipeIOTileLinkIOConverter_io_mem_req_data_valid;
  wire[127:0] MemPipeIOTileLinkIOConverter_io_mem_req_data_bits_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_req_bits = {1{$random}};
//  assign io_mem_backup_req_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = io_mem_0_resp_bits_tag;
  assign T1 = io_mem_0_resp_bits_data;
  assign T2 = io_mem_0_resp_valid;
  assign T3 = io_mem_0_req_data_ready;
  assign T4 = io_mem_0_req_cmd_ready;
  assign io_mem_0_resp_ready = T5;
  assign T5 = 1'h1;
  assign io_mem_0_req_data_bits_data = T6;
  assign T6 = MemPipeIOTileLinkIOConverter_io_mem_req_data_bits_data;
  assign io_mem_0_req_data_valid = T7;
  assign T7 = MemPipeIOTileLinkIOConverter_io_mem_req_data_valid;
  assign io_mem_0_req_cmd_bits_rw = T8;
  assign T8 = MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_rw;
  assign io_mem_0_req_cmd_bits_tag = T9;
  assign T9 = MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_tag;
  assign io_mem_0_req_cmd_bits_addr = T10;
  assign T10 = MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_addr;
  assign io_mem_0_req_cmd_valid = T11;
  assign T11 = MemPipeIOTileLinkIOConverter_io_mem_req_cmd_valid;
  assign io_htif_uncached_grant_bits_g_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  assign io_htif_uncached_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  assign io_htif_uncached_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  assign io_htif_uncached_grant_bits_client_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  assign io_htif_uncached_grant_bits_data = ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  assign io_htif_uncached_grant_bits_addr_beat = ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  assign io_htif_uncached_grant_valid = ClientTileLinkIOWrapper_1_io_in_grant_valid;
  assign io_htif_uncached_acquire_ready = ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  assign io_tiles_uncached_0_grant_bits_g_type = ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_data = ClientTileLinkIOWrapper_io_in_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_addr_beat = ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = ClientTileLinkIOWrapper_io_in_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = ClientTileLinkIOWrapper_io_in_acquire_ready;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_0_acquire_ready;
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_in_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_in_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_in_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_io_in_grant_bits_data ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_io_in_grant_bits_g_type ),
       .io_out_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_out_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_io_out_release_valid )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_data(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
  );
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper_1(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_1_io_in_acquire_ready ),
       .io_in_acquire_valid( io_htif_uncached_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_htif_uncached_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_htif_uncached_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_htif_uncached_acquire_bits_addr_beat ),
       .io_in_acquire_bits_data( io_htif_uncached_acquire_bits_data ),
       .io_in_acquire_bits_is_builtin_type( io_htif_uncached_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_htif_uncached_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_htif_uncached_acquire_bits_union ),
       .io_in_grant_ready( io_htif_uncached_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_1_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_1_io_in_grant_bits_data ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type ),
       .io_out_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_out_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_data(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
  );
  RocketChipTileLinkArbiter_0 l1tol2net(.clk(clk), .reset(reset),
       .io_clients_2_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_clients_2_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_clients_2_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_clients_2_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_clients_2_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_clients_2_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_clients_2_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_clients_2_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_clients_2_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_clients_2_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_clients_2_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_clients_2_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_clients_2_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_clients_2_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_clients_2_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_clients_2_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_clients_2_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_clients_2_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_clients_2_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_clients_2_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_clients_2_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_clients_2_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_clients_2_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid ),
       //.io_clients_2_release_bits_addr_block(  )
       //.io_clients_2_release_bits_client_xact_id(  )
       //.io_clients_2_release_bits_addr_beat(  )
       //.io_clients_2_release_bits_data(  )
       //.io_clients_2_release_bits_r_type(  )
       //.io_clients_2_release_bits_voluntary(  )
       .io_clients_1_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_clients_1_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_clients_1_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_clients_1_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_clients_1_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_clients_1_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_clients_1_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_clients_1_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_clients_1_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_clients_1_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_clients_1_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_clients_1_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_clients_1_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_clients_1_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_clients_1_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_clients_1_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_clients_1_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_clients_1_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_clients_1_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( ClientTileLinkIOWrapper_io_out_release_valid ),
       //.io_clients_1_release_bits_addr_block(  )
       //.io_clients_1_release_bits_client_xact_id(  )
       //.io_clients_1_release_bits_addr_beat(  )
       //.io_clients_1_release_bits_data(  )
       //.io_clients_1_release_bits_r_type(  )
       //.io_clients_1_release_bits_voluntary(  )
       .io_clients_0_acquire_ready( l1tol2net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_clients_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_clients_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_clients_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_clients_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_clients_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_clients_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_clients_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_clients_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_clients_0_grant_valid( l1tol2net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_addr_beat( l1tol2net_io_clients_0_grant_bits_addr_beat ),
       .io_clients_0_grant_bits_data( l1tol2net_io_clients_0_grant_bits_data ),
       .io_clients_0_grant_bits_client_xact_id( l1tol2net_io_clients_0_grant_bits_client_xact_id ),
       .io_clients_0_grant_bits_manager_xact_id( l1tol2net_io_clients_0_grant_bits_manager_xact_id ),
       .io_clients_0_grant_bits_is_builtin_type( l1tol2net_io_clients_0_grant_bits_is_builtin_type ),
       .io_clients_0_grant_bits_g_type( l1tol2net_io_clients_0_grant_bits_g_type ),
       .io_clients_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_clients_0_probe_valid( l1tol2net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_addr_block( l1tol2net_io_clients_0_probe_bits_addr_block ),
       .io_clients_0_probe_bits_p_type( l1tol2net_io_clients_0_probe_bits_p_type ),
       .io_clients_0_release_ready( l1tol2net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_clients_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_clients_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_clients_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_clients_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_clients_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_clients_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_managers_0_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_managers_0_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_managers_0_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_managers_0_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_managers_0_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_managers_0_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_managers_0_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_managers_0_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_managers_0_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_managers_0_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_managers_0_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_managers_0_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_managers_0_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_managers_0_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_managers_0_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_managers_0_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_managers_0_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_managers_0_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_managers_0_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_managers_0_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_managers_0_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_managers_0_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_managers_0_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_managers_0_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_managers_0_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_managers_0_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_managers_0_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_managers_0_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_managers_0_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_managers_0_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_managers_0_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_managers_0_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign l1tol2net.io_clients_2_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_data = {4{$random}};
    assign l1tol2net.io_clients_2_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_data = {4{$random}};
    assign l1tol2net.io_clients_1_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_voluntary = {1{$random}};
// synthesis translate_on
`endif
  L2BroadcastHub L2BroadcastHub(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_inner_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_inner_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_inner_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_inner_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_inner_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_inner_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_inner_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_inner_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_inner_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_inner_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_inner_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_inner_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_inner_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_inner_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_inner_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_inner_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_outer_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_outer_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_outer_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type )
  );
  RocketChipTileLinkArbiter_1 RocketChipTileLinkArbiter(.clk(clk), .reset(reset),
       .io_clients_0_acquire_ready( RocketChipTileLinkArbiter_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_clients_0_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_clients_0_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_clients_0_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_clients_0_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_clients_0_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_clients_0_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_clients_0_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_clients_0_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_clients_0_grant_valid( RocketChipTileLinkArbiter_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_addr_beat( RocketChipTileLinkArbiter_io_clients_0_grant_bits_addr_beat ),
       .io_clients_0_grant_bits_data( RocketChipTileLinkArbiter_io_clients_0_grant_bits_data ),
       .io_clients_0_grant_bits_client_xact_id( RocketChipTileLinkArbiter_io_clients_0_grant_bits_client_xact_id ),
       .io_clients_0_grant_bits_manager_xact_id( RocketChipTileLinkArbiter_io_clients_0_grant_bits_manager_xact_id ),
       .io_clients_0_grant_bits_is_builtin_type( RocketChipTileLinkArbiter_io_clients_0_grant_bits_is_builtin_type ),
       .io_clients_0_grant_bits_g_type( RocketChipTileLinkArbiter_io_clients_0_grant_bits_g_type ),
       .io_clients_0_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_clients_0_probe_valid( RocketChipTileLinkArbiter_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_addr_block( RocketChipTileLinkArbiter_io_clients_0_probe_bits_addr_block ),
       .io_clients_0_probe_bits_p_type( RocketChipTileLinkArbiter_io_clients_0_probe_bits_p_type ),
       .io_clients_0_release_ready( RocketChipTileLinkArbiter_io_clients_0_release_ready ),
       .io_clients_0_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid ),
       //.io_clients_0_release_bits_addr_block(  )
       //.io_clients_0_release_bits_client_xact_id(  )
       //.io_clients_0_release_bits_addr_beat(  )
       //.io_clients_0_release_bits_data(  )
       //.io_clients_0_release_bits_r_type(  )
       //.io_clients_0_release_bits_voluntary(  )
       .io_managers_0_acquire_ready( MemPipeIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_managers_0_acquire_valid( RocketChipTileLinkArbiter_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_addr_block( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_block ),
       .io_managers_0_acquire_bits_client_xact_id( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_xact_id ),
       .io_managers_0_acquire_bits_addr_beat( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_beat ),
       .io_managers_0_acquire_bits_data( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_data ),
       .io_managers_0_acquire_bits_is_builtin_type( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_is_builtin_type ),
       .io_managers_0_acquire_bits_a_type( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_a_type ),
       .io_managers_0_acquire_bits_union( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_union ),
       .io_managers_0_acquire_bits_client_id( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_id ),
       .io_managers_0_grant_ready( RocketChipTileLinkArbiter_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( MemPipeIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_managers_0_grant_bits_addr_beat( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_managers_0_grant_bits_data( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_data ),
       .io_managers_0_grant_bits_client_xact_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_managers_0_grant_bits_manager_xact_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_managers_0_grant_bits_is_builtin_type( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_managers_0_grant_bits_g_type( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_managers_0_grant_bits_client_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_id ),
       .io_managers_0_finish_ready( MemPipeIOTileLinkIOConverter_io_tl_finish_ready ),
       .io_managers_0_finish_valid( RocketChipTileLinkArbiter_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_manager_xact_id( RocketChipTileLinkArbiter_io_managers_0_finish_bits_manager_xact_id ),
       .io_managers_0_probe_ready( RocketChipTileLinkArbiter_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( MemPipeIOTileLinkIOConverter_io_tl_probe_valid ),
       //.io_managers_0_probe_bits_addr_block(  )
       //.io_managers_0_probe_bits_p_type(  )
       //.io_managers_0_probe_bits_client_id(  )
       .io_managers_0_release_ready( MemPipeIOTileLinkIOConverter_io_tl_release_ready ),
       .io_managers_0_release_valid( RocketChipTileLinkArbiter_io_managers_0_release_valid ),
       .io_managers_0_release_bits_addr_block( RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_block ),
       .io_managers_0_release_bits_client_xact_id( RocketChipTileLinkArbiter_io_managers_0_release_bits_client_xact_id ),
       .io_managers_0_release_bits_addr_beat( RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_beat ),
       .io_managers_0_release_bits_data( RocketChipTileLinkArbiter_io_managers_0_release_bits_data ),
       .io_managers_0_release_bits_r_type( RocketChipTileLinkArbiter_io_managers_0_release_bits_r_type ),
       .io_managers_0_release_bits_voluntary( RocketChipTileLinkArbiter_io_managers_0_release_bits_voluntary ),
       .io_managers_0_release_bits_client_id( RocketChipTileLinkArbiter_io_managers_0_release_bits_client_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_addr_block = {1{$random}};
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_client_xact_id = {1{$random}};
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_addr_beat = {1{$random}};
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_data = {4{$random}};
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_r_type = {1{$random}};
    assign RocketChipTileLinkArbiter.io_clients_0_release_bits_voluntary = {1{$random}};
    assign RocketChipTileLinkArbiter.io_managers_0_probe_bits_addr_block = {1{$random}};
    assign RocketChipTileLinkArbiter.io_managers_0_probe_bits_p_type = {1{$random}};
    assign RocketChipTileLinkArbiter.io_managers_0_probe_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  MemPipeIOTileLinkIOConverter MemPipeIOTileLinkIOConverter(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( MemPipeIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_tl_acquire_valid( RocketChipTileLinkArbiter_io_managers_0_acquire_valid ),
       .io_tl_acquire_bits_addr_block( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_data( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_data ),
       .io_tl_acquire_bits_is_builtin_type( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_union ),
       .io_tl_acquire_bits_client_id( RocketChipTileLinkArbiter_io_managers_0_acquire_bits_client_id ),
       .io_tl_grant_ready( RocketChipTileLinkArbiter_io_managers_0_grant_ready ),
       .io_tl_grant_valid( MemPipeIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_data( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_data ),
       .io_tl_grant_bits_client_xact_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_client_id( MemPipeIOTileLinkIOConverter_io_tl_grant_bits_client_id ),
       .io_tl_finish_ready( MemPipeIOTileLinkIOConverter_io_tl_finish_ready ),
       .io_tl_finish_valid( RocketChipTileLinkArbiter_io_managers_0_finish_valid ),
       .io_tl_finish_bits_manager_xact_id( RocketChipTileLinkArbiter_io_managers_0_finish_bits_manager_xact_id ),
       .io_tl_probe_ready( RocketChipTileLinkArbiter_io_managers_0_probe_ready ),
       .io_tl_probe_valid( MemPipeIOTileLinkIOConverter_io_tl_probe_valid ),
       //.io_tl_probe_bits_addr_block(  )
       //.io_tl_probe_bits_p_type(  )
       //.io_tl_probe_bits_client_id(  )
       .io_tl_release_ready( MemPipeIOTileLinkIOConverter_io_tl_release_ready ),
       .io_tl_release_valid( RocketChipTileLinkArbiter_io_managers_0_release_valid ),
       .io_tl_release_bits_addr_block( RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_block ),
       .io_tl_release_bits_client_xact_id( RocketChipTileLinkArbiter_io_managers_0_release_bits_client_xact_id ),
       .io_tl_release_bits_addr_beat( RocketChipTileLinkArbiter_io_managers_0_release_bits_addr_beat ),
       .io_tl_release_bits_data( RocketChipTileLinkArbiter_io_managers_0_release_bits_data ),
       .io_tl_release_bits_r_type( RocketChipTileLinkArbiter_io_managers_0_release_bits_r_type ),
       .io_tl_release_bits_voluntary( RocketChipTileLinkArbiter_io_managers_0_release_bits_voluntary ),
       .io_tl_release_bits_client_id( RocketChipTileLinkArbiter_io_managers_0_release_bits_client_id ),
       .io_mem_req_cmd_ready( T4 ),
       .io_mem_req_cmd_valid( MemPipeIOTileLinkIOConverter_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( MemPipeIOTileLinkIOConverter_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( T3 ),
       .io_mem_req_data_valid( MemPipeIOTileLinkIOConverter_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( MemPipeIOTileLinkIOConverter_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( T2 ),
       .io_mem_resp_bits_data( T1 ),
       .io_mem_resp_bits_tag( T0 )
  );
  ClientTileLinkIOWrapper_1 ClientTileLinkIOWrapper_2(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_in_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_in_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_in_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_out_acquire_ready( RocketChipTileLinkArbiter_io_clients_0_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_out_grant_valid( RocketChipTileLinkArbiter_io_clients_0_grant_valid ),
       .io_out_grant_bits_addr_beat( RocketChipTileLinkArbiter_io_clients_0_grant_bits_addr_beat ),
       .io_out_grant_bits_data( RocketChipTileLinkArbiter_io_clients_0_grant_bits_data ),
       .io_out_grant_bits_client_xact_id( RocketChipTileLinkArbiter_io_clients_0_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( RocketChipTileLinkArbiter_io_clients_0_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( RocketChipTileLinkArbiter_io_clients_0_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( RocketChipTileLinkArbiter_io_clients_0_grant_bits_g_type ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_out_probe_valid( RocketChipTileLinkArbiter_io_clients_0_probe_valid ),
       .io_out_probe_bits_addr_block( RocketChipTileLinkArbiter_io_clients_0_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( RocketChipTileLinkArbiter_io_clients_0_probe_bits_p_type ),
       .io_out_release_ready( RocketChipTileLinkArbiter_io_clients_0_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_data(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_voluntary(  )
  );
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_0_req_cmd_ready,
    output io_mem_0_req_cmd_valid,
    output[25:0] io_mem_0_req_cmd_bits_addr,
    output[5:0] io_mem_0_req_cmd_bits_tag,
    output io_mem_0_req_cmd_bits_rw,
    input  io_mem_0_req_data_ready,
    output io_mem_0_req_data_valid,
    output[127:0] io_mem_0_req_data_bits_data,
    output io_mem_0_resp_ready,
    input  io_mem_0_resp_valid,
    input [127:0] io_mem_0_resp_bits_data,
    input [5:0] io_mem_0_resp_bits_tag,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input  io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    output io_tiles_cached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input  io_tiles_cached_0_release_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [127:0] io_tiles_cached_0_release_bits_data,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input  io_tiles_cached_0_release_bits_voluntary,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input  io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_tiles_uncached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[11:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr
    //input  io_mem_backup_ctrl_en
    //input  io_mem_backup_ctrl_in_valid
    //input  io_mem_backup_ctrl_out_ready
    //output io_mem_backup_ctrl_out_valid
);

  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_pcr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire[11:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_addr_block;
  wire htif_io_mem_acquire_bits_client_xact_id;
  wire[1:0] htif_io_mem_acquire_bits_addr_beat;
  wire[127:0] htif_io_mem_acquire_bits_data;
  wire htif_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] htif_io_mem_acquire_bits_a_type;
  wire[16:0] htif_io_mem_acquire_bits_union;
  wire htif_io_mem_grant_ready;
  wire outmemsys_io_tiles_cached_0_acquire_ready;
  wire outmemsys_io_tiles_cached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire[127:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire outmemsys_io_tiles_cached_0_probe_valid;
  wire[25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire outmemsys_io_tiles_cached_0_release_ready;
  wire outmemsys_io_tiles_uncached_0_acquire_ready;
  wire outmemsys_io_tiles_uncached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[127:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire outmemsys_io_htif_uncached_acquire_ready;
  wire outmemsys_io_htif_uncached_grant_valid;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_addr_beat;
  wire[127:0] outmemsys_io_htif_uncached_grant_bits_data;
  wire outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  wire outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_g_type;
  wire outmemsys_io_mem_0_req_cmd_valid;
  wire[25:0] outmemsys_io_mem_0_req_cmd_bits_addr;
  wire[5:0] outmemsys_io_mem_0_req_cmd_bits_tag;
  wire outmemsys_io_mem_0_req_cmd_bits_rw;
  wire outmemsys_io_mem_0_req_data_valid;
  wire[127:0] outmemsys_io_mem_0_req_data_bits_data;
  wire outmemsys_io_mem_0_resp_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
  assign io_htif_0_ipi_rep_bits = {1{$random}};
//  assign io_htif_0_id = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_mem_0_resp_ready = outmemsys_io_mem_0_resp_ready;
  assign io_mem_0_req_data_bits_data = outmemsys_io_mem_0_req_data_bits_data;
  assign io_mem_0_req_data_valid = outmemsys_io_mem_0_req_data_valid;
  assign io_mem_0_req_cmd_bits_rw = outmemsys_io_mem_0_req_cmd_bits_rw;
  assign io_mem_0_req_cmd_bits_tag = outmemsys_io_mem_0_req_cmd_bits_tag;
  assign io_mem_0_req_cmd_bits_addr = outmemsys_io_mem_0_req_cmd_bits_addr;
  assign io_mem_0_req_cmd_valid = outmemsys_io_mem_0_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_mem_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_mem_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
// synthesis translate_on
`endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_cached_0_acquire_ready( outmemsys_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( outmemsys_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( outmemsys_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_data( outmemsys_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_grant_bits_client_xact_id( outmemsys_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( outmemsys_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( outmemsys_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( outmemsys_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( outmemsys_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( outmemsys_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_tiles_cached_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_tiles_uncached_0_acquire_ready( outmemsys_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( outmemsys_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( outmemsys_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_data( outmemsys_io_tiles_uncached_0_grant_bits_data ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( outmemsys_io_tiles_uncached_0_grant_bits_g_type ),
       .io_htif_uncached_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_htif_uncached_acquire_valid( htif_io_mem_acquire_valid ),
       .io_htif_uncached_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_htif_uncached_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_htif_uncached_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_htif_uncached_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_htif_uncached_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_htif_uncached_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_htif_uncached_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_htif_uncached_grant_ready( htif_io_mem_grant_ready ),
       .io_htif_uncached_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_htif_uncached_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_htif_uncached_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_htif_uncached_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_htif_uncached_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_htif_uncached_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_htif_uncached_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_incoherent_0( htif_io_cpu_0_reset ),
       .io_mem_0_req_cmd_ready( io_mem_0_req_cmd_ready ),
       .io_mem_0_req_cmd_valid( outmemsys_io_mem_0_req_cmd_valid ),
       .io_mem_0_req_cmd_bits_addr( outmemsys_io_mem_0_req_cmd_bits_addr ),
       .io_mem_0_req_cmd_bits_tag( outmemsys_io_mem_0_req_cmd_bits_tag ),
       .io_mem_0_req_cmd_bits_rw( outmemsys_io_mem_0_req_cmd_bits_rw ),
       .io_mem_0_req_data_ready( io_mem_0_req_data_ready ),
       .io_mem_0_req_data_valid( outmemsys_io_mem_0_req_data_valid ),
       .io_mem_0_req_data_bits_data( outmemsys_io_mem_0_req_data_bits_data ),
       .io_mem_0_resp_ready( outmemsys_io_mem_0_resp_ready ),
       .io_mem_0_resp_valid( io_mem_0_resp_valid ),
       .io_mem_0_resp_bits_data( io_mem_0_resp_bits_data ),
       .io_mem_0_resp_bits_tag( io_mem_0_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
endmodule

module BTB(input clk, input reset,
    input  io_req_valid,
    input [38:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output io_resp_bits_mask,
    output io_resp_bits_bridx,
    output[38:0] io_resp_bits_target,
    output[2:0] io_resp_bits_entry,
    output[3:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_btb_update_valid,
    input  io_btb_update_bits_prediction_valid,
    input  io_btb_update_bits_prediction_bits_taken,
    input  io_btb_update_bits_prediction_bits_mask,
    input  io_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_btb_update_bits_prediction_bits_target,
    input [2:0] io_btb_update_bits_prediction_bits_entry,
    input [3:0] io_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_btb_update_bits_pc,
    input [38:0] io_btb_update_bits_target,
    input  io_btb_update_bits_taken,
    input  io_btb_update_bits_isJump,
    input  io_btb_update_bits_isReturn,
    input [38:0] io_btb_update_bits_br_pc,
    input  io_bht_update_valid,
    input  io_bht_update_bits_prediction_valid,
    input  io_bht_update_bits_prediction_bits_taken,
    input  io_bht_update_bits_prediction_bits_mask,
    input  io_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_bht_update_bits_prediction_bits_target,
    input [2:0] io_bht_update_bits_prediction_bits_entry,
    input [3:0] io_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_bht_update_bits_pc,
    input  io_bht_update_bits_taken,
    input  io_bht_update_bits_mispredict,
    input  io_ras_update_valid,
    input  io_ras_update_bits_isCall,
    input  io_ras_update_bits_isReturn,
    input [38:0] io_ras_update_bits_returnAddr,
    input  io_ras_update_bits_prediction_valid,
    input  io_ras_update_bits_prediction_bits_taken,
    input  io_ras_update_bits_prediction_bits_mask,
    input  io_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_ras_update_bits_prediction_bits_target,
    input [2:0] io_ras_update_bits_prediction_bits_entry,
    input [3:0] io_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_ras_update_bits_prediction_bits_bht_value,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [38:0] R4;
  wire[38:0] T5;
  wire T6;
  reg  R7;
  wire T465;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10 [15:0];
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  reg [3:0] R25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[2:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg  isJump_7;
  wire T35;
  reg  R36;
  wire T37;
  wire T38;
  wire T39;
  wire[7:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  reg [2:0] R43;
  wire[2:0] T466;
  wire[2:0] T44;
  wire[2:0] T45;
  wire T46;
  wire T47;
  reg [2:0] R48;
  wire[2:0] T49;
  reg  updateHit;
  wire T50;
  wire T51;
  wire[7:0] hits;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[3:0] T54;
  wire[1:0] T55;
  wire T56;
  wire[3:0] T57;
  wire[3:0] pageHit;
  reg [3:0] pageValid;
  wire[3:0] T467;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T60;
  wire[3:0] pageReplEn;
  wire[3:0] tgtPageReplEn;
  wire[3:0] tgtPageRepl;
  wire[3:0] T61;
  wire[3:0] T468;
  wire T62;
  wire[3:0] T63;
  wire[2:0] T64;
  wire[3:0] idxPageUpdateOH;
  wire[3:0] idxPageRepl;
  wire[3:0] T65;
  reg [1:0] R66;
  wire[1:0] T469;
  wire[1:0] T67;
  wire[1:0] T68;
  wire T69;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire[3:0] updatePageHit;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[1:0] T72;
  wire T73;
  wire[26:0] T74;
  reg [38:0] R75;
  wire[38:0] T76;
  wire[26:0] T77;
  reg [26:0] pages [3:0];
  wire[26:0] T78;
  wire[26:0] T79;
  wire[26:0] T80;
  wire[26:0] T81;
  wire T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[26:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire[26:0] T92;
  wire[26:0] T93;
  wire[26:0] T94;
  wire[26:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[26:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire[26:0] T105;
  wire[1:0] T106;
  wire T107;
  wire[26:0] T108;
  wire T109;
  wire[26:0] T110;
  wire useUpdatePageHit;
  wire samePage;
  wire[26:0] T111;
  wire[26:0] T112;
  wire doTgtPageRepl;
  wire T113;
  wire usePageHit;
  wire[3:0] T114;
  wire[3:0] T115;
  wire T116;
  wire[3:0] idxPageReplEn;
  wire T117;
  wire[3:0] T118;
  wire[3:0] T119;
  wire[1:0] T120;
  wire T121;
  wire[26:0] T122;
  wire[26:0] T123;
  wire T124;
  wire[26:0] T125;
  wire[1:0] T126;
  wire T127;
  wire[26:0] T128;
  wire T129;
  wire[26:0] T130;
  wire[3:0] idxPagesOH_0;
  wire[3:0] T131;
  wire[1:0] T132;
  reg [1:0] idxPages [7:0];
  wire[1:0] T133;
  wire[1:0] T470;
  wire T471;
  wire[1:0] T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire T475;
  wire T134;
  wire[3:0] T135;
  wire[3:0] idxPagesOH_1;
  wire[3:0] T136;
  wire[1:0] T137;
  wire[1:0] T138;
  wire T139;
  wire[3:0] T140;
  wire[3:0] idxPagesOH_2;
  wire[3:0] T141;
  wire[1:0] T142;
  wire T143;
  wire[3:0] T144;
  wire[3:0] idxPagesOH_3;
  wire[3:0] T145;
  wire[1:0] T146;
  wire[3:0] T147;
  wire[1:0] T148;
  wire T149;
  wire[3:0] T150;
  wire[3:0] idxPagesOH_4;
  wire[3:0] T151;
  wire[1:0] T152;
  wire T153;
  wire[3:0] T154;
  wire[3:0] idxPagesOH_5;
  wire[3:0] T155;
  wire[1:0] T156;
  wire[1:0] T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] idxPagesOH_6;
  wire[3:0] T160;
  wire[1:0] T161;
  wire T162;
  wire[3:0] T163;
  wire[3:0] idxPagesOH_7;
  wire[3:0] T164;
  wire[1:0] T165;
  wire[7:0] T166;
  wire[7:0] T167;
  wire[7:0] T168;
  wire[3:0] T169;
  wire[1:0] T170;
  wire T171;
  wire[11:0] T172;
  wire[11:0] T173;
  reg [11:0] idxs [7:0];
  wire[11:0] T174;
  wire[11:0] T476;
  wire T175;
  wire[11:0] T176;
  wire[1:0] T177;
  wire T178;
  wire[11:0] T179;
  wire T180;
  wire[11:0] T181;
  wire[3:0] T182;
  wire[1:0] T183;
  wire T184;
  wire[11:0] T185;
  wire T186;
  wire[11:0] T187;
  wire[1:0] T188;
  wire T189;
  wire[11:0] T190;
  wire T191;
  wire[11:0] T192;
  reg [7:0] idxValid;
  wire[7:0] T477;
  wire[7:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[7:0] T196;
  wire[7:0] T197;
  wire[7:0] T198;
  wire[7:0] T199;
  wire[7:0] T200;
  wire[3:0] T201;
  wire[1:0] T202;
  wire T203;
  wire[3:0] T204;
  wire[3:0] T205;
  wire[3:0] tgtPagesOH_0;
  wire[3:0] T206;
  wire[1:0] T207;
  reg [1:0] tgtPages [7:0];
  wire[1:0] T208;
  wire[1:0] T478;
  wire T479;
  wire[1:0] T480;
  wire[1:0] T481;
  wire[3:0] T209;
  wire[1:0] T482;
  wire T483;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] tgtPagesOH_1;
  wire[3:0] T213;
  wire[1:0] T214;
  wire[1:0] T215;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] tgtPagesOH_2;
  wire[3:0] T219;
  wire[1:0] T220;
  wire T221;
  wire[3:0] T222;
  wire[3:0] T223;
  wire[3:0] tgtPagesOH_3;
  wire[3:0] T224;
  wire[1:0] T225;
  wire[3:0] T226;
  wire[1:0] T227;
  wire T228;
  wire[3:0] T229;
  wire[3:0] T230;
  wire[3:0] tgtPagesOH_4;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[3:0] tgtPagesOH_5;
  wire[3:0] T236;
  wire[1:0] T237;
  wire[1:0] T238;
  wire T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] tgtPagesOH_6;
  wire[3:0] T242;
  wire[1:0] T243;
  wire T244;
  wire[3:0] T245;
  wire[3:0] T246;
  wire[3:0] tgtPagesOH_7;
  wire[3:0] T247;
  wire[1:0] T248;
  wire T249;
  wire T250;
  reg  isJump_6;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  reg  isJump_5;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  reg  isJump_4;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  reg  isJump_3;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  reg  isJump_2;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  reg  isJump_1;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  reg  isJump_0;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[2:0] T292;
  wire T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[2:0] T484;
  wire[1:0] T485;
  wire T486;
  wire[1:0] T487;
  wire[1:0] T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[1:0] T492;
  wire T493;
  wire T494;
  wire[38:0] T297;
  wire[38:0] T298;
  wire[38:0] T299;
  wire[11:0] T300;
  wire[11:0] T301;
  wire[11:0] T302;
  reg [11:0] tgts [7:0];
  wire[11:0] T303;
  wire[11:0] T495;
  wire T304;
  wire[11:0] T305;
  wire[11:0] T306;
  wire[11:0] T307;
  wire T308;
  wire[11:0] T309;
  wire[11:0] T310;
  wire[11:0] T311;
  wire T312;
  wire[11:0] T313;
  wire[11:0] T314;
  wire[11:0] T315;
  wire T316;
  wire[11:0] T317;
  wire[11:0] T318;
  wire[11:0] T319;
  wire T320;
  wire[11:0] T321;
  wire[11:0] T322;
  wire[11:0] T323;
  wire T324;
  wire[11:0] T325;
  wire[11:0] T326;
  wire[11:0] T327;
  wire T328;
  wire[11:0] T329;
  wire[11:0] T330;
  wire T331;
  wire[26:0] T332;
  wire[26:0] T333;
  wire[26:0] T334;
  wire T335;
  wire[3:0] T336;
  wire[3:0] T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire T341;
  wire[3:0] T342;
  wire[3:0] T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire T350;
  wire[3:0] T351;
  wire[3:0] T352;
  wire T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire T356;
  wire[3:0] T357;
  wire T358;
  wire[26:0] T359;
  wire[26:0] T360;
  wire[26:0] T361;
  wire T362;
  wire[26:0] T363;
  wire[26:0] T364;
  wire[26:0] T365;
  wire T366;
  wire[26:0] T367;
  wire[26:0] T368;
  wire T369;
  wire[38:0] T370;
  reg [38:0] R371;
  wire[38:0] T372;
  wire T373;
  wire T374;
  wire[1:0] T375;
  wire T376;
  wire T377;
  reg  R378;
  wire T496;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  reg [1:0] R385;
  wire[1:0] T497;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  reg [38:0] R398;
  wire[38:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  reg  useRAS_7;
  wire T406;
  reg  R407;
  wire T408;
  wire T409;
  wire T410;
  wire[7:0] T411;
  wire[2:0] T412;
  wire T413;
  wire T414;
  wire T415;
  reg  useRAS_6;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  reg  useRAS_5;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  reg  useRAS_4;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  reg  useRAS_3;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  reg  useRAS_2;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  reg  useRAS_1;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  reg  useRAS_0;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  reg [0:0] brIdx [7:0];
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R7 = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      T10[initvar] = {1{$random}};
    R25 = {1{$random}};
    isJump_7 = {1{$random}};
    R36 = {1{$random}};
    R43 = {1{$random}};
    R48 = {1{$random}};
    updateHit = {1{$random}};
    pageValid = {1{$random}};
    R66 = {1{$random}};
    R75 = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    isJump_6 = {1{$random}};
    isJump_5 = {1{$random}};
    isJump_4 = {1{$random}};
    isJump_3 = {1{$random}};
    isJump_2 = {1{$random}};
    isJump_1 = {1{$random}};
    isJump_0 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R371 = {2{$random}};
    R378 = {1{$random}};
    R385 = {1{$random}};
    R398 = {2{$random}};
    useRAS_7 = {1{$random}};
    R407 = {1{$random}};
    useRAS_6 = {1{$random}};
    useRAS_5 = {1{$random}};
    useRAS_4 = {1{$random}};
    useRAS_3 = {1{$random}};
    useRAS_2 = {1{$random}};
    useRAS_1 = {1{$random}};
    useRAS_0 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      brIdx[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_btb_update_valid ? io_btb_update_bits_target : R4;
  assign T6 = R7 ^ 1'h1;
  assign T465 = reset ? 1'h0 : io_btb_update_valid;
  assign io_resp_bits_bht_value = T8;
  assign T8 = T9;
  assign T9 = T10[T24];
  assign T12 = {io_bht_update_bits_taken, T13};
  assign T13 = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = T17 | T16;
  assign T16 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T17 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T18 = T20 & T19;
  assign T19 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T20 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22 = T23 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T23 = io_bht_update_bits_pc[3'h5:2'h2];
  assign T24 = T294 ^ R25;
  assign T26 = T293 ? T291 : T27;
  assign T27 = T31 ? T28 : R25;
  assign T28 = {T30, T29};
  assign T29 = R25[2'h3:1'h1];
  assign T30 = T8[1'h0:1'h0];
  assign T31 = T290 & T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T249 | T34;
  assign T34 = T51 ? isJump_7 : 1'h0;
  assign T35 = T38 ? R36 : isJump_7;
  assign T37 = io_btb_update_valid ? io_btb_update_bits_isJump : R36;
  assign T38 = R7 & T39;
  assign T39 = T40[3'h7:3'h7];
  assign T40 = 1'h1 << T41;
  assign T41 = T42;
  assign T42 = updateHit ? R48 : R43;
  assign T466 = reset ? 3'h0 : T44;
  assign T44 = T46 ? T45 : R43;
  assign T45 = R43 + 3'h1;
  assign T46 = R7 & T47;
  assign T47 = updateHit ^ 1'h1;
  assign T49 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : R48;
  assign T50 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : updateHit;
  assign T51 = hits[3'h7:3'h7];
  assign hits = T166 & T52;
  assign T52 = T53;
  assign T53 = {T147, T54};
  assign T54 = {T138, T55};
  assign T55 = {T134, T56};
  assign T56 = T57 != 4'h0;
  assign T57 = idxPagesOH_0 & pageHit;
  assign pageHit = T118 & pageValid;
  assign T467 = reset ? 4'h0 : T58;
  assign T58 = io_invalidate ? 4'h0 : T59;
  assign T59 = T117 ? T60 : pageValid;
  assign T60 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 4'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T61;
  assign T61 = T63 | T468;
  assign T468 = {3'h0, T62};
  assign T62 = idxPageUpdateOH[2'h3:2'h3];
  assign T63 = T64 << 1'h1;
  assign T64 = idxPageUpdateOH[2'h2:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T65;
  assign T65 = 1'h1 << R66;
  assign T469 = reset ? 2'h0 : T67;
  assign T67 = T69 ? T68 : R66;
  assign T68 = R66 + 2'h1;
  assign T69 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = useUpdatePageHit ^ 1'h1;
  assign updatePageHit = T70 & pageValid;
  assign T70 = T71;
  assign T71 = {T106, T72};
  assign T72 = {T104, T73};
  assign T73 = T77 == T74;
  assign T74 = R75 >> 4'hc;
  assign T76 = io_btb_update_valid ? io_btb_update_bits_pc : R75;
  assign T77 = pages[2'h0];
  assign T79 = T82 ? T81 : T80;
  assign T80 = R75 >> 4'hc;
  assign T81 = io_req_bits_addr >> 4'hc;
  assign T82 = T83 != 4'h0;
  assign T83 = idxPageUpdateOH & 4'h5;
  assign T84 = R7 & T85;
  assign T85 = T87 & T86;
  assign T86 = pageReplEn[2'h3:2'h3];
  assign T87 = T82 ? doTgtPageRepl : doIdxPageRepl;
  assign T89 = R7 & T90;
  assign T90 = T87 & T91;
  assign T91 = pageReplEn[1'h1:1'h1];
  assign T93 = T82 ? T95 : T94;
  assign T94 = io_req_bits_addr >> 4'hc;
  assign T95 = R75 >> 4'hc;
  assign T96 = R7 & T97;
  assign T97 = T99 & T98;
  assign T98 = pageReplEn[2'h2:2'h2];
  assign T99 = T82 ? doIdxPageRepl : doTgtPageRepl;
  assign T101 = R7 & T102;
  assign T102 = T99 & T103;
  assign T103 = pageReplEn[1'h0:1'h0];
  assign T104 = T105 == T74;
  assign T105 = pages[2'h1];
  assign T106 = {T109, T107};
  assign T107 = T108 == T74;
  assign T108 = pages[2'h2];
  assign T109 = T110 == T74;
  assign T110 = pages[2'h3];
  assign useUpdatePageHit = updatePageHit != 4'h0;
  assign samePage = T112 == T111;
  assign T111 = io_req_bits_addr >> 4'hc;
  assign T112 = R75 >> 4'hc;
  assign doTgtPageRepl = T116 & T113;
  assign T113 = usePageHit ^ 1'h1;
  assign usePageHit = T114 != 4'h0;
  assign T114 = pageHit & T115;
  assign T115 = ~ idxPageReplEn;
  assign T116 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 4'h0;
  assign T117 = R7 & doPageRepl;
  assign T118 = T119;
  assign T119 = {T126, T120};
  assign T120 = {T124, T121};
  assign T121 = T123 == T122;
  assign T122 = io_req_bits_addr >> 4'hc;
  assign T123 = pages[2'h0];
  assign T124 = T125 == T122;
  assign T125 = pages[2'h1];
  assign T126 = {T129, T127};
  assign T127 = T128 == T122;
  assign T128 = pages[2'h2];
  assign T129 = T130 == T122;
  assign T130 = pages[2'h3];
  assign idxPagesOH_0 = T131[2'h3:1'h0];
  assign T131 = 1'h1 << T132;
  assign T132 = idxPages[3'h0];
  assign T470 = {T475, T471};
  assign T471 = T472[1'h1:1'h1];
  assign T472 = T474 | T473;
  assign T473 = idxPageUpdateOH[1'h1:1'h0];
  assign T474 = idxPageUpdateOH[2'h3:2'h2];
  assign T475 = T474 != 2'h0;
  assign T134 = T135 != 4'h0;
  assign T135 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T136[2'h3:1'h0];
  assign T136 = 1'h1 << T137;
  assign T137 = idxPages[3'h1];
  assign T138 = {T143, T139};
  assign T139 = T140 != 4'h0;
  assign T140 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T141[2'h3:1'h0];
  assign T141 = 1'h1 << T142;
  assign T142 = idxPages[3'h2];
  assign T143 = T144 != 4'h0;
  assign T144 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T145[2'h3:1'h0];
  assign T145 = 1'h1 << T146;
  assign T146 = idxPages[3'h3];
  assign T147 = {T157, T148};
  assign T148 = {T153, T149};
  assign T149 = T150 != 4'h0;
  assign T150 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T151[2'h3:1'h0];
  assign T151 = 1'h1 << T152;
  assign T152 = idxPages[3'h4];
  assign T153 = T154 != 4'h0;
  assign T154 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T155[2'h3:1'h0];
  assign T155 = 1'h1 << T156;
  assign T156 = idxPages[3'h5];
  assign T157 = {T162, T158};
  assign T158 = T159 != 4'h0;
  assign T159 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T160[2'h3:1'h0];
  assign T160 = 1'h1 << T161;
  assign T161 = idxPages[3'h6];
  assign T162 = T163 != 4'h0;
  assign T163 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T164[2'h3:1'h0];
  assign T164 = 1'h1 << T165;
  assign T165 = idxPages[3'h7];
  assign T166 = idxValid & T167;
  assign T167 = T168;
  assign T168 = {T182, T169};
  assign T169 = {T177, T170};
  assign T170 = {T175, T171};
  assign T171 = T173 == T172;
  assign T172 = io_req_bits_addr[4'hb:1'h0];
  assign T173 = idxs[3'h0];
  assign T476 = R75[4'hb:1'h0];
  assign T175 = T176 == T172;
  assign T176 = idxs[3'h1];
  assign T177 = {T180, T178};
  assign T178 = T179 == T172;
  assign T179 = idxs[3'h2];
  assign T180 = T181 == T172;
  assign T181 = idxs[3'h3];
  assign T182 = {T188, T183};
  assign T183 = {T186, T184};
  assign T184 = T185 == T172;
  assign T185 = idxs[3'h4];
  assign T186 = T187 == T172;
  assign T187 = idxs[3'h5];
  assign T188 = {T191, T189};
  assign T189 = T190 == T172;
  assign T190 = idxs[3'h6];
  assign T191 = T192 == T172;
  assign T192 = idxs[3'h7];
  assign T477 = reset ? 8'h0 : T193;
  assign T193 = io_invalidate ? 8'h0 : T194;
  assign T194 = R7 ? T195 : idxValid;
  assign T195 = T197 | T196;
  assign T196 = 1'h1 << T42;
  assign T197 = idxValid & T198;
  assign T198 = ~ T199;
  assign T199 = T200;
  assign T200 = {T226, T201};
  assign T201 = {T215, T202};
  assign T202 = {T210, T203};
  assign T203 = T204 != 4'h0;
  assign T204 = pageReplEn & T205;
  assign T205 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T206[2'h3:1'h0];
  assign T206 = 1'h1 << T207;
  assign T207 = tgtPages[3'h0];
  assign T478 = {T483, T479};
  assign T479 = T480[1'h1:1'h1];
  assign T480 = T482 | T481;
  assign T481 = T209[1'h1:1'h0];
  assign T209 = usePageHit ? pageHit : tgtPageRepl;
  assign T482 = T209[2'h3:2'h2];
  assign T483 = T482 != 2'h0;
  assign T210 = T211 != 4'h0;
  assign T211 = pageReplEn & T212;
  assign T212 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T213[2'h3:1'h0];
  assign T213 = 1'h1 << T214;
  assign T214 = tgtPages[3'h1];
  assign T215 = {T221, T216};
  assign T216 = T217 != 4'h0;
  assign T217 = pageReplEn & T218;
  assign T218 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T219[2'h3:1'h0];
  assign T219 = 1'h1 << T220;
  assign T220 = tgtPages[3'h2];
  assign T221 = T222 != 4'h0;
  assign T222 = pageReplEn & T223;
  assign T223 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T224[2'h3:1'h0];
  assign T224 = 1'h1 << T225;
  assign T225 = tgtPages[3'h3];
  assign T226 = {T238, T227};
  assign T227 = {T233, T228};
  assign T228 = T229 != 4'h0;
  assign T229 = pageReplEn & T230;
  assign T230 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T231[2'h3:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = tgtPages[3'h4];
  assign T233 = T234 != 4'h0;
  assign T234 = pageReplEn & T235;
  assign T235 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T236[2'h3:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = tgtPages[3'h5];
  assign T238 = {T244, T239};
  assign T239 = T240 != 4'h0;
  assign T240 = pageReplEn & T241;
  assign T241 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T242[2'h3:1'h0];
  assign T242 = 1'h1 << T243;
  assign T243 = tgtPages[3'h6];
  assign T244 = T245 != 4'h0;
  assign T245 = pageReplEn & T246;
  assign T246 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T247[2'h3:1'h0];
  assign T247 = 1'h1 << T248;
  assign T248 = tgtPages[3'h7];
  assign T249 = T255 | T250;
  assign T250 = T254 ? isJump_6 : 1'h0;
  assign T251 = T252 ? R36 : isJump_6;
  assign T252 = R7 & T253;
  assign T253 = T40[3'h6:3'h6];
  assign T254 = hits[3'h6:3'h6];
  assign T255 = T261 | T256;
  assign T256 = T260 ? isJump_5 : 1'h0;
  assign T257 = T258 ? R36 : isJump_5;
  assign T258 = R7 & T259;
  assign T259 = T40[3'h5:3'h5];
  assign T260 = hits[3'h5:3'h5];
  assign T261 = T267 | T262;
  assign T262 = T266 ? isJump_4 : 1'h0;
  assign T263 = T264 ? R36 : isJump_4;
  assign T264 = R7 & T265;
  assign T265 = T40[3'h4:3'h4];
  assign T266 = hits[3'h4:3'h4];
  assign T267 = T273 | T268;
  assign T268 = T272 ? isJump_3 : 1'h0;
  assign T269 = T270 ? R36 : isJump_3;
  assign T270 = R7 & T271;
  assign T271 = T40[2'h3:2'h3];
  assign T272 = hits[2'h3:2'h3];
  assign T273 = T279 | T274;
  assign T274 = T278 ? isJump_2 : 1'h0;
  assign T275 = T276 ? R36 : isJump_2;
  assign T276 = R7 & T277;
  assign T277 = T40[2'h2:2'h2];
  assign T278 = hits[2'h2:2'h2];
  assign T279 = T285 | T280;
  assign T280 = T284 ? isJump_1 : 1'h0;
  assign T281 = T282 ? R36 : isJump_1;
  assign T282 = R7 & T283;
  assign T283 = T40[1'h1:1'h1];
  assign T284 = hits[1'h1:1'h1];
  assign T285 = T289 ? isJump_0 : 1'h0;
  assign T286 = T287 ? R36 : isJump_0;
  assign T287 = R7 & T288;
  assign T288 = T40[1'h0:1'h0];
  assign T289 = hits[1'h0:1'h0];
  assign T290 = io_req_valid & io_resp_valid;
  assign T291 = {io_bht_update_bits_taken, T292};
  assign T292 = io_bht_update_bits_prediction_bits_bht_history[2'h3:1'h1];
  assign T293 = T21 & io_bht_update_bits_mispredict;
  assign T294 = io_req_bits_addr[3'h5:2'h2];
  assign io_resp_bits_bht_history = T295;
  assign T295 = R25;
  assign io_resp_bits_entry = T484;
  assign T484 = {T494, T485};
  assign T485 = {T493, T486};
  assign T486 = T487[1'h1:1'h1];
  assign T487 = T492 | T488;
  assign T488 = T489[1'h1:1'h0];
  assign T489 = T491 | T490;
  assign T490 = hits[2'h3:1'h0];
  assign T491 = hits[3'h7:3'h4];
  assign T492 = T489[2'h3:2'h2];
  assign T493 = T492 != 2'h0;
  assign T494 = T491 != 4'h0;
  assign io_resp_bits_target = T297;
  assign T297 = T457 ? io_ras_update_bits_returnAddr : T298;
  assign T298 = T403 ? T370 : T299;
  assign T299 = {T332, T300};
  assign T300 = T305 | T301;
  assign T301 = T304 ? T302 : 12'h0;
  assign T302 = tgts[3'h7];
  assign T495 = io_req_bits_addr[4'hb:1'h0];
  assign T304 = hits[3'h7:3'h7];
  assign T305 = T309 | T306;
  assign T306 = T308 ? T307 : 12'h0;
  assign T307 = tgts[3'h6];
  assign T308 = hits[3'h6:3'h6];
  assign T309 = T313 | T310;
  assign T310 = T312 ? T311 : 12'h0;
  assign T311 = tgts[3'h5];
  assign T312 = hits[3'h5:3'h5];
  assign T313 = T317 | T314;
  assign T314 = T316 ? T315 : 12'h0;
  assign T315 = tgts[3'h4];
  assign T316 = hits[3'h4:3'h4];
  assign T317 = T321 | T318;
  assign T318 = T320 ? T319 : 12'h0;
  assign T319 = tgts[3'h3];
  assign T320 = hits[2'h3:2'h3];
  assign T321 = T325 | T322;
  assign T322 = T324 ? T323 : 12'h0;
  assign T323 = tgts[3'h2];
  assign T324 = hits[2'h2:2'h2];
  assign T325 = T329 | T326;
  assign T326 = T328 ? T327 : 12'h0;
  assign T327 = tgts[3'h1];
  assign T328 = hits[1'h1:1'h1];
  assign T329 = T331 ? T330 : 12'h0;
  assign T330 = tgts[3'h0];
  assign T331 = hits[1'h0:1'h0];
  assign T332 = T359 | T333;
  assign T333 = T335 ? T334 : 27'h0;
  assign T334 = pages[2'h3];
  assign T335 = T336[2'h3:2'h3];
  assign T336 = T339 | T337;
  assign T337 = T338 ? tgtPagesOH_7 : 4'h0;
  assign T338 = hits[3'h7:3'h7];
  assign T339 = T342 | T340;
  assign T340 = T341 ? tgtPagesOH_6 : 4'h0;
  assign T341 = hits[3'h6:3'h6];
  assign T342 = T345 | T343;
  assign T343 = T344 ? tgtPagesOH_5 : 4'h0;
  assign T344 = hits[3'h5:3'h5];
  assign T345 = T348 | T346;
  assign T346 = T347 ? tgtPagesOH_4 : 4'h0;
  assign T347 = hits[3'h4:3'h4];
  assign T348 = T351 | T349;
  assign T349 = T350 ? tgtPagesOH_3 : 4'h0;
  assign T350 = hits[2'h3:2'h3];
  assign T351 = T354 | T352;
  assign T352 = T353 ? tgtPagesOH_2 : 4'h0;
  assign T353 = hits[2'h2:2'h2];
  assign T354 = T357 | T355;
  assign T355 = T356 ? tgtPagesOH_1 : 4'h0;
  assign T356 = hits[1'h1:1'h1];
  assign T357 = T358 ? tgtPagesOH_0 : 4'h0;
  assign T358 = hits[1'h0:1'h0];
  assign T359 = T363 | T360;
  assign T360 = T362 ? T361 : 27'h0;
  assign T361 = pages[2'h2];
  assign T362 = T336[2'h2:2'h2];
  assign T363 = T367 | T364;
  assign T364 = T366 ? T365 : 27'h0;
  assign T365 = pages[2'h1];
  assign T366 = T336[1'h1:1'h1];
  assign T367 = T369 ? T368 : 27'h0;
  assign T368 = pages[2'h0];
  assign T369 = T336[1'h0:1'h0];
  assign T370 = T402 ? R398 : R371;
  assign T372 = T373 ? io_ras_update_bits_returnAddr : R371;
  assign T373 = T397 & T374;
  assign T374 = T375[1'h0:1'h0];
  assign T375 = 1'h1 << T376;
  assign T376 = T377;
  assign T377 = R378 + 1'h1;
  assign T496 = reset ? 1'h0 : T379;
  assign T379 = T382 ? T381 : T380;
  assign T380 = T397 ? T377 : R378;
  assign T381 = R378 - 1'h1;
  assign T382 = T393 & T383;
  assign T383 = T384 ^ 1'h1;
  assign T384 = R385 == 2'h0;
  assign T497 = reset ? 2'h0 : T386;
  assign T386 = io_invalidate ? 2'h0 : T387;
  assign T387 = T382 ? T392 : T388;
  assign T388 = T390 ? T389 : R385;
  assign T389 = R385 + 2'h1;
  assign T390 = T397 & T391;
  assign T391 = R385 < 2'h2;
  assign T392 = R385 - 2'h1;
  assign T393 = io_ras_update_valid & T394;
  assign T394 = T396 & T395;
  assign T395 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T396 = io_ras_update_bits_isCall ^ 1'h1;
  assign T397 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T399 = T400 ? io_ras_update_bits_returnAddr : R398;
  assign T400 = T397 & T401;
  assign T401 = T375[1'h1:1'h1];
  assign T402 = R378;
  assign T403 = T455 & T404;
  assign T404 = T414 | T405;
  assign T405 = T413 ? useRAS_7 : 1'h0;
  assign T406 = T409 ? R407 : useRAS_7;
  assign T408 = io_btb_update_valid ? io_btb_update_bits_isReturn : R407;
  assign T409 = R7 & T410;
  assign T410 = T411[3'h7:3'h7];
  assign T411 = 1'h1 << T412;
  assign T412 = T42;
  assign T413 = hits[3'h7:3'h7];
  assign T414 = T420 | T415;
  assign T415 = T419 ? useRAS_6 : 1'h0;
  assign T416 = T417 ? R407 : useRAS_6;
  assign T417 = R7 & T418;
  assign T418 = T411[3'h6:3'h6];
  assign T419 = hits[3'h6:3'h6];
  assign T420 = T426 | T421;
  assign T421 = T425 ? useRAS_5 : 1'h0;
  assign T422 = T423 ? R407 : useRAS_5;
  assign T423 = R7 & T424;
  assign T424 = T411[3'h5:3'h5];
  assign T425 = hits[3'h5:3'h5];
  assign T426 = T432 | T427;
  assign T427 = T431 ? useRAS_4 : 1'h0;
  assign T428 = T429 ? R407 : useRAS_4;
  assign T429 = R7 & T430;
  assign T430 = T411[3'h4:3'h4];
  assign T431 = hits[3'h4:3'h4];
  assign T432 = T438 | T433;
  assign T433 = T437 ? useRAS_3 : 1'h0;
  assign T434 = T435 ? R407 : useRAS_3;
  assign T435 = R7 & T436;
  assign T436 = T411[2'h3:2'h3];
  assign T437 = hits[2'h3:2'h3];
  assign T438 = T444 | T439;
  assign T439 = T443 ? useRAS_2 : 1'h0;
  assign T440 = T441 ? R407 : useRAS_2;
  assign T441 = R7 & T442;
  assign T442 = T411[2'h2:2'h2];
  assign T443 = hits[2'h2:2'h2];
  assign T444 = T450 | T445;
  assign T445 = T449 ? useRAS_1 : 1'h0;
  assign T446 = T447 ? R407 : useRAS_1;
  assign T447 = R7 & T448;
  assign T448 = T411[1'h1:1'h1];
  assign T449 = hits[1'h1:1'h1];
  assign T450 = T454 ? useRAS_0 : 1'h0;
  assign T451 = T452 ? R407 : useRAS_0;
  assign T452 = R7 & T453;
  assign T453 = T411[1'h0:1'h0];
  assign T454 = hits[1'h0:1'h0];
  assign T455 = T456 ^ 1'h1;
  assign T456 = R385 == 2'h0;
  assign T457 = T397 & T404;
  assign io_resp_bits_bridx = T458;
  assign T458 = brIdx[io_resp_bits_entry];
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_taken = T460;
  assign T460 = T461 ? 1'h0 : io_resp_valid;
  assign T461 = T462 & T32;
  assign T462 = T463 ^ 1'h1;
  assign T463 = T8[1'h0:1'h0];
  assign io_resp_valid = T464;
  assign T464 = hits != 8'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
// synthesis translate_on
`endif
    if(io_btb_update_valid) begin
      R4 <= io_btb_update_bits_target;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_btb_update_valid;
    end
    if (T21)
      T10[T22] <= T12;
    if(T293) begin
      R25 <= T291;
    end else if(T31) begin
      R25 <= T28;
    end
    if(T38) begin
      isJump_7 <= R36;
    end
    if(io_btb_update_valid) begin
      R36 <= io_btb_update_bits_isJump;
    end
    if(reset) begin
      R43 <= 3'h0;
    end else if(T46) begin
      R43 <= T45;
    end
    if(io_btb_update_valid) begin
      R48 <= io_btb_update_bits_prediction_bits_entry;
    end
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end
    if(reset) begin
      pageValid <= 4'h0;
    end else if(io_invalidate) begin
      pageValid <= 4'h0;
    end else if(T117) begin
      pageValid <= T60;
    end
    if(reset) begin
      R66 <= 2'h0;
    end else if(T69) begin
      R66 <= T68;
    end
    if(io_btb_update_valid) begin
      R75 <= io_btb_update_bits_pc;
    end
    if (T84)
      pages[2'h3] <= T79;
    if (T89)
      pages[2'h1] <= T79;
    if (T96)
      pages[2'h2] <= T93;
    if (T101)
      pages[2'h0] <= T93;
    if (R7)
      idxPages[T42] <= T470;
    if (R7)
      idxs[T42] <= T476;
    if(reset) begin
      idxValid <= 8'h0;
    end else if(io_invalidate) begin
      idxValid <= 8'h0;
    end else if(R7) begin
      idxValid <= T195;
    end
    if (R7)
      tgtPages[T42] <= T478;
    if(T252) begin
      isJump_6 <= R36;
    end
    if(T258) begin
      isJump_5 <= R36;
    end
    if(T264) begin
      isJump_4 <= R36;
    end
    if(T270) begin
      isJump_3 <= R36;
    end
    if(T276) begin
      isJump_2 <= R36;
    end
    if(T282) begin
      isJump_1 <= R36;
    end
    if(T287) begin
      isJump_0 <= R36;
    end
    if (R7)
      tgts[T42] <= T495;
    if(T373) begin
      R371 <= io_ras_update_bits_returnAddr;
    end
    if(reset) begin
      R378 <= 1'h0;
    end else if(T382) begin
      R378 <= T381;
    end else if(T397) begin
      R378 <= T377;
    end
    if(reset) begin
      R385 <= 2'h0;
    end else if(io_invalidate) begin
      R385 <= 2'h0;
    end else if(T382) begin
      R385 <= T392;
    end else if(T390) begin
      R385 <= T389;
    end
    if(T400) begin
      R398 <= io_ras_update_bits_returnAddr;
    end
    if(T409) begin
      useRAS_7 <= R407;
    end
    if(io_btb_update_valid) begin
      R407 <= io_btb_update_bits_isReturn;
    end
    if(T417) begin
      useRAS_6 <= R407;
    end
    if(T423) begin
      useRAS_5 <= R407;
    end
    if(T429) begin
      useRAS_4 <= R407;
    end
    if(T435) begin
      useRAS_3 <= R407;
    end
    if(T441) begin
      useRAS_2 <= R407;
    end
    if(T447) begin
      useRAS_1 <= R407;
    end
    if(T452) begin
      useRAS_0 <= R407;
    end
    if (R7)
      brIdx[T42] <= 1'h0;
  end
endmodule

module FlowThroughSerializer(
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_addr_beat,
    input [127:0] io_in_bits_data,
    input  io_in_bits_client_xact_id,
    input [2:0] io_in_bits_manager_xact_id,
    input  io_in_bits_is_builtin_type,
    input [3:0] io_in_bits_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output io_out_bits_client_xact_id,
    output[2:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output io_cnt,
    output io_done
);



  assign io_done = 1'h1;
  assign io_cnt = 1'h0;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_valid = io_in_valid;
  assign io_in_ready = io_out_ready;
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [11:0] io_req_bits_idx,
    input [19:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type
);

  wire[16:0] T0;
  wire[2:0] T1;
  wire T2;
  wire[127:0] T3;
  wire[1:0] T4;
  wire T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] s2_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [11:0] s1_pgoff;
  wire[11:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s2_miss;
  wire T14;
  wire s2_any_tag_hit;
  wire T15;
  wire T16;
  wire s2_disparity_0;
  wire T17;
  reg  R18;
  wire T19;
  wire T20;
  wire T21;
  wire stall;
  wire T22;
  reg  s1_valid;
  wire T124;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  reg  R28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37_1;
  wire[5:0] T38;
  wire T39;
  reg [63:0] vb_array;
  wire[63:0] T125;
  wire[127:0] T126;
  wire[127:0] T40;
  wire[127:0] T41;
  wire[127:0] T42;
  wire[127:0] T127;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[6:0] T46;
  wire[5:0] s2_idx;
  wire[127:0] T128;
  wire T47;
  wire[127:0] T48;
  wire[127:0] T49;
  wire[127:0] T129;
  wire T50;
  wire T51;
  reg  invalidated;
  wire T52;
  wire T53;
  wire T54;
  reg [1:0] state;
  wire[1:0] T130;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire refill_done;
  wire refill_wrap;
  wire T66;
  reg [1:0] refill_cnt;
  wire[1:0] T131;
  wire[1:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire[127:0] T71;
  wire[127:0] T72;
  wire[127:0] T73;
  wire[6:0] T74;
  wire[127:0] T132;
  wire T75;
  wire[127:0] T76;
  wire[127:0] T77;
  wire[127:0] T133;
  wire T78;
  wire T79;
  wire s2_tag_hit_0;
  wire T80;
  reg  R81;
  wire T82;
  wire s1_tag_match_0;
  wire T83;
  wire[19:0] s1_tag;
  wire[19:0] T84;
  wire[19:0] T85;
  wire[19:0] tag_rdata;
  wire T94;
  wire s0_valid;
  wire T95;
  wire T96;
  wire[5:0] T92;
  wire[11:0] s0_pgoff;
  wire T93;
  wire[19:0] T87;
  wire[19:0] T88;
  wire[19:0] T89;
  wire[19:0] s2_tag;
  reg [5:0] R90;
  wire[5:0] T91;
  reg  s2_valid;
  wire T134;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  reg [127:0] s2_dout_0;
  wire[127:0] T107;
  wire[127:0] T108;
  wire T116;
  wire T117;
  wire[7:0] T115;
  wire[127:0] T110;
  wire[127:0] T111;
  wire[7:0] T112;
  reg [7:0] R113;
  wire[7:0] T114;
  wire T118;
  wire T119;
  wire T120;
  wire[31:0] s2_dout_word_0;
  wire[127:0] T121;
  wire[6:0] T122;
  wire[1:0] T123;
  wire[5:0] s2_offset;
  wire s2_hit;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R18 = {1{$random}};
    s1_valid = {1{$random}};
    R28 = {1{$random}};
    vb_array = {2{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    refill_cnt = {1{$random}};
    R81 = {1{$random}};
    R90 = {1{$random}};
    s2_valid = {1{$random}};
    s2_dout_0 = {4{$random}};
    R113 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_union = T0;
  assign T0 = 17'h1c1;
  assign io_mem_acquire_bits_a_type = T1;
  assign T1 = 3'h1;
  assign io_mem_acquire_bits_is_builtin_type = T2;
  assign T2 = 1'h1;
  assign io_mem_acquire_bits_data = T3;
  assign T3 = 128'h0;
  assign io_mem_acquire_bits_addr_beat = T4;
  assign T4 = 2'h0;
  assign io_mem_acquire_bits_client_xact_id = T5;
  assign T5 = 1'h0;
  assign io_mem_acquire_bits_addr_block = T6;
  assign T6 = T7;
  assign T7 = s2_addr >> 3'h6;
  assign T8 = T103 ? s1_addr : s2_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T102 & T13;
  assign T13 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T14;
  assign T14 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T15;
  assign T15 = s2_tag_hit_0 & T16;
  assign T16 = s2_disparity_0 ^ 1'h1;
  assign s2_disparity_0 = T17;
  assign T17 = R28 & R18;
  assign T19 = T20 ? 1'h0 : R18;
  assign T20 = T22 & T21;
  assign T21 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T22 = s1_valid & rdy;
  assign T124 = reset ? 1'h0 : T23;
  assign T23 = T27 | T24;
  assign T24 = T26 & T25;
  assign T25 = io_req_bits_kill ^ 1'h1;
  assign T26 = s1_valid & stall;
  assign T27 = io_req_valid & rdy;
  assign T29 = T20 ? T30 : R28;
  assign T30 = T79 & T31;
  assign T31 = T32;
  assign T32 = T39 & T33;
  assign T33 = T34 - 1'h1;
  assign T34 = 1'h1 << T35;
  assign T35 = T36 + 7'h1;
  assign T36 = T37_1 - T37_1;
  assign T37_1 = {1'h0, T38};
  assign T38 = s1_pgoff[4'hb:3'h6];
  assign T39 = vb_array >> T37_1;
  assign T125 = T126[6'h3f:1'h0];
  assign T126 = reset ? 128'h0 : T40;
  assign T40 = T78 ? T71 : T41;
  assign T41 = io_invalidate ? 128'h0 : T42;
  assign T42 = T50 ? T43 : T127;
  assign T127 = {64'h0, vb_array};
  assign T43 = T48 | T44;
  assign T44 = T128 & T45;
  assign T45 = 1'h1 << T46;
  assign T46 = {1'h0, s2_idx};
  assign s2_idx = s2_addr[4'hb:3'h6];
  assign T128 = T47 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T47 = 1'h1;
  assign T48 = T129 & T49;
  assign T49 = ~ T45;
  assign T129 = {64'h0, vb_array};
  assign T50 = refill_done & T51;
  assign T51 = invalidated ^ 1'h1;
  assign T52 = T54 ? 1'h0 : T53;
  assign T53 = io_invalidate ? 1'h1 : invalidated;
  assign T54 = 2'h0 == state;
  assign T130 = reset ? 2'h0 : T55;
  assign T55 = T64 ? 2'h0 : T56;
  assign T56 = T62 ? 2'h3 : T57;
  assign T57 = T60 ? 2'h2 : T58;
  assign T58 = T59 ? 2'h1 : state;
  assign T59 = T54 & s2_miss;
  assign T60 = T61 & io_mem_acquire_ready;
  assign T61 = 2'h1 == state;
  assign T62 = T63 & io_mem_grant_valid;
  assign T63 = 2'h2 == state;
  assign T64 = T65 & refill_done;
  assign T65 = 2'h3 == state;
  assign refill_done = T70 & refill_wrap;
  assign refill_wrap = T69 & T66;
  assign T66 = refill_cnt == 2'h3;
  assign T131 = reset ? 2'h0 : T67;
  assign T67 = T69 ? T68 : refill_cnt;
  assign T68 = refill_cnt + 2'h1;
  assign T69 = 1'h1 & FlowThroughSerializer_io_out_valid;
  assign T70 = state == 2'h3;
  assign T71 = T76 | T72;
  assign T72 = T132 & T73;
  assign T73 = 1'h1 << T74;
  assign T74 = {1'h0, s2_idx};
  assign T132 = T75 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T75 = 1'h0;
  assign T76 = T133 & T77;
  assign T77 = ~ T73;
  assign T133 = {64'h0, vb_array};
  assign T78 = s2_valid & s2_disparity_0;
  assign T79 = io_invalidate ^ 1'h1;
  assign s2_tag_hit_0 = T80;
  assign T80 = R28 & R81;
  assign T82 = T20 ? s1_tag_match_0 : R81;
  assign s1_tag_match_0 = T83;
  assign T83 = T84 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hc];
  assign T84 = T85[5'h13:1'h0];
  assign T85 = tag_rdata[5'h13:1'h0];
  assign T94 = T96 & s0_valid;
  assign s0_valid = io_req_valid | T95;
  assign T95 = s1_valid & stall;
  assign T96 = refill_done ^ 1'h1;
  assign T92 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T93 ? s1_pgoff : io_req_bits_idx;
  assign T93 = s1_valid & stall;
  ICache_T86 T86 (
    .CLK(clk),
    .RW0A(refill_done ? s2_idx : T92),
    .RW0E(T94 || refill_done),
    .RW0W(refill_done),
    .RW0I(T89),
    .RW0M(T88),
    .RW0O(tag_rdata)
  );
  assign T88 = 20'hfffff;
  assign T89 = s2_tag;
  assign s2_tag = s2_addr[5'h1f:4'hc];
  assign T91 = T94 ? T92 : R90;
  assign T134 = reset ? 1'h0 : T97;
  assign T97 = T99 | T98;
  assign T98 = io_resp_valid & stall;
  assign T99 = T101 & T100;
  assign T100 = io_req_bits_kill ^ 1'h1;
  assign T101 = s1_valid & rdy;
  assign T102 = state == 2'h0;
  assign T103 = T105 & T104;
  assign T104 = stall ^ 1'h1;
  assign T105 = s1_valid & rdy;
  assign io_mem_acquire_valid = T106;
  assign T106 = state == 2'h1;
  assign io_resp_bits_datablock = s2_dout_0;
  assign T107 = T118 ? T108 : s2_dout_0;
  assign T116 = T117 & s0_valid;
  assign T117 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T115 = s0_pgoff[4'hb:3'h4];
  ICache_T109 T109 (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_io_out_valid ? T112 : T115),
    .RW0E(T116 || FlowThroughSerializer_io_out_valid),
    .RW0W(FlowThroughSerializer_io_out_valid),
    .RW0I(T111),
    .RW0O(T108)
  );
  assign T111 = FlowThroughSerializer_io_out_bits_data;
  assign T112 = {s2_idx, refill_cnt};
  assign T114 = T116 ? T115 : R113;
  assign T118 = T120 & T119;
  assign T119 = stall ^ 1'h1;
  assign T120 = s1_valid & rdy;
  assign io_resp_bits_data = s2_dout_word_0;
  assign s2_dout_word_0 = T121[5'h1f:1'h0];
  assign T121 = s2_dout_0 >> T122;
  assign T122 = T123 << 3'h5;
  assign T123 = s2_offset[2'h3:2'h2];
  assign s2_offset = s2_addr[3'h5:1'h0];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_out_bits_client_xact_id(  )
       //.io_out_bits_manager_xact_id(  )
       //.io_out_bits_is_builtin_type(  )
       //.io_out_bits_g_type(  )
       //.io_cnt(  )
       //.io_done(  )
  );

  always @(posedge clk) begin
    if(T103) begin
      s2_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T20) begin
      R18 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T23;
    end
    if(T20) begin
      R28 <= T30;
    end
    vb_array <= T125;
    if(T54) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T64) begin
      state <= 2'h0;
    end else if(T62) begin
      state <= 2'h3;
    end else if(T60) begin
      state <= 2'h2;
    end else if(T59) begin
      state <= 2'h1;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T69) begin
      refill_cnt <= T68;
    end
    if(T20) begin
      R81 <= s1_tag_match_0;
    end
    if(T94) begin
      R90 <= T92;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T97;
    end
    if(T118) begin
      s2_dout_0 <= T108;
    end
    if(T116) begin
      R113 <= T115;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input [3:0] io_clear_mask,
    input [33:0] io_tag,
    output io_hit,
    output[3:0] io_hits,
    output[3:0] io_valid_bits,
    input  io_write,
    input [33:0] io_write_tag,
    input [1:0] io_write_addr
);

  reg [3:0] vb_array;
  wire[3:0] T28;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T29;
  wire T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[1:0] T12;
  wire hits_0;
  wire T13;
  wire[33:0] T14;
  reg [33:0] cam_tags [3:0];
  wire[33:0] T15;
  wire T16;
  wire hits_1;
  wire T17;
  wire[33:0] T18;
  wire T19;
  wire[1:0] T20;
  wire hits_2;
  wire T21;
  wire[33:0] T22;
  wire T23;
  wire hits_3;
  wire T24;
  wire[33:0] T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_valid_bits = vb_array;
  assign T28 = reset ? 4'h0 : T0;
  assign T0 = io_clear ? T8 : T1;
  assign T1 = io_write ? T2 : vb_array;
  assign T2 = T6 | T3;
  assign T3 = T29 & T4;
  assign T4 = 1'h1 << io_write_addr;
  assign T29 = T5 ? 4'hf : 4'h0;
  assign T5 = 1'h1;
  assign T6 = vb_array & T7;
  assign T7 = ~ T4;
  assign T8 = vb_array & T9;
  assign T9 = ~ io_clear_mask;
  assign io_hits = T10;
  assign T10 = T11;
  assign T11 = {T20, T12};
  assign T12 = {hits_1, hits_0};
  assign hits_0 = T16 & T13;
  assign T13 = T14 == io_tag;
  assign T14 = cam_tags[2'h0];
  assign T16 = vb_array[1'h0:1'h0];
  assign hits_1 = T19 & T17;
  assign T17 = T18 == io_tag;
  assign T18 = cam_tags[2'h1];
  assign T19 = vb_array[1'h1:1'h1];
  assign T20 = {hits_3, hits_2};
  assign hits_2 = T23 & T21;
  assign T21 = T22 == io_tag;
  assign T22 = cam_tags[2'h2];
  assign T23 = vb_array[2'h2:2'h2];
  assign hits_3 = T26 & T24;
  assign T24 = T25 == io_tag;
  assign T25 = cam_tags[2'h3];
  assign T26 = vb_array[2'h3:2'h3];
  assign io_hit = T27;
  assign T27 = io_hits != 4'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 4'h0;
    end else if(io_clear) begin
      vb_array <= T8;
    end else if(io_write) begin
      vb_array <= T2;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [27:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    input  io_req_bits_store,
    output io_resp_miss,
    output[19:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    output[3:0] io_resp_hit_idx,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate
);

  reg [1:0] r_refill_waddr;
  wire[1:0] T0;
  wire[1:0] repl_waddr;
  wire[1:0] T1;
  wire[2:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  reg [3:0] R9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[6:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T287;
  wire T288;
  wire[1:0] T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire T292;
  wire T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire T24;
  wire tlb_hit;
  wire tag_hit;
  wire[3:0] tag_hits;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] w_array;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[1:0] T30;
  reg  uw_array_0;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[3:0] T42;
  wire[1:0] T43;
  reg  uw_array_1;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  reg  uw_array_2;
  wire T48;
  wire T49;
  wire T50;
  reg  uw_array_3;
  wire T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[1:0] T56;
  reg  sw_array_0;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[1:0] T67;
  reg  sw_array_1;
  wire T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  reg  sw_array_2;
  wire T72;
  wire T73;
  wire T74;
  reg  sw_array_3;
  wire T75;
  wire T76;
  wire T77;
  wire priv_s;
  wire[1:0] priv;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[1:0] T82;
  reg  dirty_array_0;
  wire T83;
  wire T84;
  wire T85;
  wire[3:0] T86;
  wire[1:0] T87;
  reg  dirty_array_1;
  wire T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  reg  dirty_array_2;
  wire T92;
  wire T93;
  wire T94;
  reg  dirty_array_3;
  wire T95;
  wire T96;
  wire T97;
  wire vm_enabled;
  wire priv_uses_vm;
  wire T98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T293;
  wire[1:0] T294;
  wire[1:0] T295;
  wire T296;
  wire[3:0] T101;
  wire T297;
  wire T298;
  wire has_invalid_entry;
  wire T102;
  wire T103;
  wire tlb_miss;
  wire T104;
  wire bad_va;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[33:0] T299;
  reg [34:0] r_refill_tag;
  wire[34:0] T110;
  wire[34:0] lookup_tag;
  wire[34:0] T111;
  wire T112;
  wire T113;
  reg [1:0] state;
  wire[1:0] T300;
  wire[1:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[33:0] T301;
  wire[3:0] T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[3:0] T132;
  wire[1:0] T133;
  reg  valid_array_0;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire[3:0] T138;
  wire[1:0] T139;
  reg  valid_array_1;
  wire T140;
  wire T141;
  wire T142;
  wire[1:0] T143;
  reg  valid_array_2;
  wire T144;
  wire T145;
  wire T146;
  reg  valid_array_3;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  reg  r_req_instruction;
  wire T152;
  reg  r_req_store;
  wire T153;
  wire[26:0] T302;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[3:0] x_array;
  wire[3:0] T160;
  wire[3:0] T161;
  wire[1:0] T162;
  reg  ux_array_0;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire[3:0] T174;
  wire[1:0] T175;
  reg  ux_array_1;
  wire T176;
  wire T177;
  wire T178;
  wire[1:0] T179;
  reg  ux_array_2;
  wire T180;
  wire T181;
  wire T182;
  reg  ux_array_3;
  wire T183;
  wire T184;
  wire T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[1:0] T188;
  reg  sx_array_0;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[3:0] T198;
  wire[1:0] T199;
  reg  sx_array_1;
  wire T200;
  wire T201;
  wire T202;
  wire[1:0] T203;
  reg  sx_array_2;
  wire T204;
  wire T205;
  wire T206;
  reg  sx_array_3;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire[3:0] T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] r_array;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[1:0] T222;
  reg  ur_array_0;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[3:0] T232;
  wire[1:0] T233;
  reg  ur_array_1;
  wire T234;
  wire T235;
  wire T236;
  wire[1:0] T237;
  reg  ur_array_2;
  wire T238;
  wire T239;
  wire T240;
  reg  ur_array_3;
  wire T241;
  wire T242;
  wire T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[1:0] T246;
  reg  sr_array_0;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire[3:0] T254;
  wire[1:0] T255;
  reg  sr_array_1;
  wire T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  reg  sr_array_2;
  wire T260;
  wire T261;
  wire T262;
  reg  sr_array_3;
  wire T263;
  wire T264;
  wire T265;
  wire[19:0] T266;
  wire[19:0] T267;
  wire[19:0] T268;
  wire[19:0] T269;
  wire[19:0] T270;
  reg [19:0] tag_ram [3:0];
  wire[19:0] T271;
  wire T272;
  wire[19:0] T273;
  wire[19:0] T274;
  wire[19:0] T275;
  wire T276;
  wire[19:0] T277;
  wire[19:0] T278;
  wire[19:0] T279;
  wire T280;
  wire[19:0] T281;
  wire[19:0] T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire[3:0] tag_cam_io_hits;
  wire[3:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R9 = {1{$random}};
    uw_array_0 = {1{$random}};
    uw_array_1 = {1{$random}};
    uw_array_2 = {1{$random}};
    uw_array_3 = {1{$random}};
    sw_array_0 = {1{$random}};
    sw_array_1 = {1{$random}};
    sw_array_2 = {1{$random}};
    sw_array_3 = {1{$random}};
    dirty_array_0 = {1{$random}};
    dirty_array_1 = {1{$random}};
    dirty_array_2 = {1{$random}};
    dirty_array_3 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    valid_array_0 = {1{$random}};
    valid_array_1 = {1{$random}};
    valid_array_2 = {1{$random}};
    valid_array_3 = {1{$random}};
    r_req_instruction = {1{$random}};
    r_req_store = {1{$random}};
    ux_array_0 = {1{$random}};
    ux_array_1 = {1{$random}};
    ux_array_2 = {1{$random}};
    ux_array_3 = {1{$random}};
    sx_array_0 = {1{$random}};
    sx_array_1 = {1{$random}};
    sx_array_2 = {1{$random}};
    sx_array_3 = {1{$random}};
    ur_array_0 = {1{$random}};
    ur_array_1 = {1{$random}};
    ur_array_2 = {1{$random}};
    ur_array_3 = {1{$random}};
    sr_array_0 = {1{$random}};
    sr_array_1 = {1{$random}};
    sr_array_2 = {1{$random}};
    sr_array_3 = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T103 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T293 : T1;
  assign T1 = T2[1'h1:1'h0];
  assign T2 = {T99, T3};
  assign T3 = T8 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 2'h1;
  assign T7 = T99 - T99;
  assign T8 = R9 >> T99;
  assign T10 = T24 ? T11 : R9;
  assign T11 = T19 | T12;
  assign T12 = T18 ? 4'h0 : T13;
  assign T13 = T14[2'h3:1'h0];
  assign T14 = 4'h1 << T15;
  assign T15 = {1'h1, T16};
  assign T16 = T287[1'h1:1'h1];
  assign T287 = {T292, T288};
  assign T288 = T289[1'h1:1'h1];
  assign T289 = T291 | T290;
  assign T290 = tag_cam_io_hits[1'h1:1'h0];
  assign T291 = tag_cam_io_hits[2'h3:2'h2];
  assign T292 = T291 != 2'h0;
  assign T18 = T287[1'h0:1'h0];
  assign T19 = T21 & T20;
  assign T20 = ~ T13;
  assign T21 = T23 | T22;
  assign T22 = T16 ? 4'h0 : 4'h2;
  assign T23 = R9 & 4'hd;
  assign T24 = io_req_valid & tlb_hit;
  assign tlb_hit = vm_enabled & tag_hit;
  assign tag_hit = tag_hits != 4'h0;
  assign tag_hits = tag_cam_io_hits & T25;
  assign T25 = T80 | T26;
  assign T26 = ~ T27;
  assign T27 = io_req_bits_store ? w_array : 4'h0;
  assign w_array = priv_s ? T54 : T28;
  assign T28 = T29;
  assign T29 = {T47, T30};
  assign T30 = {uw_array_1, uw_array_0};
  assign T31 = T40 ? T32 : uw_array_0;
  assign T32 = T34 & T33;
  assign T33 = io_ptw_resp_bits_error ^ 1'h1;
  assign T34 = T36 & T35;
  assign T35 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T36 = T38 & T37;
  assign T37 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T38 = io_ptw_resp_bits_pte_v & T39;
  assign T39 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T40 = io_ptw_resp_valid & T41;
  assign T41 = T42[1'h0:1'h0];
  assign T42 = 1'h1 << T43;
  assign T43 = r_refill_waddr;
  assign T44 = T45 ? T32 : uw_array_1;
  assign T45 = io_ptw_resp_valid & T46;
  assign T46 = T42[1'h1:1'h1];
  assign T47 = {uw_array_3, uw_array_2};
  assign T48 = T49 ? T32 : uw_array_2;
  assign T49 = io_ptw_resp_valid & T50;
  assign T50 = T42[2'h2:2'h2];
  assign T51 = T52 ? T32 : uw_array_3;
  assign T52 = io_ptw_resp_valid & T53;
  assign T53 = T42[2'h3:2'h3];
  assign T54 = T55;
  assign T55 = {T71, T56};
  assign T56 = {sw_array_1, sw_array_0};
  assign T57 = T64 ? T58 : sw_array_0;
  assign T58 = T60 & T59;
  assign T59 = io_ptw_resp_bits_error ^ 1'h1;
  assign T60 = T62 & T61;
  assign T61 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T62 = io_ptw_resp_bits_pte_v & T63;
  assign T63 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T64 = io_ptw_resp_valid & T65;
  assign T65 = T66[1'h0:1'h0];
  assign T66 = 1'h1 << T67;
  assign T67 = r_refill_waddr;
  assign T68 = T69 ? T58 : sw_array_1;
  assign T69 = io_ptw_resp_valid & T70;
  assign T70 = T66[1'h1:1'h1];
  assign T71 = {sw_array_3, sw_array_2};
  assign T72 = T73 ? T58 : sw_array_2;
  assign T73 = io_ptw_resp_valid & T74;
  assign T74 = T66[2'h2:2'h2];
  assign T75 = T76 ? T58 : sw_array_3;
  assign T76 = io_ptw_resp_valid & T77;
  assign T77 = T66[2'h3:2'h3];
  assign priv_s = priv == 2'h1;
  assign priv = T78 ? io_ptw_status_prv1 : io_ptw_status_prv;
  assign T78 = io_ptw_status_mprv & T79;
  assign T79 = io_req_bits_instruction ^ 1'h1;
  assign T80 = T81;
  assign T81 = {T91, T82};
  assign T82 = {dirty_array_1, dirty_array_0};
  assign T83 = T84 ? io_ptw_resp_bits_pte_d : dirty_array_0;
  assign T84 = io_ptw_resp_valid & T85;
  assign T85 = T86[1'h0:1'h0];
  assign T86 = 1'h1 << T87;
  assign T87 = r_refill_waddr;
  assign T88 = T89 ? io_ptw_resp_bits_pte_d : dirty_array_1;
  assign T89 = io_ptw_resp_valid & T90;
  assign T90 = T86[1'h1:1'h1];
  assign T91 = {dirty_array_3, dirty_array_2};
  assign T92 = T93 ? io_ptw_resp_bits_pte_d : dirty_array_2;
  assign T93 = io_ptw_resp_valid & T94;
  assign T94 = T86[2'h2:2'h2];
  assign T95 = T96 ? io_ptw_resp_bits_pte_d : dirty_array_3;
  assign T96 = io_ptw_resp_valid & T97;
  assign T97 = T86[2'h3:2'h3];
  assign vm_enabled = T98 & priv_uses_vm;
  assign priv_uses_vm = priv <= 2'h1;
  assign T98 = io_ptw_status_vm[2'h3:2'h3];
  assign T99 = {1'h1, T100};
  assign T100 = R9[1'h1:1'h1];
  assign T293 = T298 ? 1'h0 : T294;
  assign T294 = T297 ? 1'h1 : T295;
  assign T295 = T296 ? 2'h2 : 2'h3;
  assign T296 = T101[2'h2:2'h2];
  assign T101 = ~ tag_cam_io_valid_bits;
  assign T297 = T101[1'h1:1'h1];
  assign T298 = T101[1'h0:1'h0];
  assign has_invalid_entry = T102 ^ 1'h1;
  assign T102 = tag_cam_io_valid_bits == 4'hf;
  assign T103 = T109 & tlb_miss;
  assign tlb_miss = T107 & T104;
  assign T104 = bad_va ^ 1'h1;
  assign bad_va = T106 != T105;
  assign T105 = io_req_bits_vpn[5'h1a:5'h1a];
  assign T106 = io_req_bits_vpn[5'h1b:5'h1b];
  assign T107 = vm_enabled & T108;
  assign T108 = tag_hit ^ 1'h1;
  assign T109 = io_req_ready & io_req_valid;
  assign T299 = r_refill_tag[6'h21:1'h0];
  assign T110 = T103 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T111;
  assign T111 = {io_req_bits_asid, io_req_bits_vpn};
  assign T112 = T113 & io_ptw_resp_valid;
  assign T113 = state == 2'h2;
  assign T300 = reset ? 2'h0 : T114;
  assign T114 = io_ptw_resp_valid ? 2'h0 : T115;
  assign T115 = T124 ? 2'h3 : T116;
  assign T116 = T123 ? 2'h3 : T117;
  assign T117 = T122 ? 2'h2 : T118;
  assign T118 = T120 ? 2'h0 : T119;
  assign T119 = T103 ? 2'h1 : state;
  assign T120 = T121 & io_ptw_invalidate;
  assign T121 = state == 2'h1;
  assign T122 = T121 & io_ptw_req_ready;
  assign T123 = T122 & io_ptw_invalidate;
  assign T124 = T125 & io_ptw_invalidate;
  assign T125 = state == 2'h2;
  assign T301 = lookup_tag[6'h21:1'h0];
  assign T126 = io_ptw_invalidate ? 4'hf : T127;
  assign T127 = T130 | T128;
  assign T128 = tag_cam_io_hits & T129;
  assign T129 = ~ tag_hits;
  assign T130 = ~ T131;
  assign T131 = T132;
  assign T132 = {T143, T133};
  assign T133 = {valid_array_1, valid_array_0};
  assign T134 = T136 ? T135 : valid_array_0;
  assign T135 = io_ptw_resp_bits_error ^ 1'h1;
  assign T136 = io_ptw_resp_valid & T137;
  assign T137 = T138[1'h0:1'h0];
  assign T138 = 1'h1 << T139;
  assign T139 = r_refill_waddr;
  assign T140 = T141 ? T135 : valid_array_1;
  assign T141 = io_ptw_resp_valid & T142;
  assign T142 = T138[1'h1:1'h1];
  assign T143 = {valid_array_3, valid_array_2};
  assign T144 = T145 ? T135 : valid_array_2;
  assign T145 = io_ptw_resp_valid & T146;
  assign T146 = T138[2'h2:2'h2];
  assign T147 = T148 ? T135 : valid_array_3;
  assign T148 = io_ptw_resp_valid & T149;
  assign T149 = T138[2'h3:2'h3];
  assign T150 = io_ptw_invalidate | T151;
  assign T151 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T152 = T103 ? io_req_bits_instruction : r_req_instruction;
  assign io_ptw_req_bits_store = r_req_store;
  assign T153 = T103 ? io_req_bits_store : r_req_store;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_addr = T302;
  assign T302 = r_refill_tag[5'h1a:1'h0];
  assign io_ptw_req_valid = T154;
  assign T154 = state == 2'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_xcpt_if = T155;
  assign T155 = bad_va | T156;
  assign T156 = tlb_hit & T157;
  assign T157 = T158 ^ 1'h1;
  assign T158 = T159 != 4'h0;
  assign T159 = x_array & tag_cam_io_hits;
  assign x_array = priv_s ? T186 : T160;
  assign T160 = T161;
  assign T161 = {T179, T162};
  assign T162 = {ux_array_1, ux_array_0};
  assign T163 = T172 ? T164 : ux_array_0;
  assign T164 = T166 & T165;
  assign T165 = io_ptw_resp_bits_error ^ 1'h1;
  assign T166 = T168 & T167;
  assign T167 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T168 = T170 & T169;
  assign T169 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T170 = io_ptw_resp_bits_pte_v & T171;
  assign T171 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T172 = io_ptw_resp_valid & T173;
  assign T173 = T174[1'h0:1'h0];
  assign T174 = 1'h1 << T175;
  assign T175 = r_refill_waddr;
  assign T176 = T177 ? T164 : ux_array_1;
  assign T177 = io_ptw_resp_valid & T178;
  assign T178 = T174[1'h1:1'h1];
  assign T179 = {ux_array_3, ux_array_2};
  assign T180 = T181 ? T164 : ux_array_2;
  assign T181 = io_ptw_resp_valid & T182;
  assign T182 = T174[2'h2:2'h2];
  assign T183 = T184 ? T164 : ux_array_3;
  assign T184 = io_ptw_resp_valid & T185;
  assign T185 = T174[2'h3:2'h3];
  assign T186 = T187;
  assign T187 = {T203, T188};
  assign T188 = {sx_array_1, sx_array_0};
  assign T189 = T196 ? T190 : sx_array_0;
  assign T190 = T192 & T191;
  assign T191 = io_ptw_resp_bits_error ^ 1'h1;
  assign T192 = T194 & T193;
  assign T193 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T194 = io_ptw_resp_bits_pte_v & T195;
  assign T195 = 4'h4 <= io_ptw_resp_bits_pte_typ;
  assign T196 = io_ptw_resp_valid & T197;
  assign T197 = T198[1'h0:1'h0];
  assign T198 = 1'h1 << T199;
  assign T199 = r_refill_waddr;
  assign T200 = T201 ? T190 : sx_array_1;
  assign T201 = io_ptw_resp_valid & T202;
  assign T202 = T198[1'h1:1'h1];
  assign T203 = {sx_array_3, sx_array_2};
  assign T204 = T205 ? T190 : sx_array_2;
  assign T205 = io_ptw_resp_valid & T206;
  assign T206 = T198[2'h2:2'h2];
  assign T207 = T208 ? T190 : sx_array_3;
  assign T208 = io_ptw_resp_valid & T209;
  assign T209 = T198[2'h3:2'h3];
  assign io_resp_xcpt_st = T210;
  assign T210 = bad_va | T211;
  assign T211 = tlb_hit & T212;
  assign T212 = T213 ^ 1'h1;
  assign T213 = T214 != 4'h0;
  assign T214 = w_array & tag_cam_io_hits;
  assign io_resp_xcpt_ld = T215;
  assign T215 = bad_va | T216;
  assign T216 = tlb_hit & T217;
  assign T217 = T218 ^ 1'h1;
  assign T218 = T219 != 4'h0;
  assign T219 = r_array & tag_cam_io_hits;
  assign r_array = priv_s ? T244 : T220;
  assign T220 = T221;
  assign T221 = {T237, T222};
  assign T222 = {ur_array_1, ur_array_0};
  assign T223 = T230 ? T224 : ur_array_0;
  assign T224 = T226 & T225;
  assign T225 = io_ptw_resp_bits_error ^ 1'h1;
  assign T226 = T228 & T227;
  assign T227 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T228 = io_ptw_resp_bits_pte_v & T229;
  assign T229 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T230 = io_ptw_resp_valid & T231;
  assign T231 = T232[1'h0:1'h0];
  assign T232 = 1'h1 << T233;
  assign T233 = r_refill_waddr;
  assign T234 = T235 ? T224 : ur_array_1;
  assign T235 = io_ptw_resp_valid & T236;
  assign T236 = T232[1'h1:1'h1];
  assign T237 = {ur_array_3, ur_array_2};
  assign T238 = T239 ? T224 : ur_array_2;
  assign T239 = io_ptw_resp_valid & T240;
  assign T240 = T232[2'h2:2'h2];
  assign T241 = T242 ? T224 : ur_array_3;
  assign T242 = io_ptw_resp_valid & T243;
  assign T243 = T232[2'h3:2'h3];
  assign T244 = T245;
  assign T245 = {T259, T246};
  assign T246 = {sr_array_1, sr_array_0};
  assign T247 = T252 ? T248 : sr_array_0;
  assign T248 = T250 & T249;
  assign T249 = io_ptw_resp_bits_error ^ 1'h1;
  assign T250 = io_ptw_resp_bits_pte_v & T251;
  assign T251 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T252 = io_ptw_resp_valid & T253;
  assign T253 = T254[1'h0:1'h0];
  assign T254 = 1'h1 << T255;
  assign T255 = r_refill_waddr;
  assign T256 = T257 ? T248 : sr_array_1;
  assign T257 = io_ptw_resp_valid & T258;
  assign T258 = T254[1'h1:1'h1];
  assign T259 = {sr_array_3, sr_array_2};
  assign T260 = T261 ? T248 : sr_array_2;
  assign T261 = io_ptw_resp_valid & T262;
  assign T262 = T254[2'h2:2'h2];
  assign T263 = T264 ? T248 : sr_array_3;
  assign T264 = io_ptw_resp_valid & T265;
  assign T265 = T254[2'h3:2'h3];
  assign io_resp_ppn = T266;
  assign T266 = T284 ? T268 : T267;
  assign T267 = io_req_bits_vpn[5'h13:1'h0];
  assign T268 = T273 | T269;
  assign T269 = T272 ? T270 : 20'h0;
  assign T270 = tag_ram[2'h3];
  assign T272 = tag_cam_io_hits[2'h3:2'h3];
  assign T273 = T277 | T274;
  assign T274 = T276 ? T275 : 20'h0;
  assign T275 = tag_ram[2'h2];
  assign T276 = tag_cam_io_hits[2'h2:2'h2];
  assign T277 = T281 | T278;
  assign T278 = T280 ? T279 : 20'h0;
  assign T279 = tag_ram[2'h1];
  assign T280 = tag_cam_io_hits[1'h1:1'h1];
  assign T281 = T283 ? T282 : 20'h0;
  assign T282 = tag_ram[2'h0];
  assign T283 = tag_cam_io_hits[1'h0:1'h0];
  assign T284 = vm_enabled & T285;
  assign T285 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T286;
  assign T286 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( T150 ),
       .io_clear_mask( T126 ),
       .io_tag( T301 ),
       //.io_hit(  )
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T112 ),
       .io_write_tag( T299 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T103) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T24) begin
      R9 <= T11;
    end
    if(T40) begin
      uw_array_0 <= T32;
    end
    if(T45) begin
      uw_array_1 <= T32;
    end
    if(T49) begin
      uw_array_2 <= T32;
    end
    if(T52) begin
      uw_array_3 <= T32;
    end
    if(T64) begin
      sw_array_0 <= T58;
    end
    if(T69) begin
      sw_array_1 <= T58;
    end
    if(T73) begin
      sw_array_2 <= T58;
    end
    if(T76) begin
      sw_array_3 <= T58;
    end
    if(T84) begin
      dirty_array_0 <= io_ptw_resp_bits_pte_d;
    end
    if(T89) begin
      dirty_array_1 <= io_ptw_resp_bits_pte_d;
    end
    if(T93) begin
      dirty_array_2 <= io_ptw_resp_bits_pte_d;
    end
    if(T96) begin
      dirty_array_3 <= io_ptw_resp_bits_pte_d;
    end
    if(T103) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T124) begin
      state <= 2'h3;
    end else if(T123) begin
      state <= 2'h3;
    end else if(T122) begin
      state <= 2'h2;
    end else if(T120) begin
      state <= 2'h0;
    end else if(T103) begin
      state <= 2'h1;
    end
    if(T136) begin
      valid_array_0 <= T135;
    end
    if(T141) begin
      valid_array_1 <= T135;
    end
    if(T145) begin
      valid_array_2 <= T135;
    end
    if(T148) begin
      valid_array_3 <= T135;
    end
    if(T103) begin
      r_req_instruction <= io_req_bits_instruction;
    end
    if(T103) begin
      r_req_store <= io_req_bits_store;
    end
    if(T172) begin
      ux_array_0 <= T164;
    end
    if(T177) begin
      ux_array_1 <= T164;
    end
    if(T181) begin
      ux_array_2 <= T164;
    end
    if(T184) begin
      ux_array_3 <= T164;
    end
    if(T196) begin
      sx_array_0 <= T190;
    end
    if(T201) begin
      sx_array_1 <= T190;
    end
    if(T205) begin
      sx_array_2 <= T190;
    end
    if(T208) begin
      sx_array_3 <= T190;
    end
    if(T230) begin
      ur_array_0 <= T224;
    end
    if(T235) begin
      ur_array_1 <= T224;
    end
    if(T239) begin
      ur_array_2 <= T224;
    end
    if(T242) begin
      ur_array_3 <= T224;
    end
    if(T252) begin
      sr_array_0 <= T248;
    end
    if(T257) begin
      sr_array_1 <= T248;
    end
    if(T261) begin
      sr_array_2 <= T248;
    end
    if(T264) begin
      sr_array_3 <= T248;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_pte_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data_0,
    output io_cpu_resp_bits_mask,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output io_cpu_btb_resp_bits_mask,
    output io_cpu_btb_resp_bits_bridx,
    output[38:0] io_cpu_btb_resp_bits_target,
    output[2:0] io_cpu_btb_resp_bits_entry,
    output[3:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input  io_cpu_btb_update_bits_prediction_bits_mask,
    input  io_cpu_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [2:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_btb_update_bits_pc,
    input [38:0] io_cpu_btb_update_bits_target,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isReturn,
    input [38:0] io_cpu_btb_update_bits_br_pc,
    input  io_cpu_bht_update_valid,
    input  io_cpu_bht_update_bits_prediction_valid,
    input  io_cpu_bht_update_bits_prediction_bits_taken,
    input  io_cpu_bht_update_bits_prediction_bits_mask,
    input  io_cpu_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_bht_update_bits_prediction_bits_target,
    input [2:0] io_cpu_bht_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_bht_update_bits_pc,
    input  io_cpu_bht_update_bits_taken,
    input  io_cpu_bht_update_bits_mispredict,
    input  io_cpu_ras_update_valid,
    input  io_cpu_ras_update_bits_isCall,
    input  io_cpu_ras_update_bits_isReturn,
    input [38:0] io_cpu_ras_update_bits_returnAddr,
    input  io_cpu_ras_update_bits_prediction_valid,
    input  io_cpu_ras_update_bits_prediction_bits_taken,
    input  io_cpu_ras_update_bits_prediction_bits_mask,
    input  io_cpu_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_ras_update_bits_prediction_bits_target,
    input [2:0] io_cpu_ras_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
    input  io_cpu_invalidate,
    output[39:0] io_cpu_npc,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type
);

  wire[27:0] T0;
  wire[39:0] s1_pc;
  wire[39:0] T1;
  wire[39:0] T2;
  reg [39:0] s1_pc_;
  wire[39:0] T3;
  wire[39:0] T4;
  wire[39:0] npc;
  wire[39:0] T5;
  wire[39:0] predicted_npc;
  wire[39:0] ntpc;
  wire[38:0] T6;
  wire[36:0] T7;
  wire[39:0] ntpc_0;
  wire T8;
  wire T9;
  wire T10;
  wire[39:0] btbTarget;
  wire T11;
  reg [39:0] s2_pc;
  wire[39:0] T67;
  wire[39:0] T12;
  wire T13;
  wire T14;
  wire icmiss;
  wire T15;
  reg  s2_valid;
  wire T68;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire stall;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  s1_same_block;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire s0_same_block;
  wire T30;
  wire[39:0] T31;
  wire[39:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[11:0] T69;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[38:0] T70;
  wire T46;
  wire T47;
  wire T48;
  wire[39:0] T49;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T50;
  wire T51;
  reg [3:0] s2_btb_resp_bits_bht_history;
  wire[3:0] T52;
  reg [2:0] s2_btb_resp_bits_entry;
  wire[2:0] T53;
  reg [38:0] s2_btb_resp_bits_target;
  wire[38:0] T54;
  reg  s2_btb_resp_bits_bridx;
  wire T55;
  reg  s2_btb_resp_bits_mask;
  wire T56;
  reg  s2_btb_resp_bits_taken;
  wire T57;
  reg  s2_btb_resp_valid;
  wire T71;
  wire T58;
  reg  s2_xcpt_if;
  wire T72;
  wire T59;
  wire T73;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T74;
  wire[31:0] T62;
  wire[127:0] fetch_data;
  wire[6:0] T63;
  wire[1:0] T64;
  wire T65;
  wire T66;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire btb_io_resp_bits_mask;
  wire btb_io_resp_bits_bridx;
  wire[38:0] btb_io_resp_bits_target;
  wire[2:0] btb_io_resp_bits_entry;
  wire[3:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire icache_io_mem_grant_ready;
  wire tlb_io_resp_miss;
  wire[19:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[26:0] tlb_io_ptw_req_bits_addr;
  wire[1:0] tlb_io_ptw_req_bits_prv;
  wire tlb_io_ptw_req_bits_store;
  wire tlb_io_ptw_req_bits_fetch;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_bridx = {1{$random}};
    s2_btb_resp_bits_mask = {1{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = s1_pc >> 4'hc;
  assign s1_pc = ~ T1;
  assign T1 = T2 | 40'h3;
  assign T2 = ~ s1_pc_;
  assign T3 = io_cpu_req_valid ? io_cpu_req_bits_pc : T4;
  assign T4 = T19 ? npc : s1_pc_;
  assign npc = T5;
  assign T5 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : ntpc;
  assign ntpc = {T8, T6};
  assign T6 = {T7, 2'h0};
  assign T7 = ntpc_0[6'h26:2'h2];
  assign ntpc_0 = s1_pc + 40'h4;
  assign T8 = T10 & T9;
  assign T9 = ntpc_0[6'h26:6'h26];
  assign T10 = s1_pc[6'h26:6'h26];
  assign btbTarget = {T11, btb_io_resp_bits_target};
  assign T11 = btb_io_resp_bits_target[6'h26:6'h26];
  assign T67 = reset ? 40'h200 : T12;
  assign T12 = T13 ? s1_pc : s2_pc;
  assign T13 = T19 & T14;
  assign T14 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T15;
  assign T15 = icache_io_resp_valid ^ 1'h1;
  assign T68 = reset ? 1'h1 : T16;
  assign T16 = io_cpu_req_valid ? 1'h0 : T17;
  assign T17 = T19 ? T18 : s2_valid;
  assign T18 = icmiss ^ 1'h1;
  assign T19 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T20;
  assign T20 = io_cpu_resp_ready ^ 1'h1;
  assign T21 = T23 & T22;
  assign T22 = icmiss ^ 1'h1;
  assign T23 = stall ^ 1'h1;
  assign T24 = T38 & T25;
  assign T25 = s1_same_block ^ 1'h1;
  assign T26 = io_cpu_req_valid ? 1'h0 : T27;
  assign T27 = T19 ? T28 : s1_same_block;
  assign T28 = s0_same_block & T29;
  assign T29 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T33 & T30;
  assign T30 = T32 == T31;
  assign T31 = s1_pc & 40'h10;
  assign T32 = ntpc & 40'h10;
  assign T33 = T35 & T34;
  assign T34 = btb_io_resp_bits_taken ^ 1'h1;
  assign T35 = T37 & T36;
  assign T36 = io_cpu_req_valid ^ 1'h1;
  assign T37 = icmiss ^ 1'h1;
  assign T38 = stall ^ 1'h1;
  assign T39 = T40 | io_ptw_invalidate;
  assign T40 = T41 | icmiss;
  assign T41 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T69 = io_cpu_npc[4'hb:1'h0];
  assign T42 = T44 & T43;
  assign T43 = s0_same_block ^ 1'h1;
  assign T44 = stall ^ 1'h1;
  assign T45 = io_cpu_invalidate | io_ptw_invalidate;
  assign T70 = s1_pc[6'h26:1'h0];
  assign T46 = T48 & T47;
  assign T47 = icmiss ^ 1'h1;
  assign T48 = stall ^ 1'h1;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_npc = T49;
  assign T49 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T50 = T51 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T51 = T13 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T52 = T51 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T53 = T51 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T54 = T51 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign T55 = T51 ? btb_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign T56 = T51 ? btb_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T57 = T51 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T71 = reset ? 1'h0 : T58;
  assign T58 = T13 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T72 = reset ? 1'h0 : T59;
  assign T59 = T13 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_mask = T73;
  assign T73 = T60[1'h0:1'h0];
  assign T60 = s2_btb_resp_valid ? T61 : 2'h3;
  assign T61 = 2'h3 & T74;
  assign T74 = {1'h0, s2_btb_resp_bits_mask};
  assign io_cpu_resp_bits_data_0 = T62;
  assign T62 = fetch_data[5'h1f:1'h0];
  assign fetch_data = icache_io_resp_bits_datablock >> T63;
  assign T63 = T64 << 3'h5;
  assign T64 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_valid = T65;
  assign T65 = s2_valid & T66;
  assign T66 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T46 ),
       .io_req_bits_addr( T70 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_mask( btb_io_resp_bits_mask ),
       .io_resp_bits_bridx( btb_io_resp_bits_bridx ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_btb_update_valid( io_cpu_btb_update_valid ),
       .io_btb_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_btb_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_btb_update_bits_prediction_bits_mask( io_cpu_btb_update_bits_prediction_bits_mask ),
       .io_btb_update_bits_prediction_bits_bridx( io_cpu_btb_update_bits_prediction_bits_bridx ),
       .io_btb_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_btb_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_btb_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_btb_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_btb_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_btb_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_btb_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_btb_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_btb_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_btb_update_bits_br_pc( io_cpu_btb_update_bits_br_pc ),
       .io_bht_update_valid( io_cpu_bht_update_valid ),
       .io_bht_update_bits_prediction_valid( io_cpu_bht_update_bits_prediction_valid ),
       .io_bht_update_bits_prediction_bits_taken( io_cpu_bht_update_bits_prediction_bits_taken ),
       .io_bht_update_bits_prediction_bits_mask( io_cpu_bht_update_bits_prediction_bits_mask ),
       .io_bht_update_bits_prediction_bits_bridx( io_cpu_bht_update_bits_prediction_bits_bridx ),
       .io_bht_update_bits_prediction_bits_target( io_cpu_bht_update_bits_prediction_bits_target ),
       .io_bht_update_bits_prediction_bits_entry( io_cpu_bht_update_bits_prediction_bits_entry ),
       .io_bht_update_bits_prediction_bits_bht_history( io_cpu_bht_update_bits_prediction_bits_bht_history ),
       .io_bht_update_bits_prediction_bits_bht_value( io_cpu_bht_update_bits_prediction_bits_bht_value ),
       .io_bht_update_bits_pc( io_cpu_bht_update_bits_pc ),
       .io_bht_update_bits_taken( io_cpu_bht_update_bits_taken ),
       .io_bht_update_bits_mispredict( io_cpu_bht_update_bits_mispredict ),
       .io_ras_update_valid( io_cpu_ras_update_valid ),
       .io_ras_update_bits_isCall( io_cpu_ras_update_bits_isCall ),
       .io_ras_update_bits_isReturn( io_cpu_ras_update_bits_isReturn ),
       .io_ras_update_bits_returnAddr( io_cpu_ras_update_bits_returnAddr ),
       .io_ras_update_bits_prediction_valid( io_cpu_ras_update_bits_prediction_valid ),
       .io_ras_update_bits_prediction_bits_taken( io_cpu_ras_update_bits_prediction_bits_taken ),
       .io_ras_update_bits_prediction_bits_mask( io_cpu_ras_update_bits_prediction_bits_mask ),
       .io_ras_update_bits_prediction_bits_bridx( io_cpu_ras_update_bits_prediction_bits_bridx ),
       .io_ras_update_bits_prediction_bits_target( io_cpu_ras_update_bits_prediction_bits_target ),
       .io_ras_update_bits_prediction_bits_entry( io_cpu_ras_update_bits_prediction_bits_entry ),
       .io_ras_update_bits_prediction_bits_bht_history( io_cpu_ras_update_bits_prediction_bits_bht_history ),
       .io_ras_update_bits_prediction_bits_bht_value( io_cpu_ras_update_bits_prediction_bits_bht_value ),
       .io_invalidate( T45 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T42 ),
       .io_req_bits_idx( T69 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T39 ),
       .io_resp_ready( T24 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T21 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T0 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_req_bits_store( 1'h0 ),
       .io_resp_miss( tlb_io_resp_miss ),
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( tlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( tlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( tlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( tlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T19) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 40'h200;
    end else if(T13) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T19) begin
      s2_valid <= T18;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T19) begin
      s1_same_block <= T28;
    end
    if(T51) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T51) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T51) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T51) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T51) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if(T51) begin
      s2_btb_resp_bits_mask <= btb_io_resp_bits_mask;
    end
    if(T51) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T13) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T13) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr_block,
    input  io_req_bits_client_xact_id,
    input [1:0] io_req_bits_addr_beat,
    input [127:0] io_req_bits_data,
    input [2:0] io_req_bits_r_type,
    input  io_req_bits_voluntary,
    input  io_req_bits_way_en,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr_block,
    output io_release_bits_client_xact_id,
    output[1:0] io_release_bits_addr_beat,
    output[127:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type,
    output io_release_bits_voluntary
);

  reg  req_voluntary;
  wire T0;
  wire T1;
  reg [2:0] req_r_type;
  wire[2:0] T2;
  reg [1:0] beat_cnt;
  wire[1:0] T40;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  reg  req_client_xact_id;
  wire T6;
  reg [25:0] req_addr_block;
  wire[25:0] T7;
  wire T8;
  reg  r2_data_req_fired;
  wire T41;
  wire T9;
  wire T10;
  reg  r1_data_req_fired;
  wire T42;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg  active;
  wire T43;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [2:0] data_req_cnt;
  wire[2:0] T44;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T45;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[11:0] T33;
  wire[7:0] T34;
  wire[1:0] T35;
  wire[5:0] req_idx;
  reg  req_way_en;
  wire T36;
  wire fire;
  wire T37;
  wire[19:0] T38;
  wire T39;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_voluntary = {1{$random}};
    req_r_type = {1{$random}};
    beat_cnt = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr_block = {1{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    data_req_cnt = {1{$random}};
    req_way_en = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_release_bits_voluntary = req_voluntary;
  assign T0 = T1 ? io_req_bits_voluntary : req_voluntary;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_r_type = req_r_type;
  assign T2 = T1 ? io_req_bits_r_type : req_r_type;
  assign io_release_bits_data = io_data_resp;
  assign io_release_bits_addr_beat = beat_cnt;
  assign T40 = reset ? 2'h0 : T3;
  assign T3 = T5 ? T4 : beat_cnt;
  assign T4 = beat_cnt + 2'h1;
  assign T5 = io_release_ready & io_release_valid;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T6 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr_block = req_addr_block;
  assign T7 = T1 ? io_req_bits_addr_block : req_addr_block;
  assign io_release_valid = T8;
  assign T8 = active & r2_data_req_fired;
  assign T41 = reset ? 1'h0 : T9;
  assign T9 = T18 ? 1'h0 : T10;
  assign T10 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T42 = reset ? 1'h0 : T11;
  assign T11 = T18 ? 1'h0 : T12;
  assign T12 = T14 ? 1'h1 : T13;
  assign T13 = active ? 1'h0 : r1_data_req_fired;
  assign T14 = active & T15;
  assign T15 = T17 & T16;
  assign T16 = io_meta_read_ready & io_meta_read_valid;
  assign T17 = io_data_req_ready & io_data_req_valid;
  assign T18 = T8 & T19;
  assign T19 = io_release_ready ^ 1'h1;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = T1 ? 1'h1 : T21;
  assign T21 = T31 ? T22 : active;
  assign T22 = T24 | T23;
  assign T23 = io_release_ready ^ 1'h1;
  assign T24 = data_req_cnt < 3'h4;
  assign T44 = reset ? 3'h0 : T25;
  assign T25 = T1 ? 3'h0 : T26;
  assign T26 = T18 ? T29 : T27;
  assign T27 = T14 ? T28 : data_req_cnt;
  assign T28 = data_req_cnt + 3'h1;
  assign T29 = data_req_cnt - T45;
  assign T45 = {1'h0, T30};
  assign T30 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign T31 = T8 & T32;
  assign T32 = r1_data_req_fired ^ 1'h1;
  assign io_data_req_bits_addr = T33;
  assign T33 = T34 << 3'h4;
  assign T34 = {req_idx, T35};
  assign T35 = data_req_cnt[1'h1:1'h0];
  assign req_idx = req_addr_block[3'h5:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T36 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T37;
  assign T37 = data_req_cnt < 3'h4;
  assign io_meta_read_bits_tag = T38;
  assign T38 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T39;
  assign T39 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_voluntary <= io_req_bits_voluntary;
    end
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(reset) begin
      beat_cnt <= 2'h0;
    end else if(T5) begin
      beat_cnt <= T4;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_addr_block <= io_req_bits_addr_block;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(T18) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T18) begin
      r1_data_req_fired <= 1'h0;
    end else if(T14) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T31) begin
      active <= T22;
    end
    if(reset) begin
      data_req_cnt <= 3'h0;
    end else if(T1) begin
      data_req_cnt <= 3'h0;
    end else if(T18) begin
      data_req_cnt <= T29;
    end else if(T14) begin
      data_req_cnt <= T28;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_p_type,
    //input  io_req_bits_client_xact_id
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr_block,
    output io_rep_bits_client_xact_id,
    output[1:0] io_rep_bits_addr_beat,
    output[127:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    output io_rep_bits_voluntary,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[25:0] io_wb_req_bits_addr_block,
    output io_wb_req_bits_client_xact_id,
    output[1:0] io_wb_req_bits_addr_beat,
    output[127:0] io_wb_req_bits_data,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output io_wb_req_bits_way_en,
    input  io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_block_state_state
);

  reg  way_en;
  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T63;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[2:0] T20;
  wire T21;
  reg [1:0] old_coh_state;
  wire[1:0] T22;
  wire T23;
  wire tag_matches;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire reply_voluntary;
  wire[2:0] reply_r_type;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  reg [1:0] req_p_type;
  wire[1:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire[127:0] reply_data;
  wire[1:0] reply_addr_beat;
  wire reply_client_xact_id;
  wire[25:0] reply_addr_block;
  reg [25:0] req_addr_block;
  wire[25:0] T44;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[19:0] T53;
  wire[5:0] T64;
  wire T54;
  wire[19:0] T55;
  wire[5:0] T65;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    way_en = {1{$random}};
    state = {1{$random}};
    old_coh_state = {1{$random}};
    req_p_type = {1{$random}};
    req_addr_block = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_wb_req_bits_way_en = way_en;
  assign T0 = T1 ? io_way_en : way_en;
  assign T1 = state == 3'h3;
  assign T63 = reset ? 3'h0 : T2;
  assign T2 = T29 ? 3'h1 : T3;
  assign T3 = T27 ? 3'h2 : T4;
  assign T4 = T26 ? 3'h3 : T5;
  assign T5 = T24 ? 3'h1 : T6;
  assign T6 = T1 ? 3'h4 : T7;
  assign T7 = T23 ? T20 : T8;
  assign T8 = T18 ? 3'h0 : T9;
  assign T9 = T16 ? 3'h6 : T10;
  assign T10 = T14 ? 3'h7 : T11;
  assign T11 = T12 ? 3'h0 : state;
  assign T12 = T13 & io_meta_write_ready;
  assign T13 = state == 3'h7;
  assign T14 = T15 & io_wb_req_ready;
  assign T15 = state == 3'h6;
  assign T16 = T17 & io_wb_req_ready;
  assign T17 = state == 3'h5;
  assign T18 = T19 & io_rep_ready;
  assign T19 = state == 3'h4;
  assign T20 = T21 ? 3'h5 : 3'h7;
  assign T21 = 2'h3 == old_coh_state;
  assign T22 = T1 ? io_block_state_state : old_coh_state;
  assign T23 = T18 & tag_matches;
  assign tag_matches = way_en != 1'h0;
  assign T24 = T1 & T25;
  assign T25 = io_mshr_rdy ^ 1'h1;
  assign T26 = state == 3'h2;
  assign T27 = T28 & io_meta_read_ready;
  assign T28 = state == 3'h1;
  assign T29 = T30 & io_req_valid;
  assign T30 = state == 3'h0;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign reply_voluntary = 1'h0;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign reply_r_type = T31;
  assign T31 = T43 ? T41 : T32;
  assign T32 = T40 ? T38 : T33;
  assign T33 = T36 ? T34 : 3'h3;
  assign T34 = T35 ? 3'h2 : 3'h5;
  assign T35 = 2'h3 == old_coh_state;
  assign T36 = req_p_type == 2'h2;
  assign T37 = T29 ? io_req_bits_p_type : req_p_type;
  assign T38 = T39 ? 3'h1 : 3'h4;
  assign T39 = 2'h3 == old_coh_state;
  assign T40 = req_p_type == 2'h1;
  assign T41 = T42 ? 3'h0 : 3'h3;
  assign T42 = 2'h3 == old_coh_state;
  assign T43 = req_p_type == 2'h0;
  assign io_wb_req_bits_data = reply_data;
  assign reply_data = 128'h0;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign reply_addr_beat = 2'h0;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign reply_client_xact_id = 1'h0;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign reply_addr_block = req_addr_block;
  assign T44 = T29 ? io_req_bits_addr_block : req_addr_block;
  assign io_wb_req_valid = T45;
  assign T45 = state == 3'h5;
  assign io_meta_write_bits_data_coh_state = T46;
  assign T46 = T47;
  assign T47 = T52 ? 2'h0 : T48;
  assign T48 = T51 ? 2'h1 : T49;
  assign T49 = T50 ? old_coh_state : old_coh_state;
  assign T50 = req_p_type == 2'h2;
  assign T51 = req_p_type == 2'h1;
  assign T52 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T53;
  assign T53 = req_addr_block >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T64;
  assign T64 = req_addr_block[3'h5:1'h0];
  assign io_meta_write_valid = T54;
  assign T54 = state == 3'h7;
  assign io_meta_read_bits_tag = T55;
  assign T55 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = T65;
  assign T65 = req_addr_block[3'h5:1'h0];
  assign io_meta_read_valid = T56;
  assign T56 = state == 3'h1;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_data = reply_data;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_valid = T57;
  assign T57 = T61 & T58;
  assign T58 = T59 ^ 1'h1;
  assign T59 = tag_matches & T60;
  assign T60 = 2'h3 == old_coh_state;
  assign T61 = state == 3'h4;
  assign io_req_ready = T62;
  assign T62 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      way_en <= io_way_en;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T29) begin
      state <= 3'h1;
    end else if(T27) begin
      state <= 3'h2;
    end else if(T26) begin
      state <= 3'h3;
    end else if(T24) begin
      state <= 3'h1;
    end else if(T1) begin
      state <= 3'h4;
    end else if(T23) begin
      state <= T20;
    end else if(T18) begin
      state <= 3'h0;
    end else if(T16) begin
      state <= 3'h6;
    end else if(T14) begin
      state <= 3'h7;
    end else if(T12) begin
      state <= 3'h0;
    end
    if(T1) begin
      old_coh_state <= io_block_state_state;
    end
    if(T29) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(T29) begin
      req_addr_block <= io_req_bits_addr_block;
    end
  end
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[19:0] T0;
  wire T1;
  wire[5:0] T2;
  wire T3;
  wire T4;
  wire T5;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T0;
  assign T0 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T1 = chosen;
  assign io_out_bits_idx = T2;
  assign T2 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T3;
  assign T3 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T4;
  assign T4 = T5 & io_out_ready;
  assign T5 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[1:0] T0;
  wire T1;
  wire[19:0] T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T0;
  assign T0 = T1 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T1 = chosen;
  assign io_out_bits_data_tag = T2;
  assign T2 = T1 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module LockingArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input  io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input [127:0] io_in_1_bits_data,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input  io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input [127:0] io_in_0_bits_data,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T33;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg  locked;
  wire T34;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire[1:0] T14;
  reg [1:0] R15;
  wire[1:0] T35;
  wire[1:0] T16;
  wire[16:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T20;
  wire[127:0] T21;
  wire[1:0] T22;
  wire T23;
  wire[25:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R15 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T33 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T9 & T7;
  assign T7 = io_out_bits_is_builtin_type & T8;
  assign T8 = 3'h3 == io_out_bits_a_type;
  assign T9 = io_out_ready & io_out_valid;
  assign T34 = reset ? 1'h0 : T10;
  assign T10 = T12 ? 1'h0 : T11;
  assign T11 = T4 ? 1'h1 : locked;
  assign T12 = T9 & T13;
  assign T13 = T14 == 2'h0;
  assign T14 = R15 + 2'h1;
  assign T35 = reset ? 2'h0 : T16;
  assign T16 = T6 ? T14 : R15;
  assign io_out_bits_union = T17;
  assign T17 = T18 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T18 = chosen;
  assign io_out_bits_a_type = T19;
  assign T19 = T18 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_is_builtin_type = T20;
  assign T20 = T18 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_data = T21;
  assign T21 = T18 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr_beat = T22;
  assign T22 = T18 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T23;
  assign T23 = T18 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T24;
  assign T24 = T18 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T25;
  assign T25 = T18 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = locked ? T28 : 1'h1;
  assign T28 = lockIdx == 1'h0;
  assign io_in_1_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = locked ? T32 : T31;
  assign T31 = io_in_0_valid ^ 1'h1;
  assign T32 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T12) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R15 <= 2'h0;
    end else if(T6) begin
      R15 <= T14;
    end
  end
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input  io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input [127:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    input  io_in_1_bits_voluntary,
    input  io_in_1_bits_way_en,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input  io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input [127:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_in_0_bits_voluntary,
    input  io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_out_bits_voluntary,
    output io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[127:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[25:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_way_en = T0;
  assign T0 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T1 = chosen;
  assign io_out_bits_voluntary = T2;
  assign T2 = T1 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_r_type = T3;
  assign T3 = T1 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_data = T4;
  assign T4 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr_beat = T5;
  assign T5 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T7;
  assign T7 = T1 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [39:0] io_in_1_bits_addr,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_kill,
    input  io_in_1_bits_phys,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_kill,
    input  io_in_0_bits_phys,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output io_out_bits_kill,
    output io_out_bits_phys,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[4:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire[4:0] T5;
  wire[7:0] T6;
  wire[39:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T0;
  assign T0 = T1 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T1 = chosen;
  assign io_out_bits_phys = T2;
  assign T2 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_kill = T3;
  assign T3 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_bits_typ = T4;
  assign T4 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_cmd = T5;
  assign T5 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T6;
  assign T6 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T7;
  assign T7 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits = T0;
  assign T0 = T1 ? io_in_1_bits : io_in_0_bits;
  assign T1 = chosen;
  assign io_out_valid = T2;
  assign T2 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T3;
  assign T3 = T4 & io_out_ready;
  assign T4 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[62:0] T11;
  reg [62:0] ram [15:0];
  wire[62:0] T12;
  wire[62:0] T13;
  wire[62:0] T14;
  wire[9:0] T15;
  wire[5:0] T16;
  wire[3:0] T17;
  wire[52:0] T18;
  wire[12:0] T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[4:0] T23;
  wire[7:0] T24;
  wire[39:0] T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_phys, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T18 = {io_enq_bits_addr, T19};
  assign T19 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T20;
  assign T20 = T11[3'h5:3'h5];
  assign io_deq_bits_kill = T21;
  assign T21 = T11[3'h6:3'h6];
  assign io_deq_bits_typ = T22;
  assign T22 = T11[4'h9:3'h7];
  assign io_deq_bits_cmd = T23;
  assign T23 = T11[4'he:4'ha];
  assign io_deq_bits_tag = T24;
  assign T24 = T11[5'h16:4'hf];
  assign io_deq_bits_addr = T25;
  assign T25 = T11[6'h3e:5'h17];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output[127:0] io_mem_req_bits_data,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[25:0] io_wb_req_bits_addr_block,
    output io_wb_req_bits_client_xact_id,
    output[1:0] io_wb_req_bits_addr_beat,
    output[127:0] io_wb_req_bits_data,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  req_way_en;
  wire T133;
  wire T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire[127:0] T139;
  wire[1:0] T140;
  wire T141;
  wire[25:0] T142;
  wire[25:0] T143;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[16:0] T189;
  wire[16:0] T221;
  wire[5:0] T190;
  wire[2:0] T191;
  wire[2:0] T222;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[127:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_voluntary = T134;
  assign T134 = 1'h1;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_data = T139;
  assign T139 = 128'h0;
  assign io_wb_req_bits_addr_beat = T140;
  assign T140 = 2'h0;
  assign io_wb_req_bits_client_xact_id = T141;
  assign T141 = 1'h0;
  assign io_wb_req_bits_addr_block = T142;
  assign T142 = T143;
  assign T143 = {req_old_meta_tag, req_idx};
  assign T144 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_union = T189;
  assign T189 = T221;
  assign T221 = {11'h0, T190};
  assign T190 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T191;
  assign T191 = T222;
  assign T222 = {2'h0, T192};
  assign T192 = T194 | T193;
  assign T193 = req_cmd == 5'h6;
  assign T194 = T196 | T195;
  assign T195 = req_cmd == 5'h3;
  assign T196 = T200 | T197;
  assign T197 = T199 | T198;
  assign T198 = req_cmd == 5'h4;
  assign T199 = req_cmd[2'h3:2'h3];
  assign T200 = T202 | T201;
  assign T201 = req_cmd == 5'h7;
  assign T202 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T203;
  assign T203 = 1'h0;
  assign io_mem_req_bits_data = T204;
  assign T204 = 128'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 1'h0;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_11 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output[127:0] io_mem_req_bits_data,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[25:0] io_wb_req_bits_addr_block,
    output io_wb_req_bits_client_xact_id,
    output[1:0] io_wb_req_bits_addr_beat,
    output[127:0] io_wb_req_bits_data,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  req_way_en;
  wire T133;
  wire T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire[127:0] T139;
  wire[1:0] T140;
  wire T141;
  wire[25:0] T142;
  wire[25:0] T143;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[16:0] T189;
  wire[16:0] T221;
  wire[5:0] T190;
  wire[2:0] T191;
  wire[2:0] T222;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[127:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_voluntary = T134;
  assign T134 = 1'h1;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_data = T139;
  assign T139 = 128'h0;
  assign io_wb_req_bits_addr_beat = T140;
  assign T140 = 2'h0;
  assign io_wb_req_bits_client_xact_id = T141;
  assign T141 = 1'h1;
  assign io_wb_req_bits_addr_block = T142;
  assign T142 = T143;
  assign T143 = {req_old_meta_tag, req_idx};
  assign T144 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_union = T189;
  assign T189 = T221;
  assign T221 = {11'h0, T190};
  assign T190 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T191;
  assign T191 = T222;
  assign T222 = {2'h0, T192};
  assign T192 = T194 | T193;
  assign T193 = req_cmd == 5'h6;
  assign T194 = T196 | T195;
  assign T195 = req_cmd == 5'h3;
  assign T196 = T200 | T197;
  assign T197 = T199 | T198;
  assign T198 = req_cmd == 5'h4;
  assign T199 = req_cmd[2'h3:2'h3];
  assign T200 = T202 | T201;
  assign T201 = req_cmd == 5'h7;
  assign T202 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T203;
  assign T203 = 1'h0;
  assign io_mem_req_bits_data = T204;
  assign T204 = 128'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 1'h1;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_11 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output[127:0] io_mem_req_bits_data,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[25:0] io_wb_req_bits_addr_block,
    output io_wb_req_bits_client_xact_id,
    output[1:0] io_wb_req_bits_addr_beat,
    output[127:0] io_wb_req_bits_data,
    output[2:0] io_wb_req_bits_r_type,
    output io_wb_req_bits_voluntary,
    output io_wb_req_bits_way_en,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire T0;
  wire T1;
  wire[4:0] T101;
  wire[4:0] T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[4:0] T105;
  wire[4:0] T106;
  wire[4:0] T107;
  wire[4:0] T108;
  wire[4:0] T109;
  wire[4:0] T110;
  wire[4:0] T111;
  wire[4:0] T112;
  wire[4:0] T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire[4:0] T116;
  wire T117;
  wire[16:0] T2;
  wire[16:0] T3;
  reg [16:0] sdq_val;
  wire[16:0] T118;
  wire[31:0] T119;
  wire[31:0] T4;
  wire[31:0] T120;
  wire[31:0] T5;
  wire[31:0] T121;
  wire[16:0] T6;
  wire[16:0] T7;
  wire[16:0] T122;
  wire sdq_enq;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[16:0] T16;
  wire[16:0] T17;
  wire[16:0] T18;
  wire[16:0] T19;
  wire[16:0] T20;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[16:0] T23;
  wire[16:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[31:0] T52;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T123;
  wire[16:0] T55;
  wire[16:0] T124;
  wire free_sdq;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire[31:0] T64;
  wire[31:0] T125;
  wire T65;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T66;
  wire tag_match;
  wire[27:0] T67;
  wire[27:0] T141;
  wire[19:0] T68;
  wire[19:0] T69;
  wire[19:0] tagList_1;
  wire idxMatch_1;
  wire[19:0] T70;
  wire[19:0] tagList_0;
  wire idxMatch_0;
  wire T71;
  wire sdq_rdy;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire idx_match;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire[63:0] T88;
  reg [63:0] sdq [16:0];
  wire[63:0] T89;
  wire T90;
  wire T91;
  wire[4:0] T92;
  reg [4:0] R93;
  wire[4:0] T94;
  wire[11:0] T95;
  wire[11:0] refillMux_0_addr;
  wire[11:0] refillMux_1_addr;
  wire T96;
  wire T97;
  wire refillMux_0_way_en;
  wire refillMux_1_way_en;
  wire T98;
  wire T99;
  wire pri_rdy;
  wire T100;
  wire sec_rdy;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire meta_write_arb_io_out_bits_way_en;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr_block;
  wire mem_req_arb_io_out_bits_client_xact_id;
  wire[1:0] mem_req_arb_io_out_bits_addr_beat;
  wire[127:0] mem_req_arb_io_out_bits_data;
  wire mem_req_arb_io_out_bits_is_builtin_type;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[16:0] mem_req_arb_io_out_bits_union;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[25:0] wb_req_arb_io_out_bits_addr_block;
  wire wb_req_arb_io_out_bits_client_xact_id;
  wire[1:0] wb_req_arb_io_out_bits_addr_beat;
  wire[127:0] wb_req_arb_io_out_bits_data;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire wb_req_arb_io_out_bits_voluntary;
  wire wb_req_arb_io_out_bits_way_en;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire[39:0] replay_arb_io_out_bits_addr;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_bits_phys;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire MSHR_io_req_pri_rdy;
  wire MSHR_io_req_sec_rdy;
  wire MSHR_io_idx_match;
  wire[19:0] MSHR_io_tag;
  wire MSHR_io_mem_req_valid;
  wire[25:0] MSHR_io_mem_req_bits_addr_block;
  wire MSHR_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_io_mem_req_bits_addr_beat;
  wire[127:0] MSHR_io_mem_req_bits_data;
  wire MSHR_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_io_mem_req_bits_a_type;
  wire[16:0] MSHR_io_mem_req_bits_union;
  wire MSHR_io_refill_way_en;
  wire[11:0] MSHR_io_refill_addr;
  wire MSHR_io_meta_read_valid;
  wire[5:0] MSHR_io_meta_read_bits_idx;
  wire[19:0] MSHR_io_meta_read_bits_tag;
  wire MSHR_io_meta_write_valid;
  wire[5:0] MSHR_io_meta_write_bits_idx;
  wire MSHR_io_meta_write_bits_way_en;
  wire[19:0] MSHR_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_io_meta_write_bits_data_coh_state;
  wire MSHR_io_replay_valid;
  wire[39:0] MSHR_io_replay_bits_addr;
  wire[7:0] MSHR_io_replay_bits_tag;
  wire[4:0] MSHR_io_replay_bits_cmd;
  wire[2:0] MSHR_io_replay_bits_typ;
  wire MSHR_io_replay_bits_kill;
  wire MSHR_io_replay_bits_phys;
  wire[4:0] MSHR_io_replay_bits_sdq_id;
  wire MSHR_io_wb_req_valid;
  wire[25:0] MSHR_io_wb_req_bits_addr_block;
  wire MSHR_io_wb_req_bits_client_xact_id;
  wire[1:0] MSHR_io_wb_req_bits_addr_beat;
  wire[127:0] MSHR_io_wb_req_bits_data;
  wire[2:0] MSHR_io_wb_req_bits_r_type;
  wire MSHR_io_wb_req_bits_voluntary;
  wire MSHR_io_wb_req_bits_way_en;
  wire MSHR_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[19:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr_block;
  wire MSHR_1_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_1_io_mem_req_bits_addr_beat;
  wire[127:0] MSHR_1_io_mem_req_bits_data;
  wire MSHR_1_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[16:0] MSHR_1_io_mem_req_bits_union;
  wire MSHR_1_io_refill_way_en;
  wire[11:0] MSHR_1_io_refill_addr;
  wire MSHR_1_io_meta_read_valid;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire MSHR_1_io_meta_write_bits_way_en;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire[39:0] MSHR_1_io_replay_bits_addr;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_bits_phys;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_wb_req_valid;
  wire[25:0] MSHR_1_io_wb_req_bits_addr_block;
  wire MSHR_1_io_wb_req_bits_client_xact_id;
  wire[1:0] MSHR_1_io_wb_req_bits_addr_beat;
  wire[127:0] MSHR_1_io_wb_req_bits_data;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire MSHR_1_io_wb_req_bits_voluntary;
  wire MSHR_1_io_wb_req_bits_way_en;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R93 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_grant_valid & T1;
  assign T1 = io_mem_grant_bits_client_xact_id == 1'h1;
  assign T101 = T140 ? 1'h0 : T102;
  assign T102 = T139 ? 1'h1 : T103;
  assign T103 = T138 ? 2'h2 : T104;
  assign T104 = T137 ? 2'h3 : T105;
  assign T105 = T136 ? 3'h4 : T106;
  assign T106 = T135 ? 3'h5 : T107;
  assign T107 = T134 ? 3'h6 : T108;
  assign T108 = T133 ? 3'h7 : T109;
  assign T109 = T132 ? 4'h8 : T110;
  assign T110 = T131 ? 4'h9 : T111;
  assign T111 = T130 ? 4'ha : T112;
  assign T112 = T129 ? 4'hb : T113;
  assign T113 = T128 ? 4'hc : T114;
  assign T114 = T127 ? 4'hd : T115;
  assign T115 = T126 ? 4'he : T116;
  assign T116 = T117 ? 4'hf : 5'h10;
  assign T117 = T2[4'hf:4'hf];
  assign T2 = ~ T3;
  assign T3 = sdq_val[5'h10:1'h0];
  assign T118 = T119[5'h10:1'h0];
  assign T119 = reset ? 32'h0 : T4;
  assign T4 = T65 ? T5 : T120;
  assign T120 = {15'h0, sdq_val};
  assign T5 = T52 | T121;
  assign T121 = {15'h0, T6};
  assign T6 = T16 & T7;
  assign T7 = 17'h0 - T122;
  assign T122 = {16'h0, sdq_enq};
  assign sdq_enq = T15 & T8;
  assign T8 = T12 | T9;
  assign T9 = T11 | T10;
  assign T10 = io_req_bits_cmd == 5'h4;
  assign T11 = io_req_bits_cmd[2'h3:2'h3];
  assign T12 = T14 | T13;
  assign T13 = io_req_bits_cmd == 5'h7;
  assign T14 = io_req_bits_cmd == 5'h1;
  assign T15 = io_req_valid & io_req_ready;
  assign T16 = T51 ? 17'h1 : T17;
  assign T17 = T50 ? 17'h2 : T18;
  assign T18 = T49 ? 17'h4 : T19;
  assign T19 = T48 ? 17'h8 : T20;
  assign T20 = T47 ? 17'h10 : T21;
  assign T21 = T46 ? 17'h20 : T22;
  assign T22 = T45 ? 17'h40 : T23;
  assign T23 = T44 ? 17'h80 : T24;
  assign T24 = T43 ? 17'h100 : T25;
  assign T25 = T42 ? 17'h200 : T26;
  assign T26 = T41 ? 17'h400 : T27;
  assign T27 = T40 ? 17'h800 : T28;
  assign T28 = T39 ? 17'h1000 : T29;
  assign T29 = T38 ? 17'h2000 : T30;
  assign T30 = T37 ? 17'h4000 : T31;
  assign T31 = T36 ? 17'h8000 : T32;
  assign T32 = T33 ? 17'h10000 : 17'h0;
  assign T33 = T34[5'h10:5'h10];
  assign T34 = ~ T35;
  assign T35 = sdq_val[5'h10:1'h0];
  assign T36 = T34[4'hf:4'hf];
  assign T37 = T34[4'he:4'he];
  assign T38 = T34[4'hd:4'hd];
  assign T39 = T34[4'hc:4'hc];
  assign T40 = T34[4'hb:4'hb];
  assign T41 = T34[4'ha:4'ha];
  assign T42 = T34[4'h9:4'h9];
  assign T43 = T34[4'h8:4'h8];
  assign T44 = T34[3'h7:3'h7];
  assign T45 = T34[3'h6:3'h6];
  assign T46 = T34[3'h5:3'h5];
  assign T47 = T34[3'h4:3'h4];
  assign T48 = T34[2'h3:2'h3];
  assign T49 = T34[2'h2:2'h2];
  assign T50 = T34[1'h1:1'h1];
  assign T51 = T34[1'h0:1'h0];
  assign T52 = T125 & T53;
  assign T53 = ~ T54;
  assign T54 = T64 & T123;
  assign T123 = {15'h0, T55};
  assign T55 = 17'h0 - T124;
  assign T124 = {16'h0, free_sdq};
  assign free_sdq = T63 & T56;
  assign T56 = T60 | T57;
  assign T57 = T59 | T58;
  assign T58 = io_replay_bits_cmd == 5'h4;
  assign T59 = io_replay_bits_cmd[2'h3:2'h3];
  assign T60 = T62 | T61;
  assign T61 = io_replay_bits_cmd == 5'h7;
  assign T62 = io_replay_bits_cmd == 5'h1;
  assign T63 = io_replay_ready & io_replay_valid;
  assign T64 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T125 = {15'h0, sdq_val};
  assign T65 = io_replay_valid | sdq_enq;
  assign T126 = T2[4'he:4'he];
  assign T127 = T2[4'hd:4'hd];
  assign T128 = T2[4'hc:4'hc];
  assign T129 = T2[4'hb:4'hb];
  assign T130 = T2[4'ha:4'ha];
  assign T131 = T2[4'h9:4'h9];
  assign T132 = T2[4'h8:4'h8];
  assign T133 = T2[3'h7:3'h7];
  assign T134 = T2[3'h6:3'h6];
  assign T135 = T2[3'h5:3'h5];
  assign T136 = T2[3'h4:3'h4];
  assign T137 = T2[2'h3:2'h3];
  assign T138 = T2[2'h2:2'h2];
  assign T139 = T2[1'h1:1'h1];
  assign T140 = T2[1'h0:1'h0];
  assign T66 = T71 & tag_match;
  assign tag_match = T141 == T67;
  assign T67 = io_req_bits_addr >> 4'hc;
  assign T141 = {8'h0, T68};
  assign T68 = T70 | T69;
  assign T69 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T70 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_io_tag;
  assign idxMatch_0 = MSHR_io_idx_match;
  assign T71 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T72 ^ 1'h1;
  assign T72 = sdq_val == 17'h1ffff;
  assign T73 = io_mem_grant_valid & T74;
  assign T74 = io_mem_grant_bits_client_xact_id == 1'h0;
  assign T75 = T76 & tag_match;
  assign T76 = io_req_valid & sdq_rdy;
  assign T77 = T79 & T78;
  assign T78 = idx_match ^ 1'h1;
  assign idx_match = MSHR_io_idx_match | MSHR_1_io_idx_match;
  assign T79 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T80;
  assign T80 = T83 ? 1'h0 : T81;
  assign T81 = T82 == 1'h0;
  assign T82 = MSHR_io_req_pri_rdy ^ 1'h1;
  assign T83 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T84;
  assign T84 = T87 ? 1'h0 : T85;
  assign T85 = T86 == 1'h0;
  assign T86 = MSHR_io_probe_rdy ^ 1'h1;
  assign T87 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_replay_bits_data = T88;
  assign T88 = sdq[R93];
  assign T90 = sdq_enq & T91;
  assign T91 = T92 < 5'h11;
  assign T92 = T101[3'h4:1'h0];
  assign T94 = free_sdq ? replay_arb_io_out_bits_sdq_id : R93;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_refill_addr = T95;
  assign T95 = T96 ? refillMux_1_addr : refillMux_0_addr;
  assign refillMux_0_addr = MSHR_io_refill_addr;
  assign refillMux_1_addr = MSHR_1_io_refill_addr;
  assign T96 = io_mem_grant_bits_client_xact_id;
  assign io_refill_way_en = T97;
  assign T97 = T96 ? refillMux_1_way_en : refillMux_0_way_en;
  assign refillMux_0_way_en = MSHR_io_refill_way_en;
  assign refillMux_1_way_en = MSHR_1_io_refill_way_en;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T98;
  assign T98 = T99 & sdq_rdy;
  assign T99 = idx_match ? T100 : pri_rdy;
  assign pri_rdy = MSHR_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T100 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_5 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  LockingArbiter_1 mem_req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_1_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_mem_req_valid ),
       .io_in_0_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_in_0_bits_data( MSHR_io_mem_req_bits_data ),
       .io_in_0_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_in_0_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_in_0_bits_union( MSHR_io_mem_req_bits_union ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr_block( mem_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( mem_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_is_builtin_type( mem_req_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_union( mem_req_arb_io_out_bits_union )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_1_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_wb_req_valid ),
       .io_in_0_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_data( MSHR_io_wb_req_bits_data ),
       .io_in_0_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_in_0_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_in_0_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_addr_block( wb_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( wb_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_data( wb_req_arb_io_out_bits_data ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type ),
       .io_out_bits_voluntary( wb_req_arb_io_out_bits_voluntary ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en )
       //.io_chosen(  )
  );
  Arbiter_6 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_replay_valid ),
       .io_in_0_bits_addr( MSHR_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_in_0_bits_typ( MSHR_io_replay_bits_typ ),
       .io_in_0_bits_kill( MSHR_io_replay_bits_kill ),
       .io_in_0_bits_phys( MSHR_io_replay_bits_phys ),
       .io_in_0_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_7 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T77 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  MSHR_0 MSHR(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_io_req_pri_rdy ),
       .io_req_sec_val( T75 ),
       .io_req_sec_rdy( MSHR_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T101 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_io_idx_match ),
       .io_tag( MSHR_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_data( MSHR_io_mem_req_bits_data ),
       .io_mem_req_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_io_mem_req_bits_union ),
       .io_refill_way_en( MSHR_io_refill_way_en ),
       .io_refill_addr( MSHR_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_io_replay_valid ),
       .io_replay_bits_addr( MSHR_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T73 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_io_wb_req_valid ),
       .io_wb_req_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_data( MSHR_io_wb_req_bits_data ),
       .io_wb_req_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_io_probe_rdy )
  );
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T66 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T101 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_mem_req_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_refill_way_en( MSHR_1_io_refill_way_en ),
       .io_refill_addr( MSHR_1_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T0 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );

  always @(posedge clk) begin
    sdq_val <= T118;
    if (T90)
      sdq[T101] <= io_req_bits_data;
    if(free_sdq) begin
      R93 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input  io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[21:0] tags;
  wire[21:0] T2;
  wire[21:0] T3;
  wire[21:0] T4;
  wire[21:0] T22;
  wire T5;
  wire wmask;
  wire T6;
  wire T7;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T23;
  wire[6:0] T8;
  wire[6:0] T9;
  wire[21:0] wdata;
  wire[21:0] T10;
  wire[1:0] T11;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T12;
  wire[19:0] T13;
  wire[19:0] rstVal_tag;
  wire T14;
  wire[5:0] T24;
  wire[6:0] waddr;
  wire[6:0] T25;
  reg [5:0] R15;
  wire[5:0] T16;
  wire[19:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R15 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = tags[1'h1:1'h0];
  MetadataArray_T1 T1 (
    .CLK(clk),
    .W0A(T24),
    .W0E(T14),
    .W0I(wdata),
    .W0M(T3),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(tags)
  );
  assign T3 = T4;
  assign T4 = 22'h0 - T22;
  assign T22 = {21'h0, T5};
  assign T5 = wmask;
  assign wmask = T6;
  assign T6 = rst ? 1'h1 : T7;
  assign T7 = io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T23 = reset ? 7'h0 : T8;
  assign T8 = rst ? T9 : rst_cnt;
  assign T9 = rst_cnt + 7'h1;
  assign wdata = T10;
  assign T10 = {T13, T11};
  assign T11 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T12;
  assign T12 = 2'h0;
  assign T13 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T14 = rst | io_write_valid;
  assign T24 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T25;
  assign T25 = {1'h0, io_write_bits_idx};
  assign T16 = io_read_valid ? io_read_bits_idx : R15;
  assign io_resp_0_tag = T17;
  assign T17 = tags[5'h15:2'h2];
  assign io_write_ready = T18;
  assign T18 = rst ^ 1'h1;
  assign io_read_ready = T19;
  assign T19 = T21 & T20;
  assign T20 = io_write_valid ^ 1'h1;
  assign T21 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T9;
    end
    if(io_read_valid) begin
      R15 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire[5:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[5:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T3;
  assign T3 = T11 ? io_in_4_bits_idx : T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = chosen;
  assign T8 = T9 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign T11 = T7[2'h2:2'h2];
  assign io_out_valid = T12;
  assign T12 = T19 ? io_in_4_valid : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? io_in_1_valid : io_in_0_valid;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T17 ? io_in_3_valid : io_in_2_valid;
  assign T17 = T7[1'h0:1'h0];
  assign T18 = T7[1'h1:1'h1];
  assign T19 = T7[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = T28 | io_in_2_valid;
  assign T28 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_3_valid;
  assign T32 = T33 | io_in_2_valid;
  assign T33 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input  io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire T12;
  wire[7:0] raddr;
  wire[127:0] T2;
  wire[127:0] T3;
  wire[127:0] T4;
  wire[63:0] T5;
  wire[63:0] T13;
  wire T6;
  wire[63:0] T7;
  wire[63:0] T14;
  wire T8;
  wire T9;
  wire[7:0] waddr;
  reg [7:0] R10;
  wire[7:0] T11;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R10 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0 = T0;
  assign T12 = io_read_bits_way_en & io_read_valid;
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T1 T1 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T9),
    .W0I(io_write_bits_data),
    .W0M(T3),
    .R1A(raddr),
    .R1E(T12),
    .R1O(T0)
  );
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = 64'h0 - T13;
  assign T13 = {63'h0, T6};
  assign T6 = io_write_bits_wmask[1'h0:1'h0];
  assign T7 = 64'h0 - T14;
  assign T14 = {63'h0, T8};
  assign T8 = io_write_bits_wmask[1'h1:1'h1];
  assign T9 = io_write_bits_way_en & io_write_valid;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T11 = T12 ? raddr : R10;
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T12) begin
      R10 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[11:0] T2;
  wire[11:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[11:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 2'h0 : T0;
  assign T0 = io_in_1_valid ? 2'h1 : T1;
  assign T1 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = chosen;
  assign T6 = T7 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T7 = T5[1'h0:1'h0];
  assign T8 = T5[1'h1:1'h1];
  assign io_out_bits_way_en = T9;
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T11 = T5[1'h0:1'h0];
  assign T12 = T13 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T13 = T5[1'h0:1'h0];
  assign T14 = T5[1'h1:1'h1];
  assign io_out_valid = T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T5[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T5[1'h0:1'h0];
  assign T20 = T5[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_2_valid;
  assign T29 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[127:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[11:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_wmask = T2;
  assign T2 = T1 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T3;
  assign T3 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T4;
  assign T4 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [4:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T118;
  wire[87:0] T0;
  wire[87:0] T1;
  wire[87:0] T119;
  wire[87:0] T2;
  wire[87:0] wmask;
  wire[87:0] T3;
  wire[47:0] T4;
  wire[23:0] T5;
  wire[15:0] T6;
  wire[7:0] T7;
  wire[7:0] T120;
  wire T8;
  wire[10:0] T9;
  wire[10:0] T10;
  wire[10:0] T11;
  wire[10:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[10:0] T121;
  wire[8:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire[10:0] T122;
  wire[7:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[7:0] T123;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T124;
  wire T32;
  wire[23:0] T33;
  wire[15:0] T34;
  wire[7:0] T35;
  wire[7:0] T125;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T126;
  wire T38;
  wire[7:0] T39;
  wire[7:0] T127;
  wire T40;
  wire[39:0] T41;
  wire[23:0] T42;
  wire[15:0] T43;
  wire[7:0] T44;
  wire[7:0] T128;
  wire T45;
  wire[7:0] T46;
  wire[7:0] T129;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T130;
  wire T49;
  wire[15:0] T50;
  wire[7:0] T51;
  wire[7:0] T131;
  wire T52;
  wire[7:0] T53;
  wire[7:0] T132;
  wire T54;
  wire[87:0] T55;
  wire[87:0] T133;
  wire[63:0] out;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] rhs;
  wire[63:0] T62;
  wire[31:0] T63_1;
  wire[63:0] T64;
  wire[31:0] T65_1_1;
  wire[15:0] T66_1;
  wire[63:0] T67;
  wire[31:0] T68_1_1;
  wire[15:0] T69_1_1;
  wire[7:0] T70_1;
  wire T71;
  wire max;
  wire T72;
  wire T73;
  wire min;
  wire T74;
  wire T75;
  wire less;
  wire T76;
  wire cmp_rhs;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire word;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire cmp_lhs;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire sgned;
  wire T93;
  wire T94;
  wire lt;
  wire T95;
  wire T96;
  wire lt_lo;
  wire[31:0] T97;
  wire[31:0] T98;
  wire eq_hi;
  wire[31:0] T99;
  wire[31:0] T100;
  wire lt_hi;
  wire[31:0] T101;
  wire[31:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire[63:0] T106;
  wire T107;
  wire[63:0] T108;
  wire T109;
  wire[63:0] T110;
  wire T111;
  wire[63:0] adder_out;
  wire[63:0] T112;
  wire[63:0] mask;
  wire[63:0] T134;
  wire[31:0] T113;
  wire T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire T117;


  assign io_out = T118;
  assign T118 = T0[6'h3f:1'h0];
  assign T0 = T55 | T1;
  assign T1 = T2 & T119;
  assign T119 = {24'h0, io_lhs};
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T41, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = {T29, T7};
  assign T7 = 8'h0 - T120;
  assign T120 = {7'h0, T8};
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T26 ? T122 : T10;
  assign T10 = T21 ? T121 : T11;
  assign T11 = T15 ? T12 : 11'hff;
  assign T12 = 4'hf << T13;
  assign T13 = {T14, 2'h0};
  assign T14 = io_addr[2'h2:2'h2];
  assign T15 = T17 | T16;
  assign T16 = io_typ == 3'h6;
  assign T17 = io_typ == 3'h2;
  assign T121 = {2'h0, T18};
  assign T18 = 2'h3 << T19;
  assign T19 = {T20, 1'h0};
  assign T20 = io_addr[2'h2:1'h1];
  assign T21 = T23 | T22;
  assign T22 = io_typ == 3'h5;
  assign T23 = io_typ == 3'h1;
  assign T122 = {3'h0, T24};
  assign T24 = 1'h1 << T25;
  assign T25 = io_addr[2'h2:1'h0];
  assign T26 = T28 | T27;
  assign T27 = io_typ == 3'h4;
  assign T28 = io_typ == 3'h0;
  assign T29 = 8'h0 - T123;
  assign T123 = {7'h0, T30};
  assign T30 = T9[1'h1:1'h1];
  assign T31 = 8'h0 - T124;
  assign T124 = {7'h0, T32};
  assign T32 = T9[2'h2:2'h2];
  assign T33 = {T39, T34};
  assign T34 = {T37, T35};
  assign T35 = 8'h0 - T125;
  assign T125 = {7'h0, T36};
  assign T36 = T9[2'h3:2'h3];
  assign T37 = 8'h0 - T126;
  assign T126 = {7'h0, T38};
  assign T38 = T9[3'h4:3'h4];
  assign T39 = 8'h0 - T127;
  assign T127 = {7'h0, T40};
  assign T40 = T9[3'h5:3'h5];
  assign T41 = {T50, T42};
  assign T42 = {T48, T43};
  assign T43 = {T46, T44};
  assign T44 = 8'h0 - T128;
  assign T128 = {7'h0, T45};
  assign T45 = T9[3'h6:3'h6];
  assign T46 = 8'h0 - T129;
  assign T129 = {7'h0, T47};
  assign T47 = T9[3'h7:3'h7];
  assign T48 = 8'h0 - T130;
  assign T130 = {7'h0, T49};
  assign T49 = T9[4'h8:4'h8];
  assign T50 = {T53, T51};
  assign T51 = 8'h0 - T131;
  assign T131 = {7'h0, T52};
  assign T52 = T9[4'h9:4'h9];
  assign T53 = 8'h0 - T132;
  assign T132 = {7'h0, T54};
  assign T54 = T9[4'ha:4'ha];
  assign T55 = wmask & T133;
  assign T133 = {24'h0, out};
  assign out = T117 ? adder_out : T56;
  assign T56 = T111 ? T110 : T57;
  assign T57 = T109 ? T108 : T58;
  assign T58 = T107 ? T106 : T59;
  assign T59 = T71 ? io_lhs : T60;
  assign T60 = T26 ? T67 : T61;
  assign T61 = T21 ? T64 : rhs;
  assign rhs = T15 ? T62 : io_rhs;
  assign T62 = {T63_1, T63_1};
  assign T63_1 = io_rhs[5'h1f:1'h0];
  assign T64 = {T65_1_1, T65_1_1};
  assign T65_1_1 = {T66_1, T66_1};
  assign T66_1 = io_rhs[4'hf:1'h0];
  assign T67 = {T68_1_1, T68_1_1};
  assign T68_1_1 = {T69_1_1, T69_1_1};
  assign T69_1_1 = {T70_1, T70_1};
  assign T70_1 = io_rhs[3'h7:1'h0];
  assign T71 = less ? min : max;
  assign max = T73 | T72;
  assign T72 = io_cmd == 5'hf;
  assign T73 = io_cmd == 5'hd;
  assign min = T75 | T74;
  assign T74 = io_cmd == 5'he;
  assign T75 = io_cmd == 5'hc;
  assign less = T105 ? lt : T76;
  assign T76 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T79 ? T78 : T77;
  assign T77 = rhs[6'h3f:6'h3f];
  assign T78 = rhs[5'h1f:5'h1f];
  assign T79 = word & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_addr[2'h2:2'h2];
  assign word = T83 | T82;
  assign T82 = io_typ == 3'h4;
  assign T83 = T85 | T84;
  assign T84 = io_typ == 3'h0;
  assign T85 = T87 | T86;
  assign T86 = io_typ == 3'h6;
  assign T87 = io_typ == 3'h2;
  assign cmp_lhs = T90 ? T89 : T88;
  assign T88 = io_lhs[6'h3f:6'h3f];
  assign T89 = io_lhs[5'h1f:5'h1f];
  assign T90 = word & T91;
  assign T91 = T92 ^ 1'h1;
  assign T92 = io_addr[2'h2:2'h2];
  assign sgned = T94 | T93;
  assign T93 = io_cmd == 5'hd;
  assign T94 = io_cmd == 5'hc;
  assign lt = word ? T103 : T95;
  assign T95 = lt_hi | T96;
  assign T96 = eq_hi & lt_lo;
  assign lt_lo = T98 < T97;
  assign T97 = rhs[5'h1f:1'h0];
  assign T98 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T100 == T99;
  assign T99 = rhs[6'h3f:6'h20];
  assign T100 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T102 < T101;
  assign T101 = rhs[6'h3f:6'h20];
  assign T102 = io_lhs[6'h3f:6'h20];
  assign T103 = T104 ? lt_hi : lt_lo;
  assign T104 = io_addr[2'h2:2'h2];
  assign T105 = cmp_lhs == cmp_rhs;
  assign T106 = io_lhs ^ rhs;
  assign T107 = io_cmd == 5'h9;
  assign T108 = io_lhs | rhs;
  assign T109 = io_cmd == 5'ha;
  assign T110 = io_lhs & rhs;
  assign T111 = io_cmd == 5'hb;
  assign adder_out = T115 + T112;
  assign T112 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T134;
  assign T134 = {32'h0, T113};
  assign T113 = T114 << 5'h1f;
  assign T114 = io_addr[2'h2:2'h2];
  assign T115 = T116;
  assign T116 = io_lhs & mask;
  assign T117 = io_cmd == 5'h8;
endmodule

module LockingArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input  io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input [127:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    input  io_in_1_bits_voluntary,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input  io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input [127:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_in_0_bits_voluntary,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output[127:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_out_bits_voluntary,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T35;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T36;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T37;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[127:0] T23;
  wire[1:0] T24;
  wire T25;
  wire[25:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T35 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T12 & T7;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_out_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_out_bits_r_type;
  assign T11 = 3'h0 == io_out_bits_r_type;
  assign T12 = io_out_ready & io_out_valid;
  assign T36 = reset ? 1'h0 : T13;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = T4 ? 1'h1 : locked;
  assign T15 = T12 & T16;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T37 = reset ? 2'h0 : T19;
  assign T19 = T6 ? T17 : R18;
  assign io_out_bits_voluntary = T20;
  assign T20 = T21 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign T21 = chosen;
  assign io_out_bits_r_type = T22;
  assign T22 = T21 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_data = T23;
  assign T23 = T21 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr_beat = T24;
  assign T24 = T21 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T25;
  assign T25 = T21 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T26;
  assign T26 = T21 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T27;
  assign T27 = T21 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = locked ? T30 : 1'h1;
  assign T30 = lockIdx == 1'h0;
  assign io_in_1_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T34 : T33;
  assign T33 = io_in_0_valid ^ 1'h1;
  assign T34 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T6) begin
      R18 <= T17;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_addr,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_kill,
    input  io_cpu_req_bits_phys,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_addr,
    output[7:0] io_cpu_resp_bits_tag,
    output[4:0] io_cpu_resp_bits_cmd,
    output[2:0] io_cpu_resp_bits_typ,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_invalidate_lr,
    output io_cpu_ordered,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [127:0] io_mem_grant_bits_data,
    input  io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [25:0] io_mem_probe_bits_addr_block,
    input [1:0] io_mem_probe_bits_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[25:0] io_mem_release_bits_addr_block,
    output io_mem_release_bits_client_xact_id,
    output[1:0] io_mem_release_bits_addr_beat,
    output[127:0] io_mem_release_bits_data,
    output[2:0] io_mem_release_bits_r_type,
    output io_mem_release_bits_voluntary
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg  R4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg [63:0] s2_req_data;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  s1_replay;
  wire T412;
  wire T20;
  wire T21;
  wire s1_write;
  wire T22;
  wire T23;
  reg [4:0] s1_req_cmd;
  wire[4:0] T24;
  wire[4:0] T25;
  wire[4:0] T26;
  reg [4:0] s2_req_cmd;
  wire[4:0] T27;
  wire s2_recycle;
  wire T28;
  reg  s2_recycle_next;
  wire T413;
  wire T29;
  wire T30;
  reg  s1_valid;
  wire T414;
  wire T31;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire s2_word_idx_1;
  reg [39:0] s2_req_addr;
  wire[39:0] T36;
  wire[39:0] T415;
  wire[31:0] s1_addr;
  wire[11:0] T37;
  reg [39:0] s1_req_addr;
  wire[39:0] T38;
  wire[39:0] T39;
  wire[39:0] T40;
  wire[39:0] T41;
  wire[39:0] T42;
  wire[39:0] T416;
  wire[31:0] T43;
  wire[25:0] T44;
  wire[39:0] T417;
  wire[31:0] T45;
  wire[25:0] T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire s2_hit;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  reg [1:0] s2_hit_state_state;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire s2_tag_match;
  reg  s2_tag_match_way;
  wire T82;
  wire s1_tag_match_way;
  wire T83;
  wire T84;
  wire T85;
  wire s1_tag_eq_way;
  wire T86;
  wire[19:0] T87;
  wire T88;
  wire s2_replay;
  wire T89;
  reg  R90;
  wire T418;
  reg  s2_valid;
  wire T419;
  wire s1_valid_masked;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[63:0] T98;
  wire T99;
  reg  s1_recycled;
  wire T420;
  wire T100;
  wire[63:0] T421;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[6:0] T101;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T102;
  wire[63:0] T103;
  wire[127:0] s2_data_0;
  wire[127:0] T104;
  wire[127:0] T105;
  reg [63:0] R106;
  wire[63:0] T422;
  wire[127:0] T107;
  wire[127:0] T423;
  wire[127:0] T108;
  wire T109;
  wire T110;
  reg [63:0] R111;
  wire[63:0] T112;
  wire[63:0] T113;
  wire[63:0] T114;
  wire[127:0] T424;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T115;
  wire[63:0] T116;
  wire[63:0] T117;
  reg [63:0] s4_req_data;
  wire[63:0] T118;
  wire T119;
  reg  s3_valid;
  wire T425;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire s2_sc_fail;
  wire T130;
  wire s2_lrsc_addr_match;
  wire T131;
  wire[33:0] T132;
  reg [33:0] lrsc_addr;
  wire[33:0] T133;
  wire[33:0] T134;
  wire T135;
  wire s2_lr;
  wire T136;
  wire T137;
  wire s2_valid_masked;
  wire T138;
  wire T139;
  wire s2_nack;
  wire s2_nack_miss;
  wire T140;
  wire T141;
  wire T142;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T143;
  wire s1_nack;
  wire T144;
  wire T145;
  wire T146;
  wire[5:0] T147;
  wire T148;
  wire T149;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T426;
  wire[4:0] T150;
  wire[4:0] T151;
  wire[4:0] T152;
  wire[4:0] T153;
  wire[4:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire s2_sc;
  wire T158;
  wire T159;
  reg [63:0] s3_req_data;
  wire[63:0] T427;
  wire[127:0] T160;
  wire[127:0] T428;
  wire[63:0] T161;
  wire[127:0] T162;
  wire[127:0] T429;
  wire[127:0] s2_data_corrected;
  wire[127:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  reg [4:0] s3_req_cmd;
  wire[4:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[36:0] T185;
  reg [39:0] s3_req_addr;
  wire[39:0] T186;
  wire[36:0] T430;
  wire[28:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[36:0] T198;
  wire[36:0] T431;
  wire[28:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg [4:0] s4_req_cmd;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[36:0] T216;
  reg [39:0] s4_req_addr;
  wire[39:0] T217;
  wire[36:0] T432;
  wire[28:0] T218;
  reg  s4_valid;
  wire T433;
  wire T219;
  reg  s2_store_bypass;
  wire T220;
  wire T221;
  reg [2:0] s2_req_typ;
  wire[2:0] T222;
  reg [2:0] s1_req_typ;
  wire[2:0] T223;
  wire[2:0] T224;
  wire[2:0] T225;
  wire[5:0] T434;
  wire[127:0] T226;
  wire[1:0] rowWMask;
  wire rowIdx;
  wire T227;
  wire[11:0] T435;
  reg  s3_way;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire[11:0] T436;
  wire[11:0] T437;
  wire[11:0] T438;
  wire[127:0] T239;
  wire[127:0] T240;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[5:0] T439;
  wire[33:0] T241;
  wire[5:0] T440;
  wire[33:0] T242;
  reg  s1_req_phys;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  reg  s2_req_phys;
  wire T248;
  wire[27:0] T249;
  wire T250;
  wire T251;
  wire T252;
  wire s1_readwrite;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire s1_read;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T441;
  wire[1:0] T264;
  wire[1:0] s2_replaced_way_en;
  reg  R265;
  wire T266;
  wire[1:0] T442;
  wire[1:0] T267;
  reg [1:0] s2_repl_meta_coh_state;
  wire[1:0] T268;
  wire[1:0] T269;
  wire[19:0] T270;
  reg [19:0] s2_repl_meta_tag;
  wire[19:0] T271;
  wire[19:0] T272;
  reg  s2_req_kill;
  wire T273;
  reg  s1_req_kill;
  wire T274;
  wire T275;
  wire T276;
  reg [7:0] s2_req_tag;
  wire[7:0] T277;
  reg [7:0] s1_req_tag;
  wire[7:0] T278;
  wire[7:0] T279;
  wire[7:0] T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire misaligned;
  wire T319;
  wire T320;
  wire[2:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire[1:0] T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire s1_sc;
  wire[63:0] T339;
  wire[63:0] T443;
  wire[63:0] T340;
  wire[7:0] T341;
  wire[7:0] T342;
  wire[7:0] T343;
  wire[63:0] T344;
  wire[15:0] T345;
  wire[15:0] T346;
  wire[63:0] T347;
  wire[31:0] T348;
  wire[31:0] T349;
  wire[31:0] T350;
  wire T351;
  wire[31:0] T352;
  wire[31:0] T353;
  wire[31:0] T354;
  wire[31:0] T444;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire[15:0] T367;
  wire T368;
  wire[47:0] T369;
  wire[47:0] T370;
  wire[47:0] T371;
  wire[47:0] T445;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire[7:0] T377;
  wire T378;
  wire[55:0] T379;
  wire[55:0] T380;
  wire[55:0] T381;
  wire[55:0] T446;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  reg  block_miss;
  wire T447;
  wire T410;
  wire T411;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire wb_io_data_req_bits_way_en;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[25:0] wb_io_release_bits_addr_block;
  wire wb_io_release_bits_client_xact_id;
  wire[1:0] wb_io_release_bits_addr_beat;
  wire[127:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_r_type;
  wire wb_io_release_bits_voluntary;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[25:0] prober_io_rep_bits_addr_block;
  wire prober_io_rep_bits_client_xact_id;
  wire[1:0] prober_io_rep_bits_addr_beat;
  wire[127:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_r_type;
  wire prober_io_rep_bits_voluntary;
  wire prober_io_meta_read_valid;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire prober_io_meta_write_bits_way_en;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[25:0] prober_io_wb_req_bits_addr_block;
  wire prober_io_wb_req_bits_client_xact_id;
  wire[1:0] prober_io_wb_req_bits_addr_beat;
  wire[127:0] prober_io_wb_req_bits_data;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire prober_io_wb_req_bits_voluntary;
  wire prober_io_wb_req_bits_way_en;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[19:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire metaWriteArb_io_out_bits_way_en;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire readArb_io_out_bits_way_en;
  wire[11:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire writeArb_io_out_bits_way_en;
  wire[11:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[25:0] releaseArb_io_out_bits_addr_block;
  wire releaseArb_io_out_bits_client_xact_id;
  wire[1:0] releaseArb_io_out_bits_addr_beat;
  wire[127:0] releaseArb_io_out_bits_data;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire releaseArb_io_out_bits_voluntary;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[1:0] FlowThroughSerializer_io_out_bits_addr_beat;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;
  wire FlowThroughSerializer_io_out_bits_client_xact_id;
  wire[2:0] FlowThroughSerializer_io_out_bits_manager_xact_id;
  wire FlowThroughSerializer_io_out_bits_is_builtin_type;
  wire[3:0] FlowThroughSerializer_io_out_bits_g_type;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[25:0] wbArb_io_out_bits_addr_block;
  wire wbArb_io_out_bits_client_xact_id;
  wire[1:0] wbArb_io_out_bits_addr_beat;
  wire[127:0] wbArb_io_out_bits_data;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire wbArb_io_out_bits_voluntary;
  wire wbArb_io_out_bits_way_en;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[19:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[26:0] dtlb_io_ptw_req_bits_addr;
  wire[1:0] dtlb_io_ptw_req_bits_prv;
  wire dtlb_io_ptw_req_bits_store;
  wire dtlb_io_ptw_req_bits_fetch;
  wire mshrs_io_req_ready;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr_block;
  wire mshrs_io_mem_req_bits_client_xact_id;
  wire[1:0] mshrs_io_mem_req_bits_addr_beat;
  wire[127:0] mshrs_io_mem_req_bits_data;
  wire mshrs_io_mem_req_bits_is_builtin_type;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[16:0] mshrs_io_mem_req_bits_union;
  wire mshrs_io_refill_way_en;
  wire[11:0] mshrs_io_refill_addr;
  wire mshrs_io_meta_read_valid;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire mshrs_io_meta_write_bits_way_en;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire[39:0] mshrs_io_replay_bits_addr;
  wire[7:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_kill;
  wire mshrs_io_replay_bits_phys;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_wb_req_valid;
  wire[25:0] mshrs_io_wb_req_bits_addr_block;
  wire mshrs_io_wb_req_bits_client_xact_id;
  wire[1:0] mshrs_io_wb_req_bits_addr_beat;
  wire[127:0] mshrs_io_wb_req_bits_data;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire mshrs_io_wb_req_bits_voluntary;
  wire mshrs_io_wb_req_bits_way_en;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {1{$random}};
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    s2_req_addr = {2{$random}};
    s1_req_addr = {2{$random}};
    s2_hit_state_state = {1{$random}};
    s2_tag_match_way = {1{$random}};
    R90 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R106 = {2{$random}};
    R111 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R265 = {1{$random}};
    s2_repl_meta_coh_state = {1{$random}};
    s2_repl_meta_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    block_miss = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = R4 & io_cpu_resp_valid;
  assign T5 = T6 | io_cpu_xcpt_pf_st;
  assign T6 = T7 | io_cpu_xcpt_pf_ld;
  assign T7 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T8 = writeArb_io_in_1_ready | T9;
  assign T9 = T10 ^ 1'h1;
  assign T10 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T14 : T11;
  assign T11 = T13 | T12;
  assign T12 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T13 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T14 = T16 | T15;
  assign T15 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T16 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T17 = T99 ? s1_req_data : T18;
  assign T18 = T21 ? T19 : s2_req_data;
  assign T19 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T412 = reset ? 1'h0 : T20;
  assign T20 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T21 = s1_clk_en & s1_write;
  assign s1_write = T93 | T22;
  assign T22 = T92 | T23;
  assign T23 = s1_req_cmd == 5'h4;
  assign T24 = s2_recycle ? s2_req_cmd : T25;
  assign T25 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T26;
  assign T26 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T27 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T28;
  assign T28 = s2_recycle_ecc | s2_recycle_next;
  assign T413 = reset ? 1'h0 : T29;
  assign T29 = T30 ? s2_recycle_ecc : s2_recycle_next;
  assign T30 = s1_valid | s1_replay;
  assign T414 = reset ? 1'h0 : T31;
  assign T31 = io_cpu_req_ready & io_cpu_req_valid;
  assign s2_recycle_ecc = T49 & s2_data_correctable;
  assign s2_data_correctable = T47 & T32;
  assign T32 = T33 - 1'h1;
  assign T33 = 1'h1 << T34;
  assign T34 = T35 + 1'h1;
  assign T35 = s2_word_idx_1 - s2_word_idx_1;
  assign s2_word_idx_1 = s2_req_addr[2'h3:2'h3];
  assign T36 = s1_clk_en ? T415 : s2_req_addr;
  assign T415 = {8'h0, s1_addr};
  assign s1_addr = {dtlb_io_resp_ppn, T37};
  assign T37 = s1_req_addr[4'hb:1'h0];
  assign T38 = s2_recycle ? s2_req_addr : T39;
  assign T39 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T40;
  assign T40 = prober_io_meta_read_valid ? T417 : T41;
  assign T41 = wb_io_meta_read_valid ? T416 : T42;
  assign T42 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T416 = {8'h0, T43};
  assign T43 = T44 << 3'h6;
  assign T44 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T417 = {8'h0, T45};
  assign T45 = T46 << 3'h6;
  assign T46 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T47 = T48 >> s2_word_idx_1;
  assign T48 = 2'h0;
  assign T49 = T88 & s2_hit;
  assign s2_hit = T61 & T50;
  assign T50 = s2_hit_state_state == T51;
  assign T51 = T52;
  assign T52 = T53 ? 2'h3 : s2_hit_state_state;
  assign T53 = T57 | T54;
  assign T54 = T56 | T55;
  assign T55 = s2_req_cmd == 5'h4;
  assign T56 = s2_req_cmd[2'h3:2'h3];
  assign T57 = T59 | T58;
  assign T58 = s2_req_cmd == 5'h7;
  assign T59 = s2_req_cmd == 5'h1;
  assign T60 = s1_clk_en ? meta_io_resp_0_coh_state : s2_hit_state_state;
  assign T61 = s2_tag_match & T62;
  assign T62 = T71 ? T68 : T63;
  assign T63 = T65 | T64;
  assign T64 = 2'h3 == s2_hit_state_state;
  assign T65 = T67 | T66;
  assign T66 = 2'h2 == s2_hit_state_state;
  assign T67 = 2'h1 == s2_hit_state_state;
  assign T68 = T70 | T69;
  assign T69 = 2'h3 == s2_hit_state_state;
  assign T70 = 2'h2 == s2_hit_state_state;
  assign T71 = T73 | T72;
  assign T72 = s2_req_cmd == 5'h6;
  assign T73 = T75 | T74;
  assign T74 = s2_req_cmd == 5'h3;
  assign T75 = T79 | T76;
  assign T76 = T78 | T77;
  assign T77 = s2_req_cmd == 5'h4;
  assign T78 = s2_req_cmd[2'h3:2'h3];
  assign T79 = T81 | T80;
  assign T80 = s2_req_cmd == 5'h7;
  assign T81 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 1'h0;
  assign T82 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T83;
  assign T83 = T85 & T84;
  assign T84 = meta_io_resp_0_coh_state != 2'h0;
  assign T85 = s1_tag_eq_way;
  assign s1_tag_eq_way = T86;
  assign T86 = meta_io_resp_0_tag == T87;
  assign T87 = s1_addr >> 4'hc;
  assign T88 = s2_valid | s2_replay;
  assign s2_replay = R90 & T89;
  assign T89 = s2_req_cmd != 5'h5;
  assign T418 = reset ? 1'h0 : s1_replay;
  assign T419 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T91;
  assign T91 = io_cpu_req_bits_kill ^ 1'h1;
  assign T92 = s1_req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = s1_req_cmd == 5'h7;
  assign T95 = s1_req_cmd == 5'h1;
  assign T96 = s2_recycle ? s2_req_data : T97;
  assign T97 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T98;
  assign T98 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T99 = s1_clk_en & s1_recycled;
  assign T420 = reset ? 1'h0 : T100;
  assign T100 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T421 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T424 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> T101;
  assign T101 = {s2_word_idx_1, 6'h0};
  assign s2_data_uncorrected = T102;
  assign T102 = {T114, T103};
  assign T103 = s2_data_0[6'h3f:1'h0];
  assign s2_data_0 = T104;
  assign T104 = T105;
  assign T105 = {R111, R106};
  assign T422 = T107[6'h3f:1'h0];
  assign T107 = T109 ? T108 : T423;
  assign T423 = {64'h0, R106};
  assign T108 = data_io_resp_0 >> 1'h0;
  assign T109 = s1_clk_en & T110;
  assign T110 = s1_tag_eq_way;
  assign T112 = T109 ? T113 : R111;
  assign T113 = data_io_resp_0 >> 7'h40;
  assign T114 = s2_data_0[7'h7f:7'h40];
  assign T424 = {64'h0, s2_store_bypass_data};
  assign T115 = T203 ? T116 : s2_store_bypass_data;
  assign T116 = T188 ? amoalu_io_out : T117;
  assign T117 = T174 ? s3_req_data : s4_req_data;
  assign T118 = T119 ? s3_req_data : s4_req_data;
  assign T119 = s3_valid & metaReadArb_io_out_valid;
  assign T425 = reset ? 1'h0 : T120;
  assign T120 = T128 & T121;
  assign T121 = T125 | T122;
  assign T122 = T124 | T123;
  assign T123 = s2_req_cmd == 5'h4;
  assign T124 = s2_req_cmd[2'h3:2'h3];
  assign T125 = T127 | T126;
  assign T126 = s2_req_cmd == 5'h7;
  assign T127 = s2_req_cmd == 5'h1;
  assign T128 = T158 & T129;
  assign T129 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T130;
  assign T130 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T131;
  assign T131 = lrsc_addr == T132;
  assign T132 = s2_req_addr >> 3'h6;
  assign T133 = T135 ? T134 : lrsc_addr;
  assign T134 = s2_req_addr >> 3'h6;
  assign T135 = T136 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T136 = T137 | s2_replay;
  assign T137 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T138;
  assign T138 = s2_valid & T139;
  assign T139 = s2_nack ^ 1'h1;
  assign s2_nack = T142 | s2_nack_miss;
  assign s2_nack_miss = T141 & T140;
  assign T140 = mshrs_io_req_ready ^ 1'h1;
  assign T141 = s2_hit ^ 1'h1;
  assign T142 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T143 = T149 ? s1_nack : s2_nack_hit;
  assign s1_nack = T148 | T144;
  assign T144 = T146 & T145;
  assign T145 = prober_io_req_ready ^ 1'h1;
  assign T146 = T147 == prober_io_meta_write_bits_idx;
  assign T147 = s1_req_addr[4'hb:3'h6];
  assign T148 = T250 & dtlb_io_resp_miss;
  assign T149 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T426 = reset ? 5'h0 : T150;
  assign T150 = io_cpu_invalidate_lr ? 5'h0 : T151;
  assign T151 = T157 ? 5'h0 : T152;
  assign T152 = T155 ? 5'h1f : T153;
  assign T153 = lrsc_valid ? T154 : lrsc_count;
  assign T154 = lrsc_count - 5'h1;
  assign T155 = T135 & T156;
  assign T156 = lrsc_valid ^ 1'h1;
  assign T157 = T136 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T158 = T159 | s2_replay;
  assign T159 = s2_valid_masked & s2_hit;
  assign T427 = T160[6'h3f:1'h0];
  assign T160 = T164 ? T162 : T428;
  assign T428 = {64'h0, T161};
  assign T161 = T164 ? s2_req_data : s3_req_data;
  assign T162 = s2_data_correctable ? s2_data_corrected : T429;
  assign T429 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T163;
  assign T163 = {T114, T103};
  assign T164 = T173 & T165;
  assign T165 = T166 | s2_data_correctable;
  assign T166 = T170 | T167;
  assign T167 = T169 | T168;
  assign T168 = s2_req_cmd == 5'h4;
  assign T169 = s2_req_cmd[2'h3:2'h3];
  assign T170 = T172 | T171;
  assign T171 = s2_req_cmd == 5'h7;
  assign T172 = s2_req_cmd == 5'h1;
  assign T173 = s2_valid | s2_replay;
  assign T174 = T183 & T175;
  assign T175 = T180 | T176;
  assign T176 = T179 | T177;
  assign T177 = s3_req_cmd == 5'h4;
  assign T178 = T164 ? s2_req_cmd : s3_req_cmd;
  assign T179 = s3_req_cmd[2'h3:2'h3];
  assign T180 = T182 | T181;
  assign T181 = s3_req_cmd == 5'h7;
  assign T182 = s3_req_cmd == 5'h1;
  assign T183 = s3_valid & T184;
  assign T184 = T430 == T185;
  assign T185 = s3_req_addr >> 2'h3;
  assign T186 = T164 ? s2_req_addr : s3_req_addr;
  assign T430 = {8'h0, T187};
  assign T187 = s1_addr >> 2'h3;
  assign T188 = T196 & T189;
  assign T189 = T193 | T190;
  assign T190 = T192 | T191;
  assign T191 = s2_req_cmd == 5'h4;
  assign T192 = s2_req_cmd[2'h3:2'h3];
  assign T193 = T195 | T194;
  assign T194 = s2_req_cmd == 5'h7;
  assign T195 = s2_req_cmd == 5'h1;
  assign T196 = T200 & T197;
  assign T197 = T431 == T198;
  assign T198 = s2_req_addr >> 2'h3;
  assign T431 = {8'h0, T199};
  assign T199 = s1_addr >> 2'h3;
  assign T200 = T202 & T201;
  assign T201 = s2_sc_fail ^ 1'h1;
  assign T202 = s2_valid_masked | s2_replay;
  assign T203 = s1_clk_en & T204;
  assign T204 = T219 | T205;
  assign T205 = T214 & T206;
  assign T206 = T211 | T207;
  assign T207 = T210 | T208;
  assign T208 = s4_req_cmd == 5'h4;
  assign T209 = T119 ? s3_req_cmd : s4_req_cmd;
  assign T210 = s4_req_cmd[2'h3:2'h3];
  assign T211 = T213 | T212;
  assign T212 = s4_req_cmd == 5'h7;
  assign T213 = s4_req_cmd == 5'h1;
  assign T214 = s4_valid & T215;
  assign T215 = T432 == T216;
  assign T216 = s4_req_addr >> 2'h3;
  assign T217 = T119 ? s3_req_addr : s4_req_addr;
  assign T432 = {8'h0, T218};
  assign T218 = s1_addr >> 2'h3;
  assign T433 = reset ? 1'h0 : s3_valid;
  assign T219 = T188 | T174;
  assign T220 = T203 ? 1'h1 : T221;
  assign T221 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T222 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T223 = s2_recycle ? s2_req_typ : T224;
  assign T224 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T225;
  assign T225 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T434 = s2_req_addr[3'h5:1'h0];
  assign T226 = {s3_req_data, s3_req_data};
  assign rowWMask = 1'h1 << rowIdx;
  assign rowIdx = T227;
  assign T227 = s3_req_addr[2'h3:2'h3];
  assign T435 = s3_req_addr[4'hb:1'h0];
  assign T228 = T164 ? s2_tag_match_way : s3_way;
  assign T229 = FlowThroughSerializer_io_out_valid & T230;
  assign T230 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T234 : T231;
  assign T231 = T233 | T232;
  assign T232 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T233 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T234 = T236 | T235;
  assign T235 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T236 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T237 = T238 | T8;
  assign T238 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T436 = s2_req_addr[4'hb:1'h0];
  assign T437 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T438 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T239 = T240;
  assign T240 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T439 = T241[3'h5:1'h0];
  assign T241 = s2_req_addr >> 3'h6;
  assign T440 = T242[3'h5:1'h0];
  assign T242 = io_cpu_req_bits_addr >> 3'h6;
  assign T243 = s2_recycle ? s2_req_phys : T244;
  assign T244 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T245;
  assign T245 = prober_io_meta_read_valid ? 1'h1 : T246;
  assign T246 = wb_io_meta_read_valid ? 1'h1 : T247;
  assign T247 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T248 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T249 = s1_req_addr >> 4'hc;
  assign T250 = T252 & T251;
  assign T251 = s1_req_phys ^ 1'h1;
  assign T252 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T256 | T253;
  assign T253 = T255 | T254;
  assign T254 = s1_req_cmd == 5'h3;
  assign T255 = s1_req_cmd == 5'h2;
  assign T256 = s1_read | s1_write;
  assign s1_read = T260 | T257;
  assign T257 = T259 | T258;
  assign T258 = s1_req_cmd == 5'h4;
  assign T259 = s1_req_cmd[2'h3:2'h3];
  assign T260 = T262 | T261;
  assign T261 = s1_req_cmd == 5'h6;
  assign T262 = s1_req_cmd == 5'h0;
  assign T263 = T8 & FlowThroughSerializer_io_out_valid;
  assign T441 = T264[1'h0:1'h0];
  assign T264 = s2_tag_match ? T442 : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R265;
  assign T266 = s1_clk_en ? 1'h0 : R265;
  assign T442 = {1'h0, s2_tag_match_way};
  assign T267 = s2_tag_match ? T269 : s2_repl_meta_coh_state;
  assign T268 = s1_clk_en ? meta_io_resp_0_coh_state : s2_repl_meta_coh_state;
  assign T269 = s2_hit_state_state;
  assign T270 = s2_tag_match ? T272 : s2_repl_meta_tag;
  assign T271 = s1_clk_en ? meta_io_resp_0_tag : s2_repl_meta_tag;
  assign T272 = s2_repl_meta_tag;
  assign T273 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T274 = s2_recycle ? s2_req_kill : T275;
  assign T275 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T276;
  assign T276 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T277 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T278 = s2_recycle ? s2_req_tag : T279;
  assign T279 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T280;
  assign T280 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T281 = s2_nack_hit ? 1'h0 : T282;
  assign T282 = T302 & T283;
  assign T283 = T291 | T284;
  assign T284 = T288 | T285;
  assign T285 = T287 | T286;
  assign T286 = s2_req_cmd == 5'h4;
  assign T287 = s2_req_cmd[2'h3:2'h3];
  assign T288 = T290 | T289;
  assign T289 = s2_req_cmd == 5'h7;
  assign T290 = s2_req_cmd == 5'h1;
  assign T291 = T299 | T292;
  assign T292 = T296 | T293;
  assign T293 = T295 | T294;
  assign T294 = s2_req_cmd == 5'h4;
  assign T295 = s2_req_cmd[2'h3:2'h3];
  assign T296 = T298 | T297;
  assign T297 = s2_req_cmd == 5'h6;
  assign T298 = s2_req_cmd == 5'h0;
  assign T299 = T301 | T300;
  assign T300 = s2_req_cmd == 5'h3;
  assign T301 = s2_req_cmd == 5'h2;
  assign T302 = s2_valid_masked & T303;
  assign T303 = s2_hit ^ 1'h1;
  assign T304 = io_mem_probe_valid & T305;
  assign T305 = lrsc_valid ^ 1'h1;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_probe_ready = T306;
  assign T306 = prober_io_req_ready & T307;
  assign T307 = lrsc_valid ^ 1'h1;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_ordered = T308;
  assign T308 = T310 & T309;
  assign T309 = s2_valid ^ 1'h1;
  assign T310 = mshrs_io_fence_rdy & T311;
  assign T311 = s1_valid ^ 1'h1;
  assign io_cpu_xcpt_pf_st = T312;
  assign T312 = T313 & dtlb_io_resp_xcpt_st;
  assign T313 = T314 & s1_write;
  assign T314 = s1_req_phys ^ 1'h1;
  assign io_cpu_xcpt_pf_ld = T315;
  assign T315 = T316 & dtlb_io_resp_xcpt_ld;
  assign T316 = T317 & s1_read;
  assign T317 = s1_req_phys ^ 1'h1;
  assign io_cpu_xcpt_ma_st = T318;
  assign T318 = s1_write & misaligned;
  assign misaligned = T323 | T319;
  assign T319 = T322 & T320;
  assign T320 = T321 != 3'h0;
  assign T321 = s1_req_addr[2'h2:1'h0];
  assign T322 = s1_req_typ == 3'h3;
  assign T323 = T330 | T324;
  assign T324 = T327 & T325;
  assign T325 = T326 != 2'h0;
  assign T326 = s1_req_addr[1'h1:1'h0];
  assign T327 = T329 | T328;
  assign T328 = s1_req_typ == 3'h6;
  assign T329 = s1_req_typ == 3'h2;
  assign T330 = T333 & T331;
  assign T331 = T332 != 1'h0;
  assign T332 = s1_req_addr[1'h0:1'h0];
  assign T333 = T335 | T334;
  assign T334 = s1_req_typ == 3'h5;
  assign T335 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T336;
  assign T336 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T337;
  assign T337 = s1_replay & T338;
  assign T338 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_data_subword = T339;
  assign T339 = T340 | T443;
  assign T443 = {63'h0, s2_sc_fail};
  assign T340 = {T379, T341};
  assign T341 = s2_sc ? 8'h0 : T342;
  assign T342 = T378 ? T377 : T343;
  assign T343 = T344[3'h7:1'h0];
  assign T344 = {T369, T345};
  assign T345 = T368 ? T367 : T346;
  assign T346 = T347[4'hf:1'h0];
  assign T347 = {T352, T348};
  assign T348 = T351 ? T350 : T349;
  assign T349 = s2_data_word[5'h1f:1'h0];
  assign T350 = s2_data_word[6'h3f:6'h20];
  assign T351 = s2_req_addr[2'h2:2'h2];
  assign T352 = T364 ? T354 : T353;
  assign T353 = s2_data_word[6'h3f:6'h20];
  assign T354 = 32'h0 - T444;
  assign T444 = {31'h0, T355};
  assign T355 = T357 & T356;
  assign T356 = T348[5'h1f:5'h1f];
  assign T357 = T359 | T358;
  assign T358 = s2_req_typ == 3'h3;
  assign T359 = T361 | T360;
  assign T360 = s2_req_typ == 3'h2;
  assign T361 = T363 | T362;
  assign T362 = s2_req_typ == 3'h1;
  assign T363 = s2_req_typ == 3'h0;
  assign T364 = T366 | T365;
  assign T365 = s2_req_typ == 3'h6;
  assign T366 = s2_req_typ == 3'h2;
  assign T367 = T347[5'h1f:5'h10];
  assign T368 = s2_req_addr[1'h1:1'h1];
  assign T369 = T374 ? T371 : T370;
  assign T370 = T347[6'h3f:5'h10];
  assign T371 = 48'h0 - T445;
  assign T445 = {47'h0, T372};
  assign T372 = T357 & T373;
  assign T373 = T345[4'hf:4'hf];
  assign T374 = T376 | T375;
  assign T375 = s2_req_typ == 3'h5;
  assign T376 = s2_req_typ == 3'h1;
  assign T377 = T344[4'hf:4'h8];
  assign T378 = s2_req_addr[1'h0:1'h0];
  assign T379 = T384 ? T381 : T380;
  assign T380 = T344[6'h3f:4'h8];
  assign T381 = 56'h0 - T446;
  assign T446 = {55'h0, T382};
  assign T382 = T357 & T383;
  assign T383 = T341[3'h7:3'h7];
  assign T384 = s2_sc | T385;
  assign T385 = T387 | T386;
  assign T386 = s2_req_typ == 3'h4;
  assign T387 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_has_data = T388;
  assign T388 = T389 | s2_sc;
  assign T389 = T393 | T390;
  assign T390 = T392 | T391;
  assign T391 = s2_req_cmd == 5'h4;
  assign T392 = s2_req_cmd[2'h3:2'h3];
  assign T393 = T395 | T394;
  assign T394 = s2_req_cmd == 5'h6;
  assign T395 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T396;
  assign T396 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T347;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_valid = T397;
  assign T397 = T399 & T398;
  assign T398 = s2_data_correctable ^ 1'h1;
  assign T399 = s2_replay | T400;
  assign T400 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T401;
  assign T401 = block_miss ? 1'h0 : T402;
  assign T402 = T409 ? 1'h0 : T403;
  assign T403 = T408 ? 1'h0 : T404;
  assign T404 = T405 == 1'h0;
  assign T405 = T407 & T406;
  assign T406 = io_cpu_req_bits_phys ^ 1'h1;
  assign T407 = dtlb_io_req_ready ^ 1'h1;
  assign T408 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T409 = readArb_io_in_3_ready ^ 1'h1;
  assign T447 = reset ? 1'h0 : T410;
  assign T410 = T411 & s2_nack_miss;
  assign T411 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_req_bits_data( wbArb_io_out_bits_data ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_req_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type ),
       .io_release_bits_voluntary( wb_io_release_bits_voluntary )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T304 ),
       .io_req_bits_addr_block( io_mem_probe_bits_addr_block ),
       .io_req_bits_p_type( io_mem_probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_rep_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_data( prober_io_wb_req_bits_data ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_block_state_state( s2_hit_state_state )
  );
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T281 ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T270 ),
       .io_req_bits_old_meta_coh_state( T267 ),
       .io_req_bits_way_en( T441 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( io_mem_acquire_ready ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( mshrs_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( mshrs_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_is_builtin_type( mshrs_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( mshrs_io_mem_req_bits_union ),
       .io_refill_way_en( mshrs_io_refill_way_en ),
       .io_refill_addr( mshrs_io_refill_addr ),
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T263 ),
       .io_mem_grant_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_mem_grant_bits_data( FlowThroughSerializer_io_out_bits_data ),
       .io_mem_grant_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_data( mshrs_io_wb_req_bits_data ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_wb_req_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T250 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T249 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_req_bits_store( s1_write ),
       .io_resp_miss( dtlb_io_resp_miss ),
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dtlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dtlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dtlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dtlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T440 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T439 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T239 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 1'h1 ),
       .io_in_3_bits_addr( T438 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 1'h1 ),
       .io_in_1_bits_addr( T437 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 1'h1 ),
       .io_in_0_bits_addr( T436 ),
       .io_out_ready( T237 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T229 ),
       .io_in_1_bits_way_en( mshrs_io_refill_way_en ),
       .io_in_1_bits_addr( mshrs_io_refill_addr ),
       .io_in_1_bits_wmask( 2'h1 ),
       .io_in_1_bits_data( FlowThroughSerializer_io_out_bits_data ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T435 ),
       .io_in_0_bits_wmask( rowWMask ),
       .io_in_0_bits_data( T226 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T434 ),
       .io_cmd( s2_req_cmd ),
       .io_typ( s2_req_typ ),
       .io_lhs( T421 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  LockingArbiter_0 releaseArb(.clk(clk), .reset(reset),
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_1_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_in_0_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_out_ready( io_mem_release_ready ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr_block( releaseArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( releaseArb_io_out_bits_addr_beat ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type ),
       .io_out_bits_voluntary( releaseArb_io_out_bits_voluntary )
       //.io_chosen(  )
  );
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_out_ready( T8 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data ),
       .io_out_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( FlowThroughSerializer_io_out_bits_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_data( mshrs_io_wb_req_bits_data ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_1_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_data( prober_io_wb_req_bits_data ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_in_0_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_out_bits_data( wbArb_io_out_bits_data ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_out_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "DCache exception occurred - cache response not killed.");
    $finish;
  end
// synthesis translate_on
`endif
    R4 <= T5;
    if(T99) begin
      s2_req_data <= s1_req_data;
    end else if(T21) begin
      s2_req_data <= T19;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T20;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T30) begin
      s2_recycle_next <= s2_recycle_ecc;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T31;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T415;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T417;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T416;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_hit_state_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(reset) begin
      R90 <= 1'h0;
    end else begin
      R90 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R106 <= T422;
    if(T109) begin
      R111 <= T113;
    end
    if(T203) begin
      s2_store_bypass_data <= T116;
    end
    if(T119) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T120;
    end
    if(T135) begin
      lrsc_addr <= T134;
    end
    if(T149) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_invalidate_lr) begin
      lrsc_count <= 5'h0;
    end else if(T157) begin
      lrsc_count <= 5'h0;
    end else if(T155) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T154;
    end
    s3_req_data <= T427;
    if(T164) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T164) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T119) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T119) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T203) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T164) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R265 <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_repl_meta_coh_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_repl_meta_tag <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T410;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [26:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_prv,
    input  io_in_1_bits_store,
    input  io_in_1_bits_fetch,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [26:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_prv,
    input  io_in_0_bits_store,
    input  io_in_0_bits_fetch,
    input  io_out_ready,
    output io_out_valid,
    output[26:0] io_out_bits_addr,
    output[1:0] io_out_bits_prv,
    output io_out_bits_store,
    output io_out_bits_fetch,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T28;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire[26:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T28 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_fetch = T5;
  assign T5 = T6 ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T6 = chosen;
  assign io_out_bits_store = T7;
  assign T7 = T6 ? io_in_1_bits_store : io_in_0_bits_store;
  assign io_out_bits_prv = T8;
  assign T8 = T6 ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign io_out_bits_addr = T9;
  assign T9 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = last_grant < 1'h0;
  assign T19 = last_grant < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = last_grant < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [26:0] io_requestor_1_req_bits_addr,
    input [1:0] io_requestor_1_req_bits_prv,
    input  io_requestor_1_req_bits_store,
    input  io_requestor_1_req_bits_fetch,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[19:0] io_requestor_1_resp_bits_pte_ppn,
    output[2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
    output io_requestor_1_resp_bits_pte_d,
    output io_requestor_1_resp_bits_pte_r,
    output[3:0] io_requestor_1_resp_bits_pte_typ,
    output io_requestor_1_resp_bits_pte_v,
    output io_requestor_1_status_sd,
    output[30:0] io_requestor_1_status_zero2,
    output io_requestor_1_status_sd_rv32,
    output[8:0] io_requestor_1_status_zero1,
    output[4:0] io_requestor_1_status_vm,
    output io_requestor_1_status_mprv,
    output[1:0] io_requestor_1_status_xs,
    output[1:0] io_requestor_1_status_fs,
    output[1:0] io_requestor_1_status_prv3,
    output io_requestor_1_status_ie3,
    output[1:0] io_requestor_1_status_prv2,
    output io_requestor_1_status_ie2,
    output[1:0] io_requestor_1_status_prv1,
    output io_requestor_1_status_ie1,
    output[1:0] io_requestor_1_status_prv,
    output io_requestor_1_status_ie,
    output io_requestor_1_invalidate,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [26:0] io_requestor_0_req_bits_addr,
    input [1:0] io_requestor_0_req_bits_prv,
    input  io_requestor_0_req_bits_store,
    input  io_requestor_0_req_bits_fetch,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[19:0] io_requestor_0_resp_bits_pte_ppn,
    output[2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
    output io_requestor_0_resp_bits_pte_d,
    output io_requestor_0_resp_bits_pte_r,
    output[3:0] io_requestor_0_resp_bits_pte_typ,
    output io_requestor_0_resp_bits_pte_v,
    output io_requestor_0_status_sd,
    output[30:0] io_requestor_0_status_zero2,
    output io_requestor_0_status_sd_rv32,
    output[8:0] io_requestor_0_status_zero1,
    output[4:0] io_requestor_0_status_vm,
    output io_requestor_0_status_mprv,
    output[1:0] io_requestor_0_status_xs,
    output[1:0] io_requestor_0_status_fs,
    output[1:0] io_requestor_0_status_prv3,
    output io_requestor_0_status_ie3,
    output[1:0] io_requestor_0_status_prv2,
    output io_requestor_0_status_ie2,
    output[1:0] io_requestor_0_status_prv1,
    output io_requestor_0_status_ie1,
    output[1:0] io_requestor_0_status_prv,
    output io_requestor_0_status_ie,
    output io_requestor_0_invalidate,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [7:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_status_sd,
    input [30:0] io_dpath_status_zero2,
    input  io_dpath_status_sd_rv32,
    input [8:0] io_dpath_status_zero1,
    input [4:0] io_dpath_status_vm,
    input  io_dpath_status_mprv,
    input [1:0] io_dpath_status_xs,
    input [1:0] io_dpath_status_fs,
    input [1:0] io_dpath_status_prv3,
    input  io_dpath_status_ie3,
    input [1:0] io_dpath_status_prv2,
    input  io_dpath_status_ie2,
    input [1:0] io_dpath_status_prv1,
    input  io_dpath_status_ie1,
    input [1:0] io_dpath_status_prv,
    input  io_dpath_status_ie
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T232;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] count;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire pte_cache_hit;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[1:0] T26;
  reg  R27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T233;
  wire[1:0] T234;
  wire T235;
  wire[2:0] T36;
  wire T236;
  wire[1:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  reg [2:0] R45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire[5:0] T50;
  wire[1:0] T51;
  wire T52;
  wire[1:0] T237;
  wire T238;
  wire[1:0] T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  R78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[31:0] pte_addr;
  wire[28:0] T87;
  wire[28:0] T88;
  wire[8:0] vpn_idx;
  wire[8:0] T89;
  wire[8:0] T90;
  wire[8:0] T91;
  reg [26:0] r_req_addr;
  wire[26:0] T92;
  wire T93;
  wire[8:0] T94;
  wire[17:0] T95;
  wire T96;
  wire[1:0] T97;
  wire[8:0] T98;
  wire[26:0] T99;
  wire T100;
  reg [19:0] r_pte_ppn;
  wire[19:0] T101;
  wire[19:0] T102;
  wire[19:0] T103;
  wire[19:0] T104;
  wire[19:0] T105;
  wire T106;
  wire T107;
  wire set_dirty_bit;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg  r_req_store;
  wire T112;
  wire T113;
  wire T114;
  wire perm_ok;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  r_req_fetch;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  reg [1:0] r_req_prv;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire[19:0] pte_cache_data;
  wire[19:0] T150;
  wire[19:0] T151;
  reg [19:0] T152 [2:0];
  wire[19:0] T153;
  wire T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire[19:0] T158;
  wire[19:0] T159;
  wire[19:0] T160;
  wire T161;
  wire[19:0] T162;
  wire[19:0] T163;
  wire T164;
  wire[31:0] T165;
  reg [31:0] T166 [2:0];
  wire[31:0] T167;
  wire T168;
  wire T169;
  wire[1:0] T170;
  wire T171;
  wire[31:0] T172;
  wire T173;
  wire[31:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[2:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[63:0] T243;
  wire[29:0] T198;
  wire[29:0] T199;
  wire[5:0] T200;
  wire[4:0] T201;
  wire pte_wdata_v;
  wire[3:0] pte_wdata_typ;
  wire pte_wdata_r;
  wire[23:0] T202;
  wire[3:0] T203;
  wire pte_wdata_d;
  wire[2:0] pte_wdata_reserved_for_software;
  wire[19:0] pte_wdata_ppn;
  wire[4:0] T204;
  wire T205;
  wire[39:0] T244;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  reg  r_pte_v;
  wire T210;
  reg [3:0] r_pte_typ;
  wire[3:0] T211;
  reg  r_pte_r;
  wire T212;
  reg  r_pte_d;
  wire T213;
  reg [2:0] r_pte_reserved_for_software;
  wire[2:0] T214;
  wire[2:0] T215;
  wire[19:0] T245;
  wire[27:0] resp_ppn;
  wire[27:0] T216;
  wire[27:0] T217;
  wire[17:0] T218;
  wire[9:0] T219;
  wire[27:0] T220;
  wire[8:0] T221;
  wire[18:0] T222;
  wire T223;
  wire[1:0] T224;
  wire[27:0] r_resp_ppn;
  wire T225;
  wire resp_err;
  wire T226;
  wire T227;
  reg  r_req_dest;
  wire T228;
  wire resp_val;
  wire T229;
  wire[19:0] T246;
  wire T230;
  wire T231;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[26:0] arb_io_out_bits_addr;
  wire[1:0] arb_io_out_bits_prv;
  wire arb_io_out_bits_store;
  wire arb_io_out_bits_fetch;
  wire arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    R27 = {1{$random}};
    R45 = {1{$random}};
    R73 = {1{$random}};
    R78 = {1{$random}};
    r_req_addr = {1{$random}};
    r_pte_ppn = {1{$random}};
    r_req_store = {1{$random}};
    r_req_fetch = {1{$random}};
    r_req_prv = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T152[initvar] = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T166[initvar] = {1{$random}};
    r_pte_v = {1{$random}};
    r_pte_typ = {1{$random}};
    r_pte_r = {1{$random}};
    r_pte_d = {1{$random}};
    r_pte_reserved_for_software = {1{$random}};
    r_req_dest = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
//  assign io_mem_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = state == 3'h0;
  assign T232 = reset ? 3'h0 : T1;
  assign T1 = T197 ? 3'h0 : T2;
  assign T2 = T196 ? 3'h0 : T3;
  assign T3 = T195 ? 3'h1 : T4;
  assign T4 = T193 ? 3'h3 : T5;
  assign T5 = T191 ? 3'h4 : T6;
  assign T6 = T188 ? T187 : T7;
  assign T7 = T182 ? 3'h1 : T8;
  assign T8 = T181 ? 3'h6 : T9;
  assign T9 = T179 ? 3'h1 : T10;
  assign T10 = T176 ? 3'h2 : T11;
  assign T11 = T15 ? 3'h1 : T12;
  assign T12 = T13 ? 3'h1 : state;
  assign T13 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T15 = T175 & T16;
  assign T16 = pte_cache_hit & T17;
  assign T17 = count < 2'h2;
  assign T18 = T182 ? T22 : T19;
  assign T19 = T15 ? T21 : T20;
  assign T20 = T14 ? 2'h0 : count;
  assign T21 = count + 2'h1;
  assign T22 = count + 2'h1;
  assign pte_cache_hit = T23 != 3'h0;
  assign T23 = T83 & T24;
  assign T24 = T25;
  assign T25 = {R78, T26};
  assign T26 = {R73, R27};
  assign T28 = T72 ? 1'h0 : T29;
  assign T29 = T30 ? 1'h1 : R27;
  assign T30 = T65 & T31;
  assign T31 = T32[1'h0:1'h0];
  assign T32 = 1'h1 << T33;
  assign T33 = T34;
  assign T34 = T64 ? T37 : T233;
  assign T233 = T236 ? 1'h0 : T234;
  assign T234 = T235 ? 1'h1 : 2'h2;
  assign T235 = T36[1'h1:1'h1];
  assign T36 = ~ T24;
  assign T236 = T36[1'h0:1'h0];
  assign T37 = T38[1'h1:1'h0];
  assign T38 = {T62, T39};
  assign T39 = T44 & T40;
  assign T40 = T41 - 1'h1;
  assign T41 = 1'h1 << T42;
  assign T42 = T43 + 2'h1;
  assign T43 = T62 - T62;
  assign T44 = R45 >> T62;
  assign T46 = T60 ? T47 : R45;
  assign T47 = T55 | T48;
  assign T48 = T54 ? 3'h0 : T49;
  assign T49 = T50[2'h2:1'h0];
  assign T50 = 3'h1 << T51;
  assign T51 = {1'h1, T52};
  assign T52 = T237[1'h1:1'h1];
  assign T237 = {T242, T238};
  assign T238 = T239[1'h1:1'h1];
  assign T239 = T241 | T240;
  assign T240 = T23[1'h1:1'h0];
  assign T241 = T23[2'h2:2'h2];
  assign T242 = T241 != 1'h0;
  assign T54 = T237[1'h0:1'h0];
  assign T55 = T57 & T56;
  assign T56 = ~ T49;
  assign T57 = T59 | T58;
  assign T58 = T52 ? 3'h0 : 3'h2;
  assign T59 = R45 & 3'h5;
  assign T60 = pte_cache_hit & T61;
  assign T61 = state == 3'h1;
  assign T62 = {1'h1, T63};
  assign T63 = R45[1'h1:1'h1];
  assign T64 = T24 == 3'h7;
  assign T65 = T67 & T66;
  assign T66 = pte_cache_hit ^ 1'h1;
  assign T67 = io_mem_resp_valid & T68;
  assign T68 = T71 & T69;
  assign T69 = T70 < 4'h2;
  assign T70 = io_mem_resp_bits_data[3'h4:1'h1];
  assign T71 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T72 = reset | io_dpath_invalidate;
  assign T74 = T72 ? 1'h0 : T75;
  assign T75 = T76 ? 1'h1 : R73;
  assign T76 = T65 & T77;
  assign T77 = T32[1'h1:1'h1];
  assign T79 = T72 ? 1'h0 : T80;
  assign T80 = T81 ? 1'h1 : R78;
  assign T81 = T65 & T82;
  assign T82 = T32[2'h2:2'h2];
  assign T83 = T84;
  assign T84 = {T173, T85};
  assign T85 = {T171, T86};
  assign T86 = T165 == pte_addr;
  assign pte_addr = T87 << 2'h3;
  assign T87 = T88;
  assign T88 = {r_pte_ppn, vpn_idx};
  assign vpn_idx = T100 ? T98 : T89;
  assign T89 = T96 ? T94 : T90;
  assign T90 = T91[4'h8:1'h0];
  assign T91 = r_req_addr >> 5'h12;
  assign T92 = T93 ? arb_io_out_bits_addr : r_req_addr;
  assign T93 = T0 & arb_io_out_valid;
  assign T94 = T95[4'h8:1'h0];
  assign T95 = r_req_addr >> 4'h9;
  assign T96 = T97[1'h0:1'h0];
  assign T97 = count;
  assign T98 = T99[4'h8:1'h0];
  assign T99 = r_req_addr >> 1'h0;
  assign T100 = T97[1'h1:1'h1];
  assign T101 = T15 ? pte_cache_data : T102;
  assign T102 = T106 ? T105 : T103;
  assign T103 = T93 ? T104 : r_pte_ppn;
  assign T104 = io_dpath_ptbr[5'h1f:4'hc];
  assign T105 = io_mem_resp_bits_data[5'h1d:4'ha];
  assign T106 = T148 & T107;
  assign T107 = set_dirty_bit ^ 1'h1;
  assign set_dirty_bit = perm_ok & T108;
  assign T108 = T113 | T109;
  assign T109 = r_req_store & T110;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_mem_resp_bits_data[3'h6:3'h6];
  assign T112 = T93 ? arb_io_out_bits_store : r_req_store;
  assign T113 = T114 ^ 1'h1;
  assign T114 = io_mem_resp_bits_data[3'h5:3'h5];
  assign perm_ok = T146 ? T134 : T115;
  assign T115 = r_req_fetch ? T127 : T116;
  assign T116 = r_req_store ? T121 : T117;
  assign T117 = T119 & T118;
  assign T118 = T70 < 4'h8;
  assign T119 = T71 & T120;
  assign T120 = 4'h2 <= T70;
  assign T121 = T123 & T122;
  assign T122 = T70[1'h0:1'h0];
  assign T123 = T125 & T124;
  assign T124 = T70 < 4'h8;
  assign T125 = T71 & T126;
  assign T126 = 4'h2 <= T70;
  assign T127 = T129 & T128;
  assign T128 = T70[1'h1:1'h1];
  assign T129 = T131 & T130;
  assign T130 = T70 < 4'h8;
  assign T131 = T71 & T132;
  assign T132 = 4'h2 <= T70;
  assign T133 = T93 ? arb_io_out_bits_fetch : r_req_fetch;
  assign T134 = r_req_fetch ? T142 : T135;
  assign T135 = r_req_store ? T138 : T136;
  assign T136 = T71 & T137;
  assign T137 = 4'h2 <= T70;
  assign T138 = T140 & T139;
  assign T139 = T70[1'h0:1'h0];
  assign T140 = T71 & T141;
  assign T141 = 4'h2 <= T70;
  assign T142 = T144 & T143;
  assign T143 = T70[1'h1:1'h1];
  assign T144 = T71 & T145;
  assign T145 = 4'h4 <= T70;
  assign T146 = r_req_prv[1'h0:1'h0];
  assign T147 = T93 ? arb_io_out_bits_prv : r_req_prv;
  assign T148 = io_mem_resp_valid & T149;
  assign T149 = state == 3'h2;
  assign pte_cache_data = T158 | T150;
  assign T150 = T157 ? T151 : 20'h0;
  assign T151 = T152[2'h2];
  assign T154 = T65 & T155;
  assign T155 = T156 < 2'h3;
  assign T156 = T34[1'h1:1'h0];
  assign T157 = T23[2'h2:2'h2];
  assign T158 = T162 | T159;
  assign T159 = T161 ? T160 : 20'h0;
  assign T160 = T152[2'h1];
  assign T161 = T23[1'h1:1'h1];
  assign T162 = T164 ? T163 : 20'h0;
  assign T163 = T152[2'h0];
  assign T164 = T23[1'h0:1'h0];
  assign T165 = T166[2'h0];
  assign T168 = T65 & T169;
  assign T169 = T170 < 2'h3;
  assign T170 = T34[1'h1:1'h0];
  assign T171 = T172 == pte_addr;
  assign T172 = T166[2'h1];
  assign T173 = T174 == pte_addr;
  assign T174 = T166[2'h2];
  assign T175 = 3'h1 == state;
  assign T176 = T175 & T177;
  assign T177 = T178 & io_mem_req_ready;
  assign T178 = T16 ^ 1'h1;
  assign T179 = T180 & io_mem_resp_bits_nack;
  assign T180 = 3'h2 == state;
  assign T181 = T180 & io_mem_resp_valid;
  assign T182 = T181 & T183;
  assign T183 = T185 & T184;
  assign T184 = count < 2'h2;
  assign T185 = T71 & T186;
  assign T186 = T70 < 4'h2;
  assign T187 = set_dirty_bit ? 3'h3 : 3'h5;
  assign T188 = T181 & T189;
  assign T189 = T71 & T190;
  assign T190 = 4'h2 <= T70;
  assign T191 = T192 & io_mem_req_ready;
  assign T192 = 3'h3 == state;
  assign T193 = T194 & io_mem_resp_bits_nack;
  assign T194 = 3'h4 == state;
  assign T195 = T194 & io_mem_resp_valid;
  assign T196 = 3'h5 == state;
  assign T197 = 3'h6 == state;
  assign io_mem_req_bits_data = T243;
  assign T243 = {34'h0, T198};
  assign T198 = T199;
  assign T199 = {T202, T200};
  assign T200 = {pte_wdata_r, T201};
  assign T201 = {pte_wdata_typ, pte_wdata_v};
  assign pte_wdata_v = 1'h0;
  assign pte_wdata_typ = 4'h0;
  assign pte_wdata_r = 1'h1;
  assign T202 = {pte_wdata_ppn, T203};
  assign T203 = {pte_wdata_reserved_for_software, pte_wdata_d};
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_reserved_for_software = 3'h0;
  assign pte_wdata_ppn = 20'h0;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_cmd = T204;
  assign T204 = T205 ? 5'ha : 5'h0;
  assign T205 = state == 3'h3;
  assign io_mem_req_bits_addr = T244;
  assign T244 = {8'h0, pte_addr};
  assign io_mem_req_valid = T206;
  assign T206 = T15 ? 1'h0 : T207;
  assign T207 = T209 | T208;
  assign T208 = state == 3'h3;
  assign T209 = state == 3'h1;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_ie = io_dpath_status_ie;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_0_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_0_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_0_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_0_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_0_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign T210 = T106 ? T71 : r_pte_v;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign T211 = T106 ? T70 : r_pte_typ;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign T212 = T106 ? T114 : r_pte_r;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign T213 = T106 ? T111 : r_pte_d;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign T214 = T106 ? T215 : r_pte_reserved_for_software;
  assign T215 = io_mem_resp_bits_data[4'h9:3'h7];
  assign io_requestor_0_resp_bits_pte_ppn = T245;
  assign T245 = resp_ppn[5'h13:1'h0];
  assign resp_ppn = T225 ? r_resp_ppn : T216;
  assign T216 = T223 ? T220 : T217;
  assign T217 = {T219, T218};
  assign T218 = r_req_addr[5'h11:1'h0];
  assign T219 = r_resp_ppn >> 5'h12;
  assign T220 = {T222, T221};
  assign T221 = r_req_addr[4'h8:1'h0];
  assign T222 = r_resp_ppn >> 4'h9;
  assign T223 = T224[1'h0:1'h0];
  assign T224 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hc;
  assign T225 = T224[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = state == 3'h6;
  assign io_requestor_0_resp_valid = T226;
  assign T226 = resp_val & T227;
  assign T227 = r_req_dest == 1'h0;
  assign T228 = T93 ? arb_io_chosen : r_req_dest;
  assign resp_val = T229 | resp_err;
  assign T229 = state == 3'h5;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_ie = io_dpath_status_ie;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_1_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_1_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_1_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_1_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_1_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_ppn = T246;
  assign T246 = resp_ppn[5'h13:1'h0];
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T230;
  assign T230 = resp_val & T231;
  assign T231 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits_addr( io_requestor_1_req_bits_addr ),
       .io_in_1_bits_prv( io_requestor_1_req_bits_prv ),
       .io_in_1_bits_store( io_requestor_1_req_bits_store ),
       .io_in_1_bits_fetch( io_requestor_1_req_bits_fetch ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits_addr( io_requestor_0_req_bits_addr ),
       .io_in_0_bits_prv( io_requestor_0_req_bits_prv ),
       .io_in_0_bits_store( io_requestor_0_req_bits_store ),
       .io_in_0_bits_fetch( io_requestor_0_req_bits_fetch ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits_addr( arb_io_out_bits_addr ),
       .io_out_bits_prv( arb_io_out_bits_prv ),
       .io_out_bits_store( arb_io_out_bits_store ),
       .io_out_bits_fetch( arb_io_out_bits_fetch ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T197) begin
      state <= 3'h0;
    end else if(T196) begin
      state <= 3'h0;
    end else if(T195) begin
      state <= 3'h1;
    end else if(T193) begin
      state <= 3'h3;
    end else if(T191) begin
      state <= 3'h4;
    end else if(T188) begin
      state <= T187;
    end else if(T182) begin
      state <= 3'h1;
    end else if(T181) begin
      state <= 3'h6;
    end else if(T179) begin
      state <= 3'h1;
    end else if(T176) begin
      state <= 3'h2;
    end else if(T15) begin
      state <= 3'h1;
    end else if(T13) begin
      state <= 3'h1;
    end
    if(T182) begin
      count <= T22;
    end else if(T15) begin
      count <= T21;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T72) begin
      R27 <= 1'h0;
    end else if(T30) begin
      R27 <= 1'h1;
    end
    if(T60) begin
      R45 <= T47;
    end
    if(T72) begin
      R73 <= 1'h0;
    end else if(T76) begin
      R73 <= 1'h1;
    end
    if(T72) begin
      R78 <= 1'h0;
    end else if(T81) begin
      R78 <= 1'h1;
    end
    if(T93) begin
      r_req_addr <= arb_io_out_bits_addr;
    end
    if(T15) begin
      r_pte_ppn <= pte_cache_data;
    end else if(T106) begin
      r_pte_ppn <= T105;
    end else if(T93) begin
      r_pte_ppn <= T104;
    end
    if(T93) begin
      r_req_store <= arb_io_out_bits_store;
    end
    if(T93) begin
      r_req_fetch <= arb_io_out_bits_fetch;
    end
    if(T93) begin
      r_req_prv <= arb_io_out_bits_prv;
    end
    if (T154)
      T152[T34] <= T105;
    if (T168)
      T166[T34] <= pte_addr;
    if(T106) begin
      r_pte_v <= T71;
    end
    if(T106) begin
      r_pte_typ <= T70;
    end
    if(T106) begin
      r_pte_r <= T114;
    end
    if(T106) begin
      r_pte_d <= T111;
    end
    if(T106) begin
      r_pte_reserved_for_software <= T215;
    end
    if(T93) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [11:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [2:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output io_csr_replay,
    output io_csr_stall,
    output io_csr_xcpt,
    output io_eret,
    output io_status_sd,
    output[30:0] io_status_zero2,
    output io_status_sd_rv32,
    output[8:0] io_status_zero1,
    output[4:0] io_status_vm,
    output io_status_mprv,
    output[1:0] io_status_xs,
    output[1:0] io_status_fs,
    output[1:0] io_status_prv3,
    output io_status_ie3,
    output[1:0] io_status_prv2,
    output io_status_ie2,
    output[1:0] io_status_prv1,
    output io_status_ie1,
    output[1:0] io_status_prv,
    output io_status_ie,
    output[31:0] io_ptbr,
    output[39:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input [39:0] io_pc,
    output io_fatc,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [25:0] io_rocc_imem_acquire_bits_addr_block,
    input  io_rocc_imem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_imem_acquire_bits_addr_beat,
    input [127:0] io_rocc_imem_acquire_bits_data,
    input  io_rocc_imem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_imem_acquire_bits_a_type,
    input [16:0] io_rocc_imem_acquire_bits_union,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_addr_beat
    //output[127:0] io_rocc_imem_grant_bits_data
    //output io_rocc_imem_grant_bits_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_manager_xact_id
    //output io_rocc_imem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_imem_grant_bits_g_type
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [25:0] io_rocc_dmem_acquire_bits_addr_block,
    input  io_rocc_dmem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_dmem_acquire_bits_addr_beat,
    input [127:0] io_rocc_dmem_acquire_bits_data,
    input  io_rocc_dmem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_dmem_acquire_bits_a_type,
    input [16:0] io_rocc_dmem_acquire_bits_union,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_addr_beat
    //output[127:0] io_rocc_dmem_grant_bits_data
    //output io_rocc_dmem_grant_bits_client_xact_id
    //output[2:0] io_rocc_dmem_grant_bits_manager_xact_id
    //output io_rocc_dmem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_dmem_grant_bits_g_type
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    //output io_rocc_exception
    output io_interrupt,
    output[63:0] io_interrupt_cause
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T882;
  wire csr_xcpt;
  wire insn_break;
  wire system_insn;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire insn_call;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire priv_sufficient;
  reg [1:0] reg_mstatus_prv;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  reg [1:0] reg_mstatus_prv1;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  reg [1:0] reg_mstatus_prv2;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[63:0] wdata;
  wire[63:0] T38;
  wire[63:0] T39;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T40;
  wire[63:0] T41;
  wire T42;
  wire host_pcr_req_fire;
  wire T43;
  wire cpu_ren;
  wire T44;
  wire T45;
  reg  host_pcr_req_valid;
  wire T46;
  wire T47;
  wire[63:0] T48;
  wire T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[11:0] addr;
  reg [11:0] host_pcr_bits_addr;
  wire[11:0] T62;
  wire wen;
  wire T63;
  reg  host_pcr_bits_rw;
  wire T64;
  wire T65;
  wire T66;
  wire read_only;
  wire[1:0] T67;
  wire cpu_wen;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[1:0] T883;
  wire T77;
  wire T78;
  wire T79;
  wire insn_ret;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire insn_redirect_trap;
  wire maybe_insn_redirect_trap;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[1:0] csr_addr_priv;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire fp_csr;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire addr_valid;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[2:0] T884;
  wire[3:0] T885;
  wire[1:0] T215;
  wire[1:0] T216;
  wire[1:0] T886;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] T220;
  wire[63:0] T221;
  wire T222;
  wire T223;
  wire T224;
  reg  reg_mstatus_ie;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  reg  reg_mstatus_ie1;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  reg  reg_mstatus_ie2;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  reg  reg_mip_ssip;
  wire T887;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg  reg_mie_ssip;
  wire T888;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  reg  reg_mip_msip;
  wire T889;
  wire T265;
  wire T266;
  wire T267;
  reg  reg_mie_msip;
  wire T890;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  reg  reg_mip_stip;
  wire T891;
  wire T276;
  wire T277;
  reg  reg_mie_stip;
  wire T892;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  reg  reg_mip_mtip;
  wire T893;
  wire T288;
  wire T289;
  wire T290;
  reg [63:0] reg_time;
  wire[63:0] T291;
  wire T292;
  reg [63:0] reg_mtimecmp;
  wire[63:0] T293;
  wire T294;
  reg  reg_mie_mtip;
  wire T894;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  reg [63:0] reg_fromhost;
  wire[63:0] T895;
  wire[63:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  reg [2:0] reg_frm;
  wire[2:0] T896;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T897;
  wire T312;
  wire[63:0] T898;
  wire[58:0] T313;
  wire T314;
  wire[63:0] T315;
  reg [5:0] R316;
  wire[5:0] T899;
  wire[5:0] T317;
  wire[6:0] T318;
  wire[6:0] T900;
  reg [57:0] R319;
  wire[57:0] T901;
  wire[57:0] T320;
  wire[57:0] T321;
  wire T322;
  wire insn_sfence_vm;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[39:0] T330;
  wire[39:0] T331;
  wire[39:0] T332;
  reg [39:0] reg_sepc;
  wire[39:0] T902;
  wire[63:0] T333;
  wire[63:0] T903;
  wire[39:0] T334;
  wire[63:0] T335;
  wire[63:0] T336;
  wire[63:0] T337;
  wire T338;
  reg [39:0] reg_mepc;
  wire[39:0] T904;
  wire[63:0] T339;
  wire[63:0] T905;
  wire[39:0] T340;
  wire[39:0] T341;
  wire[39:0] T342;
  wire[39:0] T343;
  wire[63:0] T344;
  wire[63:0] T345;
  wire[63:0] T346;
  wire T347;
  wire T348;
  wire[39:0] T349;
  reg [38:0] reg_stvec;
  wire[38:0] T906;
  wire[63:0] T350;
  wire[63:0] T907;
  wire[63:0] T351;
  wire[63:0] T352;
  wire[63:0] T353;
  wire T354;
  wire T355;
  wire[39:0] T908;
  wire[8:0] T356;
  wire[8:0] T909;
  wire[7:0] T357;
  wire T358;
  reg [31:0] reg_sptbr;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[19:0] T361;
  wire T362;
  reg  reg_mstatus_ie3;
  wire T363;
  reg [1:0] reg_mstatus_prv3;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[1:0] T910;
  wire T366;
  reg [1:0] reg_mstatus_fs;
  wire[1:0] T367;
  wire[1:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T911;
  wire T373;
  reg [1:0] reg_mstatus_xs;
  wire[1:0] T374;
  reg  reg_mstatus_mprv;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  reg [4:0] reg_mstatus_vm;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire T384;
  wire T385;
  wire[4:0] T386;
  wire T387;
  wire T388;
  reg [8:0] reg_mstatus_zero1;
  wire[8:0] T389;
  reg  reg_mstatus_sd_rv32;
  wire T390;
  reg [30:0] reg_mstatus_zero2;
  wire[30:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  reg  reg_wfi;
  wire T912;
  wire T396;
  wire T397;
  wire insn_wfi;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire some_interrupt_pending;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire[63:0] T421;
  wire[63:0] T422;
  wire[63:0] T423;
  reg [5:0] R424;
  wire[5:0] T913;
  wire[5:0] T425;
  wire[5:0] T426;
  wire[6:0] T427;
  wire[6:0] T914;
  wire T428;
  reg [57:0] R429;
  wire[57:0] T915;
  wire[57:0] T430;
  wire[57:0] T431;
  wire T432;
  wire T433;
  wire[63:0] T434;
  wire[63:0] T435;
  wire[63:0] T436;
  reg [5:0] R437;
  wire[5:0] T916;
  wire[5:0] T438;
  wire[5:0] T439;
  wire[6:0] T440;
  wire[6:0] T917;
  wire T441;
  reg [57:0] R442;
  wire[57:0] T918;
  wire[57:0] T443;
  wire[57:0] T444;
  wire T445;
  wire T446;
  wire[63:0] T447;
  wire[63:0] T448;
  wire[63:0] T449;
  reg [5:0] R450;
  wire[5:0] T919;
  wire[5:0] T451;
  wire[5:0] T452;
  wire[6:0] T453;
  wire[6:0] T920;
  wire T454;
  reg [57:0] R455;
  wire[57:0] T921;
  wire[57:0] T456;
  wire[57:0] T457;
  wire T458;
  wire T459;
  wire[63:0] T460;
  wire[63:0] T461;
  wire[63:0] T462;
  reg [5:0] R463;
  wire[5:0] T922;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[6:0] T466;
  wire[6:0] T923;
  wire T467;
  reg [57:0] R468;
  wire[57:0] T924;
  wire[57:0] T469;
  wire[57:0] T470;
  wire T471;
  wire T472;
  wire[63:0] T473;
  wire[63:0] T474;
  wire[63:0] T475;
  reg [5:0] R476;
  wire[5:0] T925;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[6:0] T479;
  wire[6:0] T926;
  wire T480;
  reg [57:0] R481;
  wire[57:0] T927;
  wire[57:0] T482;
  wire[57:0] T483;
  wire T484;
  wire T485;
  wire[63:0] T486;
  wire[63:0] T487;
  wire[63:0] T488;
  reg [5:0] R489;
  wire[5:0] T928;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[6:0] T492;
  wire[6:0] T929;
  wire T493;
  reg [57:0] R494;
  wire[57:0] T930;
  wire[57:0] T495;
  wire[57:0] T496;
  wire T497;
  wire T498;
  wire[63:0] T499;
  wire[63:0] T500;
  wire[63:0] T501;
  reg [5:0] R502;
  wire[5:0] T931;
  wire[5:0] T503;
  wire[5:0] T504;
  wire[6:0] T505;
  wire[6:0] T932;
  wire T506;
  reg [57:0] R507;
  wire[57:0] T933;
  wire[57:0] T508;
  wire[57:0] T509;
  wire T510;
  wire T511;
  wire[63:0] T512;
  wire[63:0] T513;
  wire[63:0] T514;
  reg [5:0] R515;
  wire[5:0] T934;
  wire[5:0] T516;
  wire[5:0] T517;
  wire[6:0] T518;
  wire[6:0] T935;
  wire T519;
  reg [57:0] R520;
  wire[57:0] T936;
  wire[57:0] T521;
  wire[57:0] T522;
  wire T523;
  wire T524;
  wire[63:0] T525;
  wire[63:0] T526;
  wire[63:0] T527;
  reg [5:0] R528;
  wire[5:0] T937;
  wire[5:0] T529;
  wire[5:0] T530;
  wire[6:0] T531;
  wire[6:0] T938;
  wire T532;
  reg [57:0] R533;
  wire[57:0] T939;
  wire[57:0] T534;
  wire[57:0] T535;
  wire T536;
  wire T537;
  wire[63:0] T538;
  wire[63:0] T539;
  wire[63:0] T540;
  reg [5:0] R541;
  wire[5:0] T940;
  wire[5:0] T542;
  wire[5:0] T543;
  wire[6:0] T544;
  wire[6:0] T941;
  wire T545;
  reg [57:0] R546;
  wire[57:0] T942;
  wire[57:0] T547;
  wire[57:0] T548;
  wire T549;
  wire T550;
  wire[63:0] T551;
  wire[63:0] T552;
  wire[63:0] T553;
  reg [5:0] R554;
  wire[5:0] T943;
  wire[5:0] T555;
  wire[5:0] T556;
  wire[6:0] T557;
  wire[6:0] T944;
  wire T558;
  reg [57:0] R559;
  wire[57:0] T945;
  wire[57:0] T560;
  wire[57:0] T561;
  wire T562;
  wire T563;
  wire[63:0] T564;
  wire[63:0] T565;
  wire[63:0] T566;
  reg [5:0] R567;
  wire[5:0] T946;
  wire[5:0] T568;
  wire[5:0] T569;
  wire[6:0] T570;
  wire[6:0] T947;
  wire T571;
  reg [57:0] R572;
  wire[57:0] T948;
  wire[57:0] T573;
  wire[57:0] T574;
  wire T575;
  wire T576;
  wire[63:0] T577;
  wire[63:0] T578;
  wire[63:0] T579;
  reg [5:0] R580;
  wire[5:0] T949;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[6:0] T583;
  wire[6:0] T950;
  wire T584;
  reg [57:0] R585;
  wire[57:0] T951;
  wire[57:0] T586;
  wire[57:0] T587;
  wire T588;
  wire T589;
  wire[63:0] T590;
  wire[63:0] T591;
  wire[63:0] T592;
  reg [5:0] R593;
  wire[5:0] T952;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[6:0] T596;
  wire[6:0] T953;
  wire T597;
  reg [57:0] R598;
  wire[57:0] T954;
  wire[57:0] T599;
  wire[57:0] T600;
  wire T601;
  wire T602;
  wire[63:0] T603;
  wire[63:0] T604;
  wire[63:0] T605;
  reg [5:0] R606;
  wire[5:0] T955;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[6:0] T609;
  wire[6:0] T956;
  wire T610;
  reg [57:0] R611;
  wire[57:0] T957;
  wire[57:0] T612;
  wire[57:0] T613;
  wire T614;
  wire T615;
  wire[63:0] T616;
  wire[63:0] T617;
  wire[63:0] T618;
  reg [5:0] R619;
  wire[5:0] T958;
  wire[5:0] T620;
  wire[5:0] T621;
  wire[6:0] T622;
  wire[6:0] T959;
  wire T623;
  reg [57:0] R624;
  wire[57:0] T960;
  wire[57:0] T625;
  wire[57:0] T626;
  wire T627;
  wire T628;
  wire[63:0] T629;
  wire[63:0] T630;
  wire[63:0] T631;
  wire[24:0] T632;
  wire[24:0] T961;
  wire T633;
  wire[63:0] T634;
  wire[63:0] T635;
  wire[63:0] T636;
  wire[23:0] T637;
  wire[23:0] T962;
  wire T638;
  wire[63:0] T639;
  wire[63:0] T640;
  wire[63:0] T963;
  wire[31:0] T641;
  wire[63:0] T642;
  wire[63:0] T643;
  wire[63:0] T644;
  reg [39:0] reg_sbadaddr;
  wire[39:0] T645;
  reg [39:0] reg_mbadaddr;
  wire[39:0] T646;
  wire[39:0] T647;
  wire[39:0] T648;
  wire[39:0] T649;
  wire[38:0] T650;
  wire T651;
  wire T652;
  wire[24:0] T653;
  wire T654;
  wire T655;
  wire[38:0] T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire[39:0] T665;
  wire T666;
  wire[23:0] T667;
  wire[23:0] T964;
  wire T668;
  wire[63:0] T669;
  wire[63:0] T670;
  reg [63:0] reg_scause;
  wire[63:0] T671;
  reg [63:0] reg_mcause;
  wire[63:0] T672;
  wire[63:0] T673;
  wire[63:0] T674;
  wire[63:0] T675;
  wire[63:0] T676;
  wire T677;
  wire T678;
  wire[63:0] T965;
  wire[3:0] T679;
  wire[3:0] T966;
  wire T680;
  wire[63:0] T681;
  wire T682;
  wire[63:0] T683;
  wire[63:0] T684;
  reg [63:0] reg_sscratch;
  wire[63:0] T685;
  wire T686;
  wire[63:0] T687;
  wire[63:0] T967;
  wire[7:0] T688;
  wire[7:0] T689;
  wire[7:0] T690;
  wire[3:0] T691;
  wire[1:0] T692;
  wire T693;
  wire T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire[3:0] T698;
  wire[1:0] T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire T703;
  wire T704;
  wire[63:0] T705;
  wire[63:0] T968;
  wire[7:0] T706;
  wire[7:0] T707;
  wire[7:0] T708;
  wire[3:0] T709;
  wire[1:0] T710;
  wire T711;
  wire T712;
  wire[1:0] T713;
  wire T714;
  wire T715;
  wire[3:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire[1:0] T720;
  wire T721;
  wire T722;
  wire[63:0] T723;
  wire[63:0] T724;
  wire[63:0] T725;
  wire[63:0] T726;
  wire[13:0] T727;
  wire[3:0] T728;
  wire[2:0] T729;
  wire T730;
  wire T731;
  wire[63:0] read_mstatus;
  wire[63:0] T732;
  wire[11:0] T733;
  wire[5:0] T734;
  wire[2:0] T735;
  wire[2:0] T736;
  wire[5:0] T737;
  wire[2:0] T738;
  wire[2:0] T739;
  wire[51:0] T740;
  wire[9:0] T741;
  wire[3:0] T742;
  wire[5:0] T743;
  wire[41:0] T744;
  wire[9:0] T745;
  wire[31:0] T746;
  wire[1:0] T747;
  wire T748;
  wire T749;
  wire[9:0] T750;
  wire[7:0] T751;
  wire T752;
  wire T753;
  wire[6:0] T754;
  wire[1:0] T755;
  wire[1:0] T756;
  wire[49:0] T757;
  wire[16:0] T758;
  wire[2:0] T759;
  wire[1:0] T760;
  wire[1:0] T761;
  wire T762;
  wire T763;
  wire[13:0] T764;
  wire[32:0] T765;
  wire[31:0] T766;
  wire T767;
  wire T768;
  wire[30:0] T769;
  wire T770;
  wire T771;
  wire[63:0] T772;
  wire[63:0] T773;
  wire[63:0] T774;
  wire[63:0] T775;
  reg [63:0] reg_tohost;
  wire[63:0] T969;
  wire[63:0] T776;
  wire[63:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire[63:0] T785;
  wire[63:0] T970;
  wire T786;
  reg  reg_stats;
  wire T971;
  wire T787;
  wire T788;
  wire T789;
  wire[63:0] T790;
  wire[63:0] T972;
  wire T791;
  wire[63:0] T792;
  wire[63:0] T973;
  wire T793;
  wire[63:0] T794;
  wire[63:0] T795;
  wire[63:0] T796;
  wire[63:0] T797;
  wire[63:0] T798;
  wire[63:0] T799;
  wire[63:0] T800;
  wire[23:0] T801;
  wire[23:0] T974;
  wire T802;
  wire[63:0] T803;
  wire[63:0] T804;
  wire[63:0] T805;
  wire[23:0] T806;
  wire[23:0] T975;
  wire T807;
  wire[63:0] T808;
  wire[63:0] T809;
  reg [63:0] reg_mscratch;
  wire[63:0] T810;
  wire T811;
  wire[63:0] T812;
  wire[63:0] T976;
  wire[7:0] T813;
  wire[7:0] T814;
  wire[7:0] T815;
  wire[3:0] T816;
  wire[1:0] T817;
  reg  reg_mie_usip;
  wire T977;
  wire[1:0] T818;
  reg  reg_mie_hsip;
  wire T978;
  wire[3:0] T819;
  wire[1:0] T820;
  reg  reg_mie_utip;
  wire T979;
  wire[1:0] T821;
  reg  reg_mie_htip;
  wire T980;
  wire[63:0] T822;
  wire[63:0] T981;
  wire[7:0] T823;
  wire[7:0] T824;
  wire[7:0] T825;
  wire[3:0] T826;
  wire[1:0] T827;
  reg  reg_mip_usip;
  wire T982;
  wire[1:0] T828;
  reg  reg_mip_hsip;
  wire T983;
  wire[3:0] T829;
  wire[1:0] T830;
  reg  reg_mip_utip;
  wire T984;
  wire[1:0] T831;
  reg  reg_mip_htip;
  wire T985;
  wire[63:0] T832;
  wire[63:0] T986;
  wire[8:0] T833;
  wire[63:0] T834;
  wire[63:0] T835;
  wire[63:0] T836;
  wire[63:0] T837;
  wire[63:0] T838;
  wire[63:0] T987;
  wire[63:0] T839;
  wire[63:0] T840;
  wire[63:0] T841;
  wire[63:0] T842;
  wire[63:0] T843;
  wire[63:0] T844;
  wire[63:0] T845;
  wire[63:0] T846;
  wire[63:0] T847;
  wire[63:0] T848;
  wire[63:0] T849;
  wire[63:0] T850;
  wire[63:0] T851;
  wire[63:0] T852;
  wire[63:0] T853;
  reg [5:0] R854;
  wire[5:0] T988;
  wire[5:0] T855;
  wire[5:0] T856;
  wire[5:0] T857;
  wire[6:0] T858;
  wire[6:0] T989;
  wire T859;
  wire[5:0] T860;
  wire T861;
  reg [57:0] R862;
  wire[57:0] T990;
  wire[57:0] T863;
  wire[57:0] T864;
  wire[57:0] T865;
  wire T866;
  wire T867;
  wire[57:0] T868;
  wire[63:0] T869;
  wire[63:0] T870;
  wire[63:0] T871;
  wire[63:0] T872;
  wire[63:0] T873;
  wire[63:0] T874;
  wire T991;
  wire T875;
  reg  host_pcr_rep_valid;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    reg_mstatus_prv = {1{$random}};
    reg_mstatus_prv1 = {1{$random}};
    reg_mstatus_prv2 = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    reg_mstatus_ie = {1{$random}};
    reg_mstatus_ie1 = {1{$random}};
    reg_mstatus_ie2 = {1{$random}};
    reg_mip_ssip = {1{$random}};
    reg_mie_ssip = {1{$random}};
    reg_mip_msip = {1{$random}};
    reg_mie_msip = {1{$random}};
    reg_mip_stip = {1{$random}};
    reg_mie_stip = {1{$random}};
    reg_mip_mtip = {1{$random}};
    reg_time = {2{$random}};
    reg_mtimecmp = {2{$random}};
    reg_mie_mtip = {1{$random}};
    reg_fromhost = {2{$random}};
    reg_frm = {1{$random}};
    R316 = {1{$random}};
    R319 = {2{$random}};
    reg_sepc = {2{$random}};
    reg_mepc = {2{$random}};
    reg_stvec = {2{$random}};
    reg_sptbr = {1{$random}};
    reg_mstatus_ie3 = {1{$random}};
    reg_mstatus_prv3 = {1{$random}};
    reg_mstatus_fs = {1{$random}};
    reg_mstatus_xs = {1{$random}};
    reg_mstatus_mprv = {1{$random}};
    reg_mstatus_vm = {1{$random}};
    reg_mstatus_zero1 = {1{$random}};
    reg_mstatus_sd_rv32 = {1{$random}};
    reg_mstatus_zero2 = {1{$random}};
    reg_wfi = {1{$random}};
    R424 = {1{$random}};
    R429 = {2{$random}};
    R437 = {1{$random}};
    R442 = {2{$random}};
    R450 = {1{$random}};
    R455 = {2{$random}};
    R463 = {1{$random}};
    R468 = {2{$random}};
    R476 = {1{$random}};
    R481 = {2{$random}};
    R489 = {1{$random}};
    R494 = {2{$random}};
    R502 = {1{$random}};
    R507 = {2{$random}};
    R515 = {1{$random}};
    R520 = {2{$random}};
    R528 = {1{$random}};
    R533 = {2{$random}};
    R541 = {1{$random}};
    R546 = {2{$random}};
    R554 = {1{$random}};
    R559 = {2{$random}};
    R567 = {1{$random}};
    R572 = {2{$random}};
    R580 = {1{$random}};
    R585 = {2{$random}};
    R593 = {1{$random}};
    R598 = {2{$random}};
    R606 = {1{$random}};
    R611 = {2{$random}};
    R619 = {1{$random}};
    R624 = {2{$random}};
    reg_sbadaddr = {2{$random}};
    reg_mbadaddr = {2{$random}};
    reg_scause = {2{$random}};
    reg_mcause = {2{$random}};
    reg_sscratch = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_mscratch = {2{$random}};
    reg_mie_usip = {1{$random}};
    reg_mie_hsip = {1{$random}};
    reg_mie_utip = {1{$random}};
    reg_mie_htip = {1{$random}};
    reg_mip_usip = {1{$random}};
    reg_mip_hsip = {1{$random}};
    reg_mip_utip = {1{$random}};
    reg_mip_htip = {1{$random}};
    R854 = {1{$random}};
    R862 = {2{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_data = {4{$random}};
//  assign io_rocc_dmem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_data = {4{$random}};
//  assign io_rocc_imem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
//  assign io_rocc_cmd_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 <= 4'h1;
  assign T3 = T885 + T4;
  assign T4 = {1'h0, T5};
  assign T5 = T884 + T6;
  assign T6 = {1'h0, T7};
  assign T7 = T882 + T8;
  assign T8 = {1'h0, io_csr_replay};
  assign T882 = {1'h0, csr_xcpt};
  assign csr_xcpt = T13 | insn_break;
  assign insn_break = T9 & system_insn;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T9 = T11 & T10;
  assign T10 = io_rw_addr[1'h0:1'h0];
  assign T11 = T12 ^ 1'h1;
  assign T12 = io_rw_addr[4'h8:4'h8];
  assign T13 = T19 | insn_call;
  assign insn_call = T14 & system_insn;
  assign T14 = T17 & T15;
  assign T15 = T16 ^ 1'h1;
  assign T16 = io_rw_addr[1'h0:1'h0];
  assign T17 = T18 ^ 1'h1;
  assign T18 = io_rw_addr[4'h8:4'h8];
  assign T19 = T96 | T20;
  assign T20 = system_insn & T21;
  assign T21 = priv_sufficient ^ 1'h1;
  assign priv_sufficient = csr_addr_priv <= reg_mstatus_prv;
  assign T22 = reset ? 2'h3 : T23;
  assign T23 = T90 ? T89 : T24;
  assign T24 = insn_redirect_trap ? 2'h1 : T25;
  assign T25 = insn_ret ? reg_mstatus_prv1 : T26;
  assign T26 = T27 ? 2'h3 : reg_mstatus_prv;
  assign T27 = io_exception | csr_xcpt;
  assign T28 = reset ? 2'h3 : T29;
  assign T29 = T78 ? T883 : T30;
  assign T30 = T71 ? T70 : T31;
  assign T31 = insn_ret ? reg_mstatus_prv2 : T32;
  assign T32 = T27 ? reg_mstatus_prv : reg_mstatus_prv1;
  assign T33 = reset ? 2'h0 : T34;
  assign T34 = T54 ? T37 : T35;
  assign T35 = insn_ret ? 2'h0 : T36;
  assign T36 = T27 ? reg_mstatus_prv1 : reg_mstatus_prv2;
  assign T37 = wdata[4'h8:3'h7];
  assign wdata = T53 ? io_rw_wdata : T38;
  assign T38 = T52 ? T50 : T39;
  assign T39 = T49 ? T48 : host_pcr_bits_data;
  assign T40 = host_pcr_req_fire ? io_rw_rdata : T41;
  assign T41 = T42 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T42 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T43;
  assign T43 = cpu_ren ^ 1'h1;
  assign cpu_ren = T45 & T44;
  assign T44 = system_insn ^ 1'h1;
  assign T45 = io_rw_cmd != 3'h0;
  assign T46 = host_pcr_req_fire ? 1'h0 : T47;
  assign T47 = T42 ? 1'h1 : host_pcr_req_valid;
  assign T48 = io_rw_rdata | io_rw_wdata;
  assign T49 = io_rw_cmd == 3'h2;
  assign T50 = io_rw_rdata & T51;
  assign T51 = ~ io_rw_wdata;
  assign T52 = io_rw_cmd == 3'h3;
  assign T53 = io_rw_cmd == 3'h1;
  assign T54 = T60 & T55;
  assign T55 = T57 | T56;
  assign T56 = 2'h1 == T37;
  assign T57 = T59 | T58;
  assign T58 = 2'h0 == T37;
  assign T59 = 2'h3 == T37;
  assign T60 = wen & T61;
  assign T61 = addr == 12'h300;
  assign addr = cpu_ren ? io_rw_addr : host_pcr_bits_addr;
  assign T62 = T42 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign wen = T65 | T63;
  assign T63 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T64 = T42 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T65 = cpu_wen & T66;
  assign T66 = read_only ^ 1'h1;
  assign read_only = T67 == 2'h3;
  assign T67 = io_rw_addr[4'hb:4'ha];
  assign cpu_wen = T68 & priv_sufficient;
  assign T68 = cpu_ren & T69;
  assign T69 = io_rw_cmd != 3'h5;
  assign T70 = wdata[3'h5:3'h4];
  assign T71 = T60 & T72;
  assign T72 = T74 | T73;
  assign T73 = 2'h1 == T70;
  assign T74 = T76 | T75;
  assign T75 = 2'h0 == T70;
  assign T76 = 2'h3 == T70;
  assign T883 = {1'h0, T77};
  assign T77 = wdata[3'h4:3'h4];
  assign T78 = wen & T79;
  assign T79 = addr == 12'h100;
  assign insn_ret = T80 & priv_sufficient;
  assign T80 = T81 & system_insn;
  assign T81 = T84 & T82;
  assign T82 = T83 ^ 1'h1;
  assign T83 = io_rw_addr[1'h0:1'h0];
  assign T84 = T87 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = io_rw_addr[1'h1:1'h1];
  assign T87 = io_rw_addr[4'h8:4'h8];
  assign insn_redirect_trap = maybe_insn_redirect_trap & priv_sufficient;
  assign maybe_insn_redirect_trap = T88 & system_insn;
  assign T88 = io_rw_addr[2'h2:2'h2];
  assign T89 = wdata[2'h2:1'h1];
  assign T90 = T60 & T91;
  assign T91 = T93 | T92;
  assign T92 = 2'h1 == T89;
  assign T93 = T95 | T94;
  assign T94 = 2'h0 == T89;
  assign T95 = 2'h3 == T89;
  assign csr_addr_priv = io_rw_addr[4'h9:4'h8];
  assign T96 = T214 | T97;
  assign T97 = cpu_ren & T98;
  assign T98 = T106 | T99;
  assign T99 = fp_csr & T100;
  assign T100 = T101 ^ 1'h1;
  assign T101 = io_status_fs != 2'h0;
  assign fp_csr = T103 | T102;
  assign T102 = addr == 12'h3;
  assign T103 = T105 | T104;
  assign T104 = addr == 12'h2;
  assign T105 = addr == 12'h1;
  assign T106 = T213 | T107;
  assign T107 = addr_valid ^ 1'h1;
  assign addr_valid = T109 | T108;
  assign T108 = addr == 12'hccf;
  assign T109 = T111 | T110;
  assign T110 = addr == 12'hcce;
  assign T111 = T113 | T112;
  assign T112 = addr == 12'hccd;
  assign T113 = T115 | T114;
  assign T114 = addr == 12'hccc;
  assign T115 = T117 | T116;
  assign T116 = addr == 12'hccb;
  assign T117 = T119 | T118;
  assign T118 = addr == 12'hcca;
  assign T119 = T121 | T120;
  assign T120 = addr == 12'hcc9;
  assign T121 = T123 | T122;
  assign T122 = addr == 12'hcc8;
  assign T123 = T125 | T124;
  assign T124 = addr == 12'hcc7;
  assign T125 = T127 | T126;
  assign T126 = addr == 12'hcc6;
  assign T127 = T129 | T128;
  assign T128 = addr == 12'hcc5;
  assign T129 = T131 | T130;
  assign T130 = addr == 12'hcc4;
  assign T131 = T133 | T132;
  assign T132 = addr == 12'hcc3;
  assign T133 = T135 | T134;
  assign T134 = addr == 12'hcc2;
  assign T135 = T137 | T136;
  assign T136 = addr == 12'hcc1;
  assign T137 = T139 | T138;
  assign T138 = addr == 12'hcc0;
  assign T139 = T141 | T140;
  assign T140 = addr == 12'h101;
  assign T141 = T143 | T142;
  assign T142 = addr == 12'h141;
  assign T143 = T145 | T144;
  assign T144 = addr == 12'h181;
  assign T145 = T147 | T146;
  assign T146 = addr == 12'h180;
  assign T147 = T149 | T148;
  assign T148 = addr == 12'hd43;
  assign T149 = T151 | T150;
  assign T150 = addr == 12'hd42;
  assign T151 = T153 | T152;
  assign T152 = addr == 12'h140;
  assign T153 = T155 | T154;
  assign T154 = addr == 12'h104;
  assign T155 = T157 | T156;
  assign T156 = addr == 12'h144;
  assign T157 = T158 | T79;
  assign T158 = T160 | T159;
  assign T159 = addr == 12'h781;
  assign T160 = T162 | T161;
  assign T161 = addr == 12'h780;
  assign T162 = T164 | T163;
  assign T163 = addr == 12'hc0;
  assign T164 = T166 | T165;
  assign T165 = addr == 12'h783;
  assign T166 = T168 | T167;
  assign T167 = addr == 12'hf10;
  assign T168 = T170 | T169;
  assign T169 = addr == 12'h321;
  assign T170 = T172 | T171;
  assign T171 = addr == 12'h342;
  assign T172 = T174 | T173;
  assign T173 = addr == 12'h343;
  assign T174 = T176 | T175;
  assign T175 = addr == 12'h341;
  assign T176 = T178 | T177;
  assign T177 = addr == 12'h340;
  assign T178 = T180 | T179;
  assign T179 = addr == 12'h304;
  assign T180 = T182 | T181;
  assign T181 = addr == 12'h344;
  assign T182 = T184 | T183;
  assign T183 = addr == 12'h301;
  assign T184 = T186 | T185;
  assign T185 = addr == 12'h782;
  assign T186 = T188 | T187;
  assign T187 = addr == 12'h302;
  assign T188 = T189 | T61;
  assign T189 = T191 | T190;
  assign T190 = addr == 12'hf01;
  assign T191 = T193 | T192;
  assign T192 = addr == 12'hf00;
  assign T193 = T195 | T194;
  assign T194 = addr == 12'h701;
  assign T195 = T197 | T196;
  assign T196 = addr == 12'ha01;
  assign T197 = T199 | T198;
  assign T198 = addr == 12'hd01;
  assign T199 = T201 | T200;
  assign T200 = addr == 12'h901;
  assign T201 = T203 | T202;
  assign T202 = addr == 12'hc01;
  assign T203 = T205 | T204;
  assign T204 = addr == 12'h902;
  assign T205 = T207 | T206;
  assign T206 = addr == 12'hc02;
  assign T207 = T209 | T208;
  assign T208 = addr == 12'h900;
  assign T209 = T211 | T210;
  assign T210 = addr == 12'hc00;
  assign T211 = T212 | T102;
  assign T212 = T105 | T104;
  assign T213 = priv_sufficient ^ 1'h1;
  assign T214 = cpu_wen & read_only;
  assign T884 = {2'h0, io_exception};
  assign T885 = {2'h0, T215};
  assign T215 = T886 + T216;
  assign T216 = {1'h0, insn_redirect_trap};
  assign T886 = {1'h0, insn_ret};
  assign io_interrupt_cause = T217;
  assign T217 = T297 ? 64'h8000000000000002 : T218;
  assign T218 = T282 ? 64'h8000000000000001 : T219;
  assign T219 = T270 ? 64'h8000000000000001 : T220;
  assign T220 = T259 ? 64'h8000000000000000 : T221;
  assign T221 = T222 ? 64'h8000000000000000 : 64'h0;
  assign T222 = T246 & T223;
  assign T223 = T245 | T224;
  assign T224 = T244 & reg_mstatus_ie;
  assign T225 = reset ? 1'h0 : T226;
  assign T226 = T78 ? T243 : T227;
  assign T227 = T60 ? T242 : T228;
  assign T228 = insn_ret ? reg_mstatus_ie1 : T229;
  assign T229 = T27 ? 1'h0 : reg_mstatus_ie;
  assign T230 = reset ? 1'h0 : T231;
  assign T231 = T78 ? T241 : T232;
  assign T232 = T60 ? T240 : T233;
  assign T233 = insn_ret ? reg_mstatus_ie2 : T234;
  assign T234 = T27 ? reg_mstatus_ie : reg_mstatus_ie1;
  assign T235 = reset ? 1'h0 : T236;
  assign T236 = T60 ? T239 : T237;
  assign T237 = insn_ret ? 1'h1 : T238;
  assign T238 = T27 ? reg_mstatus_ie1 : reg_mstatus_ie2;
  assign T239 = wdata[3'h6:3'h6];
  assign T240 = wdata[2'h3:2'h3];
  assign T241 = wdata[2'h3:2'h3];
  assign T242 = wdata[1'h0:1'h0];
  assign T243 = wdata[1'h0:1'h0];
  assign T244 = reg_mstatus_prv == 2'h1;
  assign T245 = reg_mstatus_prv < 2'h1;
  assign T246 = reg_mie_ssip & reg_mip_ssip;
  assign T887 = reset ? 1'h0 : T247;
  assign T247 = T252 ? T251 : T248;
  assign T248 = T250 ? T249 : reg_mip_ssip;
  assign T249 = wdata[1'h1:1'h1];
  assign T250 = wen & T181;
  assign T251 = wdata[1'h1:1'h1];
  assign T252 = wen & T156;
  assign T888 = reset ? 1'h0 : T253;
  assign T253 = T258 ? T257 : T254;
  assign T254 = T256 ? T255 : reg_mie_ssip;
  assign T255 = wdata[1'h1:1'h1];
  assign T256 = wen & T179;
  assign T257 = wdata[1'h1:1'h1];
  assign T258 = wen & T154;
  assign T259 = T264 & T260;
  assign T260 = T263 | T261;
  assign T261 = T262 & reg_mstatus_ie;
  assign T262 = reg_mstatus_prv == 2'h3;
  assign T263 = reg_mstatus_prv < 2'h3;
  assign T264 = reg_mie_msip & reg_mip_msip;
  assign T889 = reset ? 1'h0 : T265;
  assign T265 = io_host_ipi_rep_valid ? 1'h1 : T266;
  assign T266 = T250 ? T267 : reg_mip_msip;
  assign T267 = wdata[2'h3:2'h3];
  assign T890 = reset ? 1'h0 : T268;
  assign T268 = T256 ? T269 : reg_mie_msip;
  assign T269 = wdata[2'h3:2'h3];
  assign T270 = T275 & T271;
  assign T271 = T274 | T272;
  assign T272 = T273 & reg_mstatus_ie;
  assign T273 = reg_mstatus_prv == 2'h1;
  assign T274 = reg_mstatus_prv < 2'h1;
  assign T275 = reg_mie_stip & reg_mip_stip;
  assign T891 = reset ? 1'h0 : T276;
  assign T276 = T250 ? T277 : reg_mip_stip;
  assign T277 = wdata[3'h5:3'h5];
  assign T892 = reset ? 1'h0 : T278;
  assign T278 = T258 ? T281 : T279;
  assign T279 = T256 ? T280 : reg_mie_stip;
  assign T280 = wdata[3'h5:3'h5];
  assign T281 = wdata[3'h5:3'h5];
  assign T282 = T287 & T283;
  assign T283 = T286 | T284;
  assign T284 = T285 & reg_mstatus_ie;
  assign T285 = reg_mstatus_prv == 2'h3;
  assign T286 = reg_mstatus_prv < 2'h3;
  assign T287 = reg_mie_mtip & reg_mip_mtip;
  assign T893 = reset ? 1'h0 : T288;
  assign T288 = T294 ? 1'h0 : T289;
  assign T289 = T290 ? 1'h1 : reg_mip_mtip;
  assign T290 = reg_mtimecmp <= reg_time;
  assign T291 = T292 ? wdata : reg_time;
  assign T292 = wen & T185;
  assign T293 = T294 ? wdata : reg_mtimecmp;
  assign T294 = wen & T169;
  assign T894 = reset ? 1'h0 : T295;
  assign T295 = T256 ? T296 : reg_mie_mtip;
  assign T296 = wdata[3'h7:3'h7];
  assign T297 = T302 & T298;
  assign T298 = T301 | T299;
  assign T299 = T300 & reg_mstatus_ie;
  assign T300 = reg_mstatus_prv == 2'h3;
  assign T301 = reg_mstatus_prv < 2'h3;
  assign T302 = reg_fromhost != 64'h0;
  assign T895 = reset ? 64'h0 : T303;
  assign T303 = T304 ? wdata : reg_fromhost;
  assign T304 = T308 & T305;
  assign T305 = T307 | T306;
  assign T306 = host_pcr_req_fire ^ 1'h1;
  assign T307 = reg_fromhost == 64'h0;
  assign T308 = wen & T159;
  assign io_interrupt = T309;
  assign T309 = io_interrupt_cause[6'h3f:6'h3f];
  assign io_fcsr_rm = reg_frm;
  assign T896 = T310[2'h2:1'h0];
  assign T310 = T314 ? T898 : T311;
  assign T311 = T312 ? wdata : T897;
  assign T897 = {61'h0, reg_frm};
  assign T312 = wen & T104;
  assign T898 = {5'h0, T313};
  assign T313 = wdata >> 3'h5;
  assign T314 = wen & T102;
  assign io_time = T315;
  assign T315 = {R319, R316};
  assign T899 = reset ? 6'h0 : T317;
  assign T317 = T318[3'h5:1'h0];
  assign T318 = T900 + 7'h1;
  assign T900 = {1'h0, R316};
  assign T901 = reset ? 58'h0 : T320;
  assign T320 = T322 ? T321 : R319;
  assign T321 = R319 + 58'h1;
  assign T322 = T318[3'h6:3'h6];
  assign io_fatc = insn_sfence_vm;
  assign insn_sfence_vm = T323 & priv_sufficient;
  assign T323 = T324 & system_insn;
  assign T324 = T326 & T325;
  assign T325 = io_rw_addr[1'h0:1'h0];
  assign T326 = T329 & T327;
  assign T327 = T328 ^ 1'h1;
  assign T328 = io_rw_addr[1'h1:1'h1];
  assign T329 = io_rw_addr[4'h8:4'h8];
  assign io_evec = T330;
  assign T330 = T358 ? T908 : T331;
  assign T331 = maybe_insn_redirect_trap ? T349 : T332;
  assign T332 = T348 ? reg_mepc : reg_sepc;
  assign T902 = T333[6'h27:1'h0];
  assign T333 = T338 ? T335 : T903;
  assign T903 = {24'h0, T334};
  assign T334 = insn_redirect_trap ? reg_mepc : reg_sepc;
  assign T335 = ~ T336;
  assign T336 = T337 | 64'h3;
  assign T337 = ~ wdata;
  assign T338 = wen & T142;
  assign T904 = T339[6'h27:1'h0];
  assign T339 = T347 ? T344 : T905;
  assign T905 = {24'h0, T340};
  assign T340 = T27 ? T341 : reg_mepc;
  assign T341 = ~ T342;
  assign T342 = T343 | 40'h3;
  assign T343 = ~ io_pc;
  assign T344 = ~ T345;
  assign T345 = T346 | 64'h3;
  assign T346 = ~ wdata;
  assign T347 = wen & T175;
  assign T348 = reg_mstatus_prv[1'h1:1'h1];
  assign T349 = {T355, reg_stvec};
  assign T906 = T350[6'h26:1'h0];
  assign T350 = T354 ? T351 : T907;
  assign T907 = {25'h0, reg_stvec};
  assign T351 = ~ T352;
  assign T352 = T353 | 64'h3;
  assign T353 = ~ wdata;
  assign T354 = wen & T140;
  assign T355 = reg_stvec[6'h26:6'h26];
  assign T908 = {31'h0, T356};
  assign T356 = T909 + 9'h100;
  assign T909 = {1'h0, T357};
  assign T357 = reg_mstatus_prv << 3'h6;
  assign T358 = io_exception | csr_xcpt;
  assign io_ptbr = reg_sptbr;
  assign T359 = T362 ? T360 : reg_sptbr;
  assign T360 = {T361, 12'h0};
  assign T361 = wdata[5'h1f:4'hc];
  assign T362 = wen & T146;
  assign io_status_ie = reg_mstatus_ie;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_ie1 = reg_mstatus_ie1;
  assign io_status_prv1 = reg_mstatus_prv1;
  assign io_status_ie2 = reg_mstatus_ie2;
  assign io_status_prv2 = reg_mstatus_prv2;
  assign io_status_ie3 = reg_mstatus_ie3;
  assign T363 = reset ? 1'h0 : reg_mstatus_ie3;
  assign io_status_prv3 = reg_mstatus_prv3;
  assign T364 = reset ? 2'h0 : reg_mstatus_prv3;
  assign io_status_fs = T365;
  assign T365 = 2'h0 - T910;
  assign T910 = {1'h0, T366};
  assign T366 = reg_mstatus_fs != 2'h0;
  assign T367 = reset ? 2'h0 : T368;
  assign T368 = T78 ? T371 : T369;
  assign T369 = T60 ? T370 : reg_mstatus_fs;
  assign T370 = wdata[4'hd:4'hc];
  assign T371 = wdata[4'hd:4'hc];
  assign io_status_xs = T372;
  assign T372 = 2'h0 - T911;
  assign T911 = {1'h0, T373};
  assign T373 = reg_mstatus_xs != 2'h0;
  assign T374 = reset ? 2'h0 : reg_mstatus_xs;
  assign io_status_mprv = reg_mstatus_mprv;
  assign T375 = reset ? 1'h0 : T376;
  assign T376 = T78 ? T380 : T377;
  assign T377 = T60 ? T379 : T378;
  assign T378 = T27 ? 1'h0 : reg_mstatus_mprv;
  assign T379 = wdata[5'h10:5'h10];
  assign T380 = wdata[5'h10:5'h10];
  assign io_status_vm = reg_mstatus_vm;
  assign T381 = reset ? 5'h0 : T382;
  assign T382 = T387 ? 5'h9 : T383;
  assign T383 = T384 ? 5'h0 : reg_mstatus_vm;
  assign T384 = T60 & T385;
  assign T385 = T386 == 5'h0;
  assign T386 = wdata[5'h15:5'h11];
  assign T387 = T60 & T388;
  assign T388 = T386 == 5'h9;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign T389 = reset ? 9'h0 : reg_mstatus_zero1;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign T390 = reset ? 1'h0 : reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign T391 = reset ? 31'h0 : reg_mstatus_zero2;
  assign io_status_sd = T392;
  assign T392 = T394 | T393;
  assign T393 = io_status_xs == 2'h3;
  assign T394 = io_status_fs == 2'h3;
  assign io_eret = T395;
  assign T395 = insn_ret | insn_redirect_trap;
  assign io_csr_xcpt = csr_xcpt;
  assign io_csr_stall = reg_wfi;
  assign T912 = reset ? 1'h0 : T396;
  assign T396 = some_interrupt_pending ? 1'h0 : T397;
  assign T397 = insn_wfi ? 1'h1 : reg_wfi;
  assign insn_wfi = T398 & priv_sufficient;
  assign T398 = T399 & system_insn;
  assign T399 = T402 & T400;
  assign T400 = T401 ^ 1'h1;
  assign T401 = io_rw_addr[1'h0:1'h0];
  assign T402 = T404 & T403;
  assign T403 = io_rw_addr[1'h1:1'h1];
  assign T404 = io_rw_addr[4'h8:4'h8];
  assign some_interrupt_pending = T405;
  assign T405 = T417 ? 1'h1 : T406;
  assign T406 = T415 ? 1'h1 : T407;
  assign T407 = T413 ? 1'h1 : T408;
  assign T408 = T411 ? 1'h1 : T409;
  assign T409 = T246 & T410;
  assign T410 = reg_mstatus_prv <= 2'h1;
  assign T411 = T264 & T412;
  assign T412 = reg_mstatus_prv <= 2'h3;
  assign T413 = T275 & T414;
  assign T414 = reg_mstatus_prv <= 2'h1;
  assign T415 = T287 & T416;
  assign T416 = reg_mstatus_prv <= 2'h3;
  assign T417 = T302 & T418;
  assign T418 = reg_mstatus_prv <= 2'h3;
  assign io_csr_replay = T419;
  assign T419 = io_host_ipi_req_valid & T420;
  assign T420 = io_host_ipi_req_ready ^ 1'h1;
  assign io_rw_rdata = T421;
  assign T421 = T434 | T422;
  assign T422 = T108 ? T423 : 64'h0;
  assign T423 = {R429, R424};
  assign T913 = reset ? 6'h0 : T425;
  assign T425 = T428 ? T426 : R424;
  assign T426 = T427[3'h5:1'h0];
  assign T427 = T914 + 7'h1;
  assign T914 = {1'h0, R424};
  assign T428 = io_uarch_counters_15 != 1'h0;
  assign T915 = reset ? 58'h0 : T430;
  assign T430 = T432 ? T431 : R429;
  assign T431 = R429 + 58'h1;
  assign T432 = T428 & T433;
  assign T433 = T427[3'h6:3'h6];
  assign T434 = T447 | T435;
  assign T435 = T110 ? T436 : 64'h0;
  assign T436 = {R442, R437};
  assign T916 = reset ? 6'h0 : T438;
  assign T438 = T441 ? T439 : R437;
  assign T439 = T440[3'h5:1'h0];
  assign T440 = T917 + 7'h1;
  assign T917 = {1'h0, R437};
  assign T441 = io_uarch_counters_14 != 1'h0;
  assign T918 = reset ? 58'h0 : T443;
  assign T443 = T445 ? T444 : R442;
  assign T444 = R442 + 58'h1;
  assign T445 = T441 & T446;
  assign T446 = T440[3'h6:3'h6];
  assign T447 = T460 | T448;
  assign T448 = T112 ? T449 : 64'h0;
  assign T449 = {R455, R450};
  assign T919 = reset ? 6'h0 : T451;
  assign T451 = T454 ? T452 : R450;
  assign T452 = T453[3'h5:1'h0];
  assign T453 = T920 + 7'h1;
  assign T920 = {1'h0, R450};
  assign T454 = io_uarch_counters_13 != 1'h0;
  assign T921 = reset ? 58'h0 : T456;
  assign T456 = T458 ? T457 : R455;
  assign T457 = R455 + 58'h1;
  assign T458 = T454 & T459;
  assign T459 = T453[3'h6:3'h6];
  assign T460 = T473 | T461;
  assign T461 = T114 ? T462 : 64'h0;
  assign T462 = {R468, R463};
  assign T922 = reset ? 6'h0 : T464;
  assign T464 = T467 ? T465 : R463;
  assign T465 = T466[3'h5:1'h0];
  assign T466 = T923 + 7'h1;
  assign T923 = {1'h0, R463};
  assign T467 = io_uarch_counters_12 != 1'h0;
  assign T924 = reset ? 58'h0 : T469;
  assign T469 = T471 ? T470 : R468;
  assign T470 = R468 + 58'h1;
  assign T471 = T467 & T472;
  assign T472 = T466[3'h6:3'h6];
  assign T473 = T486 | T474;
  assign T474 = T116 ? T475 : 64'h0;
  assign T475 = {R481, R476};
  assign T925 = reset ? 6'h0 : T477;
  assign T477 = T480 ? T478 : R476;
  assign T478 = T479[3'h5:1'h0];
  assign T479 = T926 + 7'h1;
  assign T926 = {1'h0, R476};
  assign T480 = io_uarch_counters_11 != 1'h0;
  assign T927 = reset ? 58'h0 : T482;
  assign T482 = T484 ? T483 : R481;
  assign T483 = R481 + 58'h1;
  assign T484 = T480 & T485;
  assign T485 = T479[3'h6:3'h6];
  assign T486 = T499 | T487;
  assign T487 = T118 ? T488 : 64'h0;
  assign T488 = {R494, R489};
  assign T928 = reset ? 6'h0 : T490;
  assign T490 = T493 ? T491 : R489;
  assign T491 = T492[3'h5:1'h0];
  assign T492 = T929 + 7'h1;
  assign T929 = {1'h0, R489};
  assign T493 = io_uarch_counters_10 != 1'h0;
  assign T930 = reset ? 58'h0 : T495;
  assign T495 = T497 ? T496 : R494;
  assign T496 = R494 + 58'h1;
  assign T497 = T493 & T498;
  assign T498 = T492[3'h6:3'h6];
  assign T499 = T512 | T500;
  assign T500 = T120 ? T501 : 64'h0;
  assign T501 = {R507, R502};
  assign T931 = reset ? 6'h0 : T503;
  assign T503 = T506 ? T504 : R502;
  assign T504 = T505[3'h5:1'h0];
  assign T505 = T932 + 7'h1;
  assign T932 = {1'h0, R502};
  assign T506 = io_uarch_counters_9 != 1'h0;
  assign T933 = reset ? 58'h0 : T508;
  assign T508 = T510 ? T509 : R507;
  assign T509 = R507 + 58'h1;
  assign T510 = T506 & T511;
  assign T511 = T505[3'h6:3'h6];
  assign T512 = T525 | T513;
  assign T513 = T122 ? T514 : 64'h0;
  assign T514 = {R520, R515};
  assign T934 = reset ? 6'h0 : T516;
  assign T516 = T519 ? T517 : R515;
  assign T517 = T518[3'h5:1'h0];
  assign T518 = T935 + 7'h1;
  assign T935 = {1'h0, R515};
  assign T519 = io_uarch_counters_8 != 1'h0;
  assign T936 = reset ? 58'h0 : T521;
  assign T521 = T523 ? T522 : R520;
  assign T522 = R520 + 58'h1;
  assign T523 = T519 & T524;
  assign T524 = T518[3'h6:3'h6];
  assign T525 = T538 | T526;
  assign T526 = T124 ? T527 : 64'h0;
  assign T527 = {R533, R528};
  assign T937 = reset ? 6'h0 : T529;
  assign T529 = T532 ? T530 : R528;
  assign T530 = T531[3'h5:1'h0];
  assign T531 = T938 + 7'h1;
  assign T938 = {1'h0, R528};
  assign T532 = io_uarch_counters_7 != 1'h0;
  assign T939 = reset ? 58'h0 : T534;
  assign T534 = T536 ? T535 : R533;
  assign T535 = R533 + 58'h1;
  assign T536 = T532 & T537;
  assign T537 = T531[3'h6:3'h6];
  assign T538 = T551 | T539;
  assign T539 = T126 ? T540 : 64'h0;
  assign T540 = {R546, R541};
  assign T940 = reset ? 6'h0 : T542;
  assign T542 = T545 ? T543 : R541;
  assign T543 = T544[3'h5:1'h0];
  assign T544 = T941 + 7'h1;
  assign T941 = {1'h0, R541};
  assign T545 = io_uarch_counters_6 != 1'h0;
  assign T942 = reset ? 58'h0 : T547;
  assign T547 = T549 ? T548 : R546;
  assign T548 = R546 + 58'h1;
  assign T549 = T545 & T550;
  assign T550 = T544[3'h6:3'h6];
  assign T551 = T564 | T552;
  assign T552 = T128 ? T553 : 64'h0;
  assign T553 = {R559, R554};
  assign T943 = reset ? 6'h0 : T555;
  assign T555 = T558 ? T556 : R554;
  assign T556 = T557[3'h5:1'h0];
  assign T557 = T944 + 7'h1;
  assign T944 = {1'h0, R554};
  assign T558 = io_uarch_counters_5 != 1'h0;
  assign T945 = reset ? 58'h0 : T560;
  assign T560 = T562 ? T561 : R559;
  assign T561 = R559 + 58'h1;
  assign T562 = T558 & T563;
  assign T563 = T557[3'h6:3'h6];
  assign T564 = T577 | T565;
  assign T565 = T130 ? T566 : 64'h0;
  assign T566 = {R572, R567};
  assign T946 = reset ? 6'h0 : T568;
  assign T568 = T571 ? T569 : R567;
  assign T569 = T570[3'h5:1'h0];
  assign T570 = T947 + 7'h1;
  assign T947 = {1'h0, R567};
  assign T571 = io_uarch_counters_4 != 1'h0;
  assign T948 = reset ? 58'h0 : T573;
  assign T573 = T575 ? T574 : R572;
  assign T574 = R572 + 58'h1;
  assign T575 = T571 & T576;
  assign T576 = T570[3'h6:3'h6];
  assign T577 = T590 | T578;
  assign T578 = T132 ? T579 : 64'h0;
  assign T579 = {R585, R580};
  assign T949 = reset ? 6'h0 : T581;
  assign T581 = T584 ? T582 : R580;
  assign T582 = T583[3'h5:1'h0];
  assign T583 = T950 + 7'h1;
  assign T950 = {1'h0, R580};
  assign T584 = io_uarch_counters_3 != 1'h0;
  assign T951 = reset ? 58'h0 : T586;
  assign T586 = T588 ? T587 : R585;
  assign T587 = R585 + 58'h1;
  assign T588 = T584 & T589;
  assign T589 = T583[3'h6:3'h6];
  assign T590 = T603 | T591;
  assign T591 = T134 ? T592 : 64'h0;
  assign T592 = {R598, R593};
  assign T952 = reset ? 6'h0 : T594;
  assign T594 = T597 ? T595 : R593;
  assign T595 = T596[3'h5:1'h0];
  assign T596 = T953 + 7'h1;
  assign T953 = {1'h0, R593};
  assign T597 = io_uarch_counters_2 != 1'h0;
  assign T954 = reset ? 58'h0 : T599;
  assign T599 = T601 ? T600 : R598;
  assign T600 = R598 + 58'h1;
  assign T601 = T597 & T602;
  assign T602 = T596[3'h6:3'h6];
  assign T603 = T616 | T604;
  assign T604 = T136 ? T605 : 64'h0;
  assign T605 = {R611, R606};
  assign T955 = reset ? 6'h0 : T607;
  assign T607 = T610 ? T608 : R606;
  assign T608 = T609[3'h5:1'h0];
  assign T609 = T956 + 7'h1;
  assign T956 = {1'h0, R606};
  assign T610 = io_uarch_counters_1 != 1'h0;
  assign T957 = reset ? 58'h0 : T612;
  assign T612 = T614 ? T613 : R611;
  assign T613 = R611 + 58'h1;
  assign T614 = T610 & T615;
  assign T615 = T609[3'h6:3'h6];
  assign T616 = T629 | T617;
  assign T617 = T138 ? T618 : 64'h0;
  assign T618 = {R624, R619};
  assign T958 = reset ? 6'h0 : T620;
  assign T620 = T623 ? T621 : R619;
  assign T621 = T622[3'h5:1'h0];
  assign T622 = T959 + 7'h1;
  assign T959 = {1'h0, R619};
  assign T623 = io_uarch_counters_0 != 1'h0;
  assign T960 = reset ? 58'h0 : T625;
  assign T625 = T627 ? T626 : R624;
  assign T626 = R624 + 58'h1;
  assign T627 = T623 & T628;
  assign T628 = T622[3'h6:3'h6];
  assign T629 = T634 | T630;
  assign T630 = T140 ? T631 : 64'h0;
  assign T631 = {T632, reg_stvec};
  assign T632 = 25'h0 - T961;
  assign T961 = {24'h0, T633};
  assign T633 = reg_stvec[6'h26:6'h26];
  assign T634 = T639 | T635;
  assign T635 = T142 ? T636 : 64'h0;
  assign T636 = {T637, reg_sepc};
  assign T637 = 24'h0 - T962;
  assign T962 = {23'h0, T638};
  assign T638 = reg_sepc[6'h27:6'h27];
  assign T639 = T640 | 64'h0;
  assign T640 = T642 | T963;
  assign T963 = {32'h0, T641};
  assign T641 = T146 ? reg_sptbr : 32'h0;
  assign T642 = T669 | T643;
  assign T643 = T148 ? T644 : 64'h0;
  assign T644 = {T667, reg_sbadaddr};
  assign T645 = insn_redirect_trap ? reg_mbadaddr : reg_sbadaddr;
  assign T646 = T666 ? T665 : T647;
  assign T647 = T657 ? T649 : T648;
  assign T648 = T27 ? io_pc : reg_mbadaddr;
  assign T649 = {T651, T650};
  assign T650 = io_rw_wdata[6'h26:1'h0];
  assign T651 = T655 ? T654 : T652;
  assign T652 = T653 != 25'h0;
  assign T653 = io_rw_wdata[6'h3f:6'h27];
  assign T654 = T653 == 25'h1ffffff;
  assign T655 = $signed(T656) < $signed(1'h0);
  assign T656 = T650;
  assign T657 = T27 & T658;
  assign T658 = T660 | T659;
  assign T659 = io_cause == 64'h6;
  assign T660 = T662 | T661;
  assign T661 = io_cause == 64'h7;
  assign T662 = T664 | T663;
  assign T663 = io_cause == 64'h4;
  assign T664 = io_cause == 64'h5;
  assign T665 = wdata[6'h27:1'h0];
  assign T666 = wen & T173;
  assign T667 = 24'h0 - T964;
  assign T964 = {23'h0, T668};
  assign T668 = reg_sbadaddr[6'h27:6'h27];
  assign T669 = T683 | T670;
  assign T670 = T150 ? reg_scause : 64'h0;
  assign T671 = insn_redirect_trap ? reg_mcause : reg_scause;
  assign T672 = T682 ? T681 : T673;
  assign T673 = T680 ? T965 : T674;
  assign T674 = T678 ? 64'h3 : T675;
  assign T675 = T677 ? 64'h2 : T676;
  assign T676 = T27 ? io_cause : reg_mcause;
  assign T677 = T27 & csr_xcpt;
  assign T678 = T677 & insn_break;
  assign T965 = {60'h0, T679};
  assign T679 = T966 + 4'h8;
  assign T966 = {2'h0, reg_mstatus_prv};
  assign T680 = T677 & insn_call;
  assign T681 = wdata & 64'h800000000000001f;
  assign T682 = wen & T171;
  assign T683 = T687 | T684;
  assign T684 = T152 ? reg_sscratch : 64'h0;
  assign T685 = T686 ? wdata : reg_sscratch;
  assign T686 = wen & T152;
  assign T687 = T705 | T967;
  assign T967 = {56'h0, T688};
  assign T688 = T154 ? T689 : 8'h0;
  assign T689 = T690;
  assign T690 = {T698, T691};
  assign T691 = {T695, T692};
  assign T692 = {T694, T693};
  assign T693 = 1'h0;
  assign T694 = reg_mie_ssip;
  assign T695 = {T697, T696};
  assign T696 = 1'h0;
  assign T697 = 1'h0;
  assign T698 = {T702, T699};
  assign T699 = {T701, T700};
  assign T700 = 1'h0;
  assign T701 = reg_mie_stip;
  assign T702 = {T704, T703};
  assign T703 = 1'h0;
  assign T704 = 1'h0;
  assign T705 = T723 | T968;
  assign T968 = {56'h0, T706};
  assign T706 = T156 ? T707 : 8'h0;
  assign T707 = T708;
  assign T708 = {T716, T709};
  assign T709 = {T713, T710};
  assign T710 = {T712, T711};
  assign T711 = 1'h0;
  assign T712 = reg_mip_ssip;
  assign T713 = {T715, T714};
  assign T714 = 1'h0;
  assign T715 = 1'h0;
  assign T716 = {T720, T717};
  assign T717 = {T719, T718};
  assign T718 = 1'h0;
  assign T719 = reg_mip_stip;
  assign T720 = {T722, T721};
  assign T721 = 1'h0;
  assign T722 = 1'h0;
  assign T723 = T772 | T724;
  assign T724 = T79 ? T725 : 64'h0;
  assign T725 = T726;
  assign T726 = {T757, T727};
  assign T727 = {T750, T728};
  assign T728 = {T748, T729};
  assign T729 = {T747, T730};
  assign T730 = T731;
  assign T731 = read_mstatus[1'h0:1'h0];
  assign read_mstatus = T732;
  assign T732 = {T740, T733};
  assign T733 = {T737, T734};
  assign T734 = {T736, T735};
  assign T735 = {io_status_prv, io_status_ie};
  assign T736 = {io_status_prv1, io_status_ie1};
  assign T737 = {T739, T738};
  assign T738 = {io_status_prv2, io_status_ie2};
  assign T739 = {io_status_prv3, io_status_ie3};
  assign T740 = {T744, T741};
  assign T741 = {T743, T742};
  assign T742 = {io_status_xs, io_status_fs};
  assign T743 = {io_status_vm, io_status_mprv};
  assign T744 = {T746, T745};
  assign T745 = {io_status_sd_rv32, io_status_zero1};
  assign T746 = {io_status_sd, io_status_zero2};
  assign T747 = 2'h0;
  assign T748 = T749;
  assign T749 = read_mstatus[2'h3:2'h3];
  assign T750 = {T755, T751};
  assign T751 = {T754, T752};
  assign T752 = T753;
  assign T753 = read_mstatus[3'h4:3'h4];
  assign T754 = 7'h0;
  assign T755 = T756;
  assign T756 = read_mstatus[4'hd:4'hc];
  assign T757 = {T765, T758};
  assign T758 = {T764, T759};
  assign T759 = {T762, T760};
  assign T760 = T761;
  assign T761 = read_mstatus[4'hf:4'he];
  assign T762 = T763;
  assign T763 = read_mstatus[5'h10:5'h10];
  assign T764 = 14'h0;
  assign T765 = {T770, T766};
  assign T766 = {T769, T767};
  assign T767 = T768;
  assign T768 = read_mstatus[5'h1f:5'h1f];
  assign T769 = 31'h0;
  assign T770 = T771;
  assign T771 = read_mstatus[6'h3f:6'h3f];
  assign T772 = T774 | T773;
  assign T773 = T159 ? reg_fromhost : 64'h0;
  assign T774 = T785 | T775;
  assign T775 = T161 ? reg_tohost : 64'h0;
  assign T969 = reset ? 64'h0 : T776;
  assign T776 = T781 ? wdata : T777;
  assign T777 = T778 ? 64'h0 : reg_tohost;
  assign T778 = T779 & T161;
  assign T779 = host_pcr_req_fire & T780;
  assign T780 = host_pcr_bits_rw ^ 1'h1;
  assign T781 = T784 & T782;
  assign T782 = T783 | host_pcr_req_fire;
  assign T783 = reg_tohost == 64'h0;
  assign T784 = wen & T161;
  assign T785 = T790 | T970;
  assign T970 = {63'h0, T786};
  assign T786 = T163 ? reg_stats : 1'h0;
  assign T971 = reset ? 1'h0 : T787;
  assign T787 = T789 ? T788 : reg_stats;
  assign T788 = wdata[1'h0:1'h0];
  assign T789 = wen & T163;
  assign T790 = T792 | T972;
  assign T972 = {63'h0, T791};
  assign T791 = T165 ? io_host_id : 1'h0;
  assign T792 = T794 | T973;
  assign T973 = {63'h0, T793};
  assign T793 = T167 ? io_host_id : 1'h0;
  assign T794 = T796 | T795;
  assign T795 = T169 ? reg_mtimecmp : 64'h0;
  assign T796 = T798 | T797;
  assign T797 = T171 ? reg_mcause : 64'h0;
  assign T798 = T803 | T799;
  assign T799 = T173 ? T800 : 64'h0;
  assign T800 = {T801, reg_mbadaddr};
  assign T801 = 24'h0 - T974;
  assign T974 = {23'h0, T802};
  assign T802 = reg_mbadaddr[6'h27:6'h27];
  assign T803 = T808 | T804;
  assign T804 = T175 ? T805 : 64'h0;
  assign T805 = {T806, reg_mepc};
  assign T806 = 24'h0 - T975;
  assign T975 = {23'h0, T807};
  assign T807 = reg_mepc[6'h27:6'h27];
  assign T808 = T812 | T809;
  assign T809 = T177 ? reg_mscratch : 64'h0;
  assign T810 = T811 ? wdata : reg_mscratch;
  assign T811 = wen & T177;
  assign T812 = T822 | T976;
  assign T976 = {56'h0, T813};
  assign T813 = T179 ? T814 : 8'h0;
  assign T814 = T815;
  assign T815 = {T819, T816};
  assign T816 = {T818, T817};
  assign T817 = {reg_mie_ssip, reg_mie_usip};
  assign T977 = reset ? 1'h0 : reg_mie_usip;
  assign T818 = {reg_mie_msip, reg_mie_hsip};
  assign T978 = reset ? 1'h0 : reg_mie_hsip;
  assign T819 = {T821, T820};
  assign T820 = {reg_mie_stip, reg_mie_utip};
  assign T979 = reset ? 1'h0 : reg_mie_utip;
  assign T821 = {reg_mie_mtip, reg_mie_htip};
  assign T980 = reset ? 1'h0 : reg_mie_htip;
  assign T822 = T832 | T981;
  assign T981 = {56'h0, T823};
  assign T823 = T181 ? T824 : 8'h0;
  assign T824 = T825;
  assign T825 = {T829, T826};
  assign T826 = {T828, T827};
  assign T827 = {reg_mip_ssip, reg_mip_usip};
  assign T982 = reset ? 1'h0 : reg_mip_usip;
  assign T828 = {reg_mip_msip, reg_mip_hsip};
  assign T983 = reset ? 1'h0 : reg_mip_hsip;
  assign T829 = {T831, T830};
  assign T830 = {reg_mip_stip, reg_mip_utip};
  assign T984 = reset ? 1'h0 : reg_mip_utip;
  assign T831 = {reg_mip_mtip, reg_mip_htip};
  assign T985 = reset ? 1'h0 : reg_mip_htip;
  assign T832 = T834 | T986;
  assign T986 = {55'h0, T833};
  assign T833 = T183 ? 9'h100 : 9'h0;
  assign T834 = T835 | 64'h0;
  assign T835 = T836 | 64'h0;
  assign T836 = T838 | T837;
  assign T837 = T61 ? read_mstatus : 64'h0;
  assign T838 = T839 | T987;
  assign T987 = {63'h0, T190};
  assign T839 = T841 | T840;
  assign T840 = T192 ? 64'h8000000000041101 : 64'h0;
  assign T841 = T843 | T842;
  assign T842 = T194 ? reg_time : 64'h0;
  assign T843 = T845 | T844;
  assign T844 = T196 ? reg_time : 64'h0;
  assign T845 = T847 | T846;
  assign T846 = T198 ? reg_time : 64'h0;
  assign T847 = T849 | T848;
  assign T848 = T200 ? reg_time : 64'h0;
  assign T849 = T851 | T850;
  assign T850 = T202 ? reg_time : 64'h0;
  assign T851 = T869 | T852;
  assign T852 = T204 ? T853 : 64'h0;
  assign T853 = {R862, R854};
  assign T988 = reset ? 6'h0 : T855;
  assign T855 = T861 ? T860 : T856;
  assign T856 = T859 ? T857 : R854;
  assign T857 = T858[3'h5:1'h0];
  assign T858 = T989 + 7'h1;
  assign T989 = {1'h0, R854};
  assign T859 = io_retire != 1'h0;
  assign T860 = wdata[3'h5:1'h0];
  assign T861 = wen & T204;
  assign T990 = reset ? 58'h0 : T863;
  assign T863 = T861 ? T868 : T864;
  assign T864 = T866 ? T865 : R862;
  assign T865 = R862 + 58'h1;
  assign T866 = T859 & T867;
  assign T867 = T858[3'h6:3'h6];
  assign T868 = wdata[6'h3f:3'h6];
  assign T869 = T871 | T870;
  assign T870 = T206 ? T853 : 64'h0;
  assign T871 = T873 | T872;
  assign T872 = T208 ? T315 : 64'h0;
  assign T873 = 64'h0 | T874;
  assign T874 = T210 ? T315 : 64'h0;
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T991;
  assign T991 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T875;
  assign T875 = cpu_wen & T165;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T876 = T878 ? 1'h0 : T877;
  assign T877 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T878 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T879;
  assign T879 = T881 & T880;
  assign T880 = host_pcr_rep_valid ^ 1'h1;
  assign T881 = host_pcr_req_valid ^ 1'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "these conditions must be mutually exclusive");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if(T90) begin
      reg_mstatus_prv <= T89;
    end else if(insn_redirect_trap) begin
      reg_mstatus_prv <= 2'h1;
    end else if(insn_ret) begin
      reg_mstatus_prv <= reg_mstatus_prv1;
    end else if(T27) begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_prv1 <= 2'h3;
    end else if(T78) begin
      reg_mstatus_prv1 <= T883;
    end else if(T71) begin
      reg_mstatus_prv1 <= T70;
    end else if(insn_ret) begin
      reg_mstatus_prv1 <= reg_mstatus_prv2;
    end else if(T27) begin
      reg_mstatus_prv1 <= reg_mstatus_prv;
    end
    if(reset) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T54) begin
      reg_mstatus_prv2 <= T37;
    end else if(insn_ret) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T27) begin
      reg_mstatus_prv2 <= reg_mstatus_prv1;
    end
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T42) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T42) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T42) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T42) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(reset) begin
      reg_mstatus_ie <= 1'h0;
    end else if(T78) begin
      reg_mstatus_ie <= T243;
    end else if(T60) begin
      reg_mstatus_ie <= T242;
    end else if(insn_ret) begin
      reg_mstatus_ie <= reg_mstatus_ie1;
    end else if(T27) begin
      reg_mstatus_ie <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_ie1 <= 1'h0;
    end else if(T78) begin
      reg_mstatus_ie1 <= T241;
    end else if(T60) begin
      reg_mstatus_ie1 <= T240;
    end else if(insn_ret) begin
      reg_mstatus_ie1 <= reg_mstatus_ie2;
    end else if(T27) begin
      reg_mstatus_ie1 <= reg_mstatus_ie;
    end
    if(reset) begin
      reg_mstatus_ie2 <= 1'h0;
    end else if(T60) begin
      reg_mstatus_ie2 <= T239;
    end else if(insn_ret) begin
      reg_mstatus_ie2 <= 1'h1;
    end else if(T27) begin
      reg_mstatus_ie2 <= reg_mstatus_ie1;
    end
    if(reset) begin
      reg_mip_ssip <= 1'h0;
    end else if(T252) begin
      reg_mip_ssip <= T251;
    end else if(T250) begin
      reg_mip_ssip <= T249;
    end
    if(reset) begin
      reg_mie_ssip <= 1'h0;
    end else if(T258) begin
      reg_mie_ssip <= T257;
    end else if(T256) begin
      reg_mie_ssip <= T255;
    end
    if(reset) begin
      reg_mip_msip <= 1'h0;
    end else if(io_host_ipi_rep_valid) begin
      reg_mip_msip <= 1'h1;
    end else if(T250) begin
      reg_mip_msip <= T267;
    end
    if(reset) begin
      reg_mie_msip <= 1'h0;
    end else if(T256) begin
      reg_mie_msip <= T269;
    end
    if(reset) begin
      reg_mip_stip <= 1'h0;
    end else if(T250) begin
      reg_mip_stip <= T277;
    end
    if(reset) begin
      reg_mie_stip <= 1'h0;
    end else if(T258) begin
      reg_mie_stip <= T281;
    end else if(T256) begin
      reg_mie_stip <= T280;
    end
    if(reset) begin
      reg_mip_mtip <= 1'h0;
    end else if(T294) begin
      reg_mip_mtip <= 1'h0;
    end else if(T290) begin
      reg_mip_mtip <= 1'h1;
    end
    if(T292) begin
      reg_time <= wdata;
    end
    if(T294) begin
      reg_mtimecmp <= wdata;
    end
    if(reset) begin
      reg_mie_mtip <= 1'h0;
    end else if(T256) begin
      reg_mie_mtip <= T296;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T304) begin
      reg_fromhost <= wdata;
    end
    reg_frm <= T896;
    if(reset) begin
      R316 <= 6'h0;
    end else begin
      R316 <= T317;
    end
    if(reset) begin
      R319 <= 58'h0;
    end else if(T322) begin
      R319 <= T321;
    end
    reg_sepc <= T902;
    reg_mepc <= T904;
    reg_stvec <= T906;
    if(T362) begin
      reg_sptbr <= T360;
    end
    if(reset) begin
      reg_mstatus_ie3 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_prv3 <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if(T78) begin
      reg_mstatus_fs <= T371;
    end else if(T60) begin
      reg_mstatus_fs <= T370;
    end
    if(reset) begin
      reg_mstatus_xs <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if(T78) begin
      reg_mstatus_mprv <= T380;
    end else if(T60) begin
      reg_mstatus_mprv <= T379;
    end else if(T27) begin
      reg_mstatus_mprv <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_vm <= 5'h0;
    end else if(T387) begin
      reg_mstatus_vm <= 5'h9;
    end else if(T384) begin
      reg_mstatus_vm <= 5'h0;
    end
    if(reset) begin
      reg_mstatus_zero1 <= 9'h0;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_zero2 <= 31'h0;
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else if(some_interrupt_pending) begin
      reg_wfi <= 1'h0;
    end else if(insn_wfi) begin
      reg_wfi <= 1'h1;
    end
    if(reset) begin
      R424 <= 6'h0;
    end else if(T428) begin
      R424 <= T426;
    end
    if(reset) begin
      R429 <= 58'h0;
    end else if(T432) begin
      R429 <= T431;
    end
    if(reset) begin
      R437 <= 6'h0;
    end else if(T441) begin
      R437 <= T439;
    end
    if(reset) begin
      R442 <= 58'h0;
    end else if(T445) begin
      R442 <= T444;
    end
    if(reset) begin
      R450 <= 6'h0;
    end else if(T454) begin
      R450 <= T452;
    end
    if(reset) begin
      R455 <= 58'h0;
    end else if(T458) begin
      R455 <= T457;
    end
    if(reset) begin
      R463 <= 6'h0;
    end else if(T467) begin
      R463 <= T465;
    end
    if(reset) begin
      R468 <= 58'h0;
    end else if(T471) begin
      R468 <= T470;
    end
    if(reset) begin
      R476 <= 6'h0;
    end else if(T480) begin
      R476 <= T478;
    end
    if(reset) begin
      R481 <= 58'h0;
    end else if(T484) begin
      R481 <= T483;
    end
    if(reset) begin
      R489 <= 6'h0;
    end else if(T493) begin
      R489 <= T491;
    end
    if(reset) begin
      R494 <= 58'h0;
    end else if(T497) begin
      R494 <= T496;
    end
    if(reset) begin
      R502 <= 6'h0;
    end else if(T506) begin
      R502 <= T504;
    end
    if(reset) begin
      R507 <= 58'h0;
    end else if(T510) begin
      R507 <= T509;
    end
    if(reset) begin
      R515 <= 6'h0;
    end else if(T519) begin
      R515 <= T517;
    end
    if(reset) begin
      R520 <= 58'h0;
    end else if(T523) begin
      R520 <= T522;
    end
    if(reset) begin
      R528 <= 6'h0;
    end else if(T532) begin
      R528 <= T530;
    end
    if(reset) begin
      R533 <= 58'h0;
    end else if(T536) begin
      R533 <= T535;
    end
    if(reset) begin
      R541 <= 6'h0;
    end else if(T545) begin
      R541 <= T543;
    end
    if(reset) begin
      R546 <= 58'h0;
    end else if(T549) begin
      R546 <= T548;
    end
    if(reset) begin
      R554 <= 6'h0;
    end else if(T558) begin
      R554 <= T556;
    end
    if(reset) begin
      R559 <= 58'h0;
    end else if(T562) begin
      R559 <= T561;
    end
    if(reset) begin
      R567 <= 6'h0;
    end else if(T571) begin
      R567 <= T569;
    end
    if(reset) begin
      R572 <= 58'h0;
    end else if(T575) begin
      R572 <= T574;
    end
    if(reset) begin
      R580 <= 6'h0;
    end else if(T584) begin
      R580 <= T582;
    end
    if(reset) begin
      R585 <= 58'h0;
    end else if(T588) begin
      R585 <= T587;
    end
    if(reset) begin
      R593 <= 6'h0;
    end else if(T597) begin
      R593 <= T595;
    end
    if(reset) begin
      R598 <= 58'h0;
    end else if(T601) begin
      R598 <= T600;
    end
    if(reset) begin
      R606 <= 6'h0;
    end else if(T610) begin
      R606 <= T608;
    end
    if(reset) begin
      R611 <= 58'h0;
    end else if(T614) begin
      R611 <= T613;
    end
    if(reset) begin
      R619 <= 6'h0;
    end else if(T623) begin
      R619 <= T621;
    end
    if(reset) begin
      R624 <= 58'h0;
    end else if(T627) begin
      R624 <= T626;
    end
    if(insn_redirect_trap) begin
      reg_sbadaddr <= reg_mbadaddr;
    end
    if(T666) begin
      reg_mbadaddr <= T665;
    end else if(T657) begin
      reg_mbadaddr <= T649;
    end else if(T27) begin
      reg_mbadaddr <= io_pc;
    end
    if(insn_redirect_trap) begin
      reg_scause <= reg_mcause;
    end
    if(T682) begin
      reg_mcause <= T681;
    end else if(T680) begin
      reg_mcause <= T965;
    end else if(T678) begin
      reg_mcause <= 64'h3;
    end else if(T677) begin
      reg_mcause <= 64'h2;
    end else if(T27) begin
      reg_mcause <= io_cause;
    end
    if(T686) begin
      reg_sscratch <= wdata;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T781) begin
      reg_tohost <= wdata;
    end else if(T778) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T789) begin
      reg_stats <= T788;
    end
    if(T811) begin
      reg_mscratch <= wdata;
    end
    if(reset) begin
      reg_mie_usip <= 1'h0;
    end
    if(reset) begin
      reg_mie_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mie_utip <= 1'h0;
    end
    if(reset) begin
      reg_mie_htip <= 1'h0;
    end
    if(reset) begin
      reg_mip_usip <= 1'h0;
    end
    if(reset) begin
      reg_mip_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mip_utip <= 1'h0;
    end
    if(reset) begin
      reg_mip_htip <= 1'h0;
    end
    if(reset) begin
      R854 <= 6'h0;
    end else if(T861) begin
      R854 <= T860;
    end else if(T859) begin
      R854 <= T857;
    end
    if(reset) begin
      R862 <= 58'h0;
    end else if(T861) begin
      R862 <= T868;
    end else if(T866) begin
      R862 <= T865;
    end
    if(T878) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T136;
  wire cmp;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] T29;
  wire T30;
  wire[63:0] shout_l;
  wire[63:0] T31;
  wire[63:0] T32;
  wire[62:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[61:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[59:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[55:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[47:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T137;
  wire[31:0] T55;
  wire[63:0] T56;
  wire[63:0] T138;
  wire[47:0] T57;
  wire[63:0] T58;
  wire[63:0] T139;
  wire[55:0] T59;
  wire[63:0] T60;
  wire[63:0] T140;
  wire[59:0] T61;
  wire[63:0] T62;
  wire[63:0] T141;
  wire[61:0] T63;
  wire[63:0] T64;
  wire[63:0] T142;
  wire[62:0] T65;
  wire T66;
  wire[63:0] shout_r;
  wire[64:0] T67;
  wire[5:0] shamt;
  wire[5:0] T68;
  wire[4:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[64:0] T74;
  wire[64:0] T75;
  wire[63:0] shin;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[62:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[61:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[59:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[63:0] T90;
  wire[55:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[63:0] T94;
  wire[47:0] T95;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[63:0] T98;
  wire[31:0] T99;
  wire[63:0] T100;
  wire[63:0] T143;
  wire[31:0] T101;
  wire[63:0] T102;
  wire[63:0] T144;
  wire[47:0] T103;
  wire[63:0] T104;
  wire[63:0] T145;
  wire[55:0] T105;
  wire[63:0] T106;
  wire[63:0] T146;
  wire[59:0] T107;
  wire[63:0] T108;
  wire[63:0] T147;
  wire[61:0] T109;
  wire[63:0] T110;
  wire[63:0] T148;
  wire[62:0] T111;
  wire[63:0] shin_r;
  wire[31:0] T112;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T113;
  wire[31:0] T149;
  wire T114;
  wire T115;
  wire[31:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire[31:0] out_hi;
  wire[31:0] T131;
  wire[31:0] T150;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T128 ? sum : T6;
  assign T6 = T125 ? shout_r : T7;
  assign T7 = T66 ? shout_l : T8;
  assign T8 = T30 ? T29 : T9;
  assign T9 = T28 ? T27 : T10;
  assign T10 = T26 ? T25 : T136;
  assign T136 = {63'h0, cmp};
  assign cmp = T24 ^ T11;
  assign T11 = T22 ? T21 : T12;
  assign T12 = T18 ? T17 : T13;
  assign T13 = T16 ? T15 : T14;
  assign T14 = io_in1[6'h3f:6'h3f];
  assign T15 = io_in2[6'h3f:6'h3f];
  assign T16 = io_fn[1'h1:1'h1];
  assign T17 = sum[6'h3f:6'h3f];
  assign T18 = T20 == T19;
  assign T19 = io_in2[6'h3f:6'h3f];
  assign T20 = io_in1[6'h3f:6'h3f];
  assign T21 = sum == 64'h0;
  assign T22 = T23 ^ 1'h1;
  assign T23 = io_fn[2'h2:2'h2];
  assign T24 = io_fn[1'h0:1'h0];
  assign T25 = io_in1 ^ io_in2;
  assign T26 = io_fn == 4'h4;
  assign T27 = io_in1 | io_in2;
  assign T28 = io_fn == 4'h6;
  assign T29 = io_in1 & io_in2;
  assign T30 = io_fn == 4'h7;
  assign shout_l = T64 | T31;
  assign T31 = T32 & 64'haaaaaaaaaaaaaaaa;
  assign T32 = T33 << 1'h1;
  assign T33 = T34[6'h3e:1'h0];
  assign T34 = T62 | T35;
  assign T35 = T36 & 64'hcccccccccccccccc;
  assign T36 = T37 << 2'h2;
  assign T37 = T38[6'h3d:1'h0];
  assign T38 = T60 | T39;
  assign T39 = T40 & 64'hf0f0f0f0f0f0f0f0;
  assign T40 = T41 << 3'h4;
  assign T41 = T42[6'h3b:1'h0];
  assign T42 = T58 | T43;
  assign T43 = T44 & 64'hff00ff00ff00ff00;
  assign T44 = T45 << 4'h8;
  assign T45 = T46[6'h37:1'h0];
  assign T46 = T56 | T47;
  assign T47 = T48 & 64'hffff0000ffff0000;
  assign T48 = T49 << 5'h10;
  assign T49 = T50[6'h2f:1'h0];
  assign T50 = T54 | T51;
  assign T51 = T52 & 64'hffffffff00000000;
  assign T52 = T53 << 6'h20;
  assign T53 = shout_r[5'h1f:1'h0];
  assign T54 = T137 & 64'hffffffff;
  assign T137 = {32'h0, T55};
  assign T55 = shout_r >> 6'h20;
  assign T56 = T138 & 64'hffff0000ffff;
  assign T138 = {16'h0, T57};
  assign T57 = T50 >> 5'h10;
  assign T58 = T139 & 64'hff00ff00ff00ff;
  assign T139 = {8'h0, T59};
  assign T59 = T46 >> 4'h8;
  assign T60 = T140 & 64'hf0f0f0f0f0f0f0f;
  assign T140 = {4'h0, T61};
  assign T61 = T42 >> 3'h4;
  assign T62 = T141 & 64'h3333333333333333;
  assign T141 = {2'h0, T63};
  assign T63 = T38 >> 2'h2;
  assign T64 = T142 & 64'h5555555555555555;
  assign T142 = {1'h0, T65};
  assign T65 = T34 >> 1'h1;
  assign T66 = io_fn == 4'h1;
  assign shout_r = T67[6'h3f:1'h0];
  assign T67 = $signed(T74) >>> shamt;
  assign shamt = T68;
  assign T68 = {T70, T69};
  assign T69 = io_in2[3'h4:1'h0];
  assign T70 = T73 & T71;
  assign T71 = 1'h1 == T72;
  assign T72 = io_dw & 1'h1;
  assign T73 = io_in2[3'h5:3'h5];
  assign T74 = T75;
  assign T75 = {T122, shin};
  assign shin = T119 ? shin_r : T76;
  assign T76 = T110 | T77;
  assign T77 = T78 & 64'haaaaaaaaaaaaaaaa;
  assign T78 = T79 << 1'h1;
  assign T79 = T80[6'h3e:1'h0];
  assign T80 = T108 | T81;
  assign T81 = T82 & 64'hcccccccccccccccc;
  assign T82 = T83 << 2'h2;
  assign T83 = T84[6'h3d:1'h0];
  assign T84 = T106 | T85;
  assign T85 = T86 & 64'hf0f0f0f0f0f0f0f0;
  assign T86 = T87 << 3'h4;
  assign T87 = T88[6'h3b:1'h0];
  assign T88 = T104 | T89;
  assign T89 = T90 & 64'hff00ff00ff00ff00;
  assign T90 = T91 << 4'h8;
  assign T91 = T92[6'h37:1'h0];
  assign T92 = T102 | T93;
  assign T93 = T94 & 64'hffff0000ffff0000;
  assign T94 = T95 << 5'h10;
  assign T95 = T96[6'h2f:1'h0];
  assign T96 = T100 | T97;
  assign T97 = T98 & 64'hffffffff00000000;
  assign T98 = T99 << 6'h20;
  assign T99 = shin_r[5'h1f:1'h0];
  assign T100 = T143 & 64'hffffffff;
  assign T143 = {32'h0, T101};
  assign T101 = shin_r >> 6'h20;
  assign T102 = T144 & 64'hffff0000ffff;
  assign T144 = {16'h0, T103};
  assign T103 = T96 >> 5'h10;
  assign T104 = T145 & 64'hff00ff00ff00ff;
  assign T145 = {8'h0, T105};
  assign T105 = T92 >> 4'h8;
  assign T106 = T146 & 64'hf0f0f0f0f0f0f0f;
  assign T146 = {4'h0, T107};
  assign T107 = T88 >> 3'h4;
  assign T108 = T147 & 64'h3333333333333333;
  assign T147 = {2'h0, T109};
  assign T109 = T84 >> 2'h2;
  assign T110 = T148 & 64'h5555555555555555;
  assign T148 = {1'h0, T111};
  assign T111 = T80 >> 1'h1;
  assign shin_r = {shin_hi, T112};
  assign T112 = io_in1[5'h1f:1'h0];
  assign shin_hi = T117 ? T116 : shin_hi_32;
  assign shin_hi_32 = T115 ? T113 : 32'h0;
  assign T113 = 32'h0 - T149;
  assign T149 = {31'h0, T114};
  assign T114 = io_in1[5'h1f:5'h1f];
  assign T115 = io_fn[2'h3:2'h3];
  assign T116 = io_in1[6'h3f:6'h20];
  assign T117 = 1'h1 == T118;
  assign T118 = io_dw & 1'h1;
  assign T119 = T121 | T120;
  assign T120 = io_fn == 4'hb;
  assign T121 = io_fn == 4'h5;
  assign T122 = T124 & T123;
  assign T123 = shin[6'h3f:6'h3f];
  assign T124 = io_fn[2'h3:2'h3];
  assign T125 = T127 | T126;
  assign T126 = io_fn == 4'hb;
  assign T127 = io_fn == 4'h5;
  assign T128 = T130 | T129;
  assign T129 = io_fn == 4'ha;
  assign T130 = io_fn == 4'h0;
  assign out_hi = T134 ? T133 : T131;
  assign T131 = 32'h0 - T150;
  assign T150 = {31'h0, T132};
  assign T132 = out64[5'h1f:5'h1f];
  assign T133 = out64[6'h3f:6'h20];
  assign T134 = 1'h1 == T135;
  assign T135 = io_dw & 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T148;
  wire[63:0] negated_remainder;
  wire[63:0] T95;
  wire T10;
  wire T11;
  reg  isMul;
  wire T12;
  wire cmdMul;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  reg [2:0] state;
  wire[2:0] T149;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  reg  neg_out;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  isHi;
  wire T33;
  wire cmdHi;
  wire T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire[3:0] T39;
  wire T40;
  wire T41;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T42;
  wire[64:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[64:0] T47;
  wire[63:0] rhs_in;
  wire[31:0] T48;
  wire[31:0] T49;
  wire[31:0] T50;
  wire[31:0] T150;
  wire[31:0] T51;
  wire T52;
  wire T53;
  wire rhs_sign;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire rhsSigned;
  wire T59;
  wire T60;
  wire[3:0] T61;
  wire[64:0] T62;
  wire T63;
  reg [6:0] count;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[6:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire lhs_sign;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire lhsSigned;
  wire T77;
  wire T78;
  wire[3:0] T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire T83;
  wire T84;
  wire[2:0] T85;
  wire[2:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire[129:0] T151;
  wire T96;
  wire[129:0] T152;
  wire[63:0] T97;
  wire T98;
  wire[129:0] T99;
  wire[64:0] T100;
  wire[63:0] T101;
  wire[128:0] T102;
  wire[63:0] T103;
  wire[128:0] T104;
  wire[128:0] T105;
  wire[62:0] T106;
  wire[63:0] T107;
  wire[128:0] T108;
  wire[63:0] T109;
  wire[64:0] T110;
  wire[65:0] T111;
  wire[65:0] T153;
  wire[64:0] T112;
  wire[64:0] T113;
  wire T154;
  wire[65:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire[64:0] T118;
  wire[64:0] T119;
  wire[64:0] T120;
  wire T121;
  wire T122;
  wire[129:0] T155;
  wire[128:0] T123;
  wire[64:0] T124;
  wire T125;
  wire[63:0] T126;
  wire[63:0] T127;
  wire[63:0] T128;
  wire[63:0] T129;
  wire T130;
  wire T131;
  wire T132;
  wire[129:0] T156;
  wire[63:0] lhs_in;
  wire[31:0] T133;
  wire[31:0] T134;
  wire[31:0] T135;
  wire[31:0] T157;
  wire[31:0] T136;
  wire T137;
  wire T138;
  wire[63:0] T139;
  wire[31:0] T140;
  wire[31:0] T141;
  wire[31:0] T158;
  wire T142;
  wire T143;
  wire T144;
  reg  req_dw;
  wire T145;
  wire T146;
  wire T147;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T143 ? T139 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T156 : T5;
  assign T5 = T130 ? T155 : T6;
  assign T6 = T121 ? T99 : T7;
  assign T7 = T98 ? T152 : T8;
  assign T8 = T96 ? T151 : T9;
  assign T9 = T10 ? T148 : remainder;
  assign T148 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T95;
  assign T95 = remainder[6'h3f:1'h0];
  assign T10 = T19 & T11;
  assign T11 = T18 | isMul;
  assign T12 = T1 ? cmdMul : isMul;
  assign cmdMul = T13;
  assign T13 = T16 | T14;
  assign T14 = T15 == 4'h8;
  assign T15 = io_req_bits_fn & 4'h8;
  assign T16 = T17 == 4'h0;
  assign T17 = io_req_bits_fn & 4'h4;
  assign T18 = remainder[6'h3f:6'h3f];
  assign T19 = state == 3'h1;
  assign T149 = reset ? 3'h0 : T20;
  assign T20 = T1 ? T91 : T21;
  assign T21 = T89 ? 3'h0 : T22;
  assign T22 = T87 ? T85 : T23;
  assign T23 = T83 ? T82 : T24;
  assign T24 = T98 ? T27 : T25;
  assign T25 = T96 ? 3'h5 : T26;
  assign T26 = T19 ? 3'h2 : state;
  assign T27 = neg_out ? 3'h4 : 3'h5;
  assign T28 = T1 ? T69 : T29;
  assign T29 = T30 ? 1'h0 : neg_out;
  assign T30 = T130 & T31;
  assign T31 = T40 & T32;
  assign T32 = isHi ^ 1'h1;
  assign T33 = T1 ? cmdHi : isHi;
  assign cmdHi = T34;
  assign T34 = T35 | T14;
  assign T35 = T38 | T36;
  assign T36 = T37 == 4'h2;
  assign T37 = io_req_bits_fn & 4'h2;
  assign T38 = T39 == 4'h1;
  assign T39 = io_req_bits_fn & 4'h5;
  assign T40 = T63 & T41;
  assign T41 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T62 - divisor;
  assign T42 = T1 ? T47 : T43;
  assign T43 = T44 ? subtractor : divisor;
  assign T44 = T19 & T45;
  assign T45 = T46 | isMul;
  assign T46 = divisor[6'h3f:6'h3f];
  assign T47 = {rhs_sign, rhs_in};
  assign rhs_in = {T49, T48};
  assign T48 = io_req_bits_in2[5'h1f:1'h0];
  assign T49 = T52 ? T51 : T50;
  assign T50 = 32'h0 - T150;
  assign T150 = {31'h0, rhs_sign};
  assign T51 = io_req_bits_in2[6'h3f:6'h20];
  assign T52 = 1'h1 == T53;
  assign T53 = io_req_bits_dw & 1'h1;
  assign rhs_sign = rhsSigned & T54;
  assign T54 = T57 ? T56 : T55;
  assign T55 = io_req_bits_in2[5'h1f:5'h1f];
  assign T56 = io_req_bits_in2[6'h3f:6'h3f];
  assign T57 = 1'h1 == T58;
  assign T58 = io_req_bits_dw & 1'h1;
  assign rhsSigned = T59;
  assign T59 = T60 | T16;
  assign T60 = T61 == 4'h0;
  assign T61 = io_req_bits_fn & 4'h9;
  assign T62 = remainder[8'h80:7'h40];
  assign T63 = count == 7'h0;
  assign T64 = T1 ? 7'h0 : T65;
  assign T65 = T130 ? T68 : T66;
  assign T66 = T121 ? T67 : count;
  assign T67 = count + 7'h1;
  assign T68 = count + 7'h1;
  assign T69 = T81 & T70;
  assign T70 = cmdHi ? lhs_sign : T71;
  assign T71 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T72;
  assign T72 = T75 ? T74 : T73;
  assign T73 = io_req_bits_in1[5'h1f:5'h1f];
  assign T74 = io_req_bits_in1[6'h3f:6'h3f];
  assign T75 = 1'h1 == T76;
  assign T76 = io_req_bits_dw & 1'h1;
  assign lhsSigned = T77;
  assign T77 = T80 | T78;
  assign T78 = T79 == 4'h0;
  assign T79 = io_req_bits_fn & 4'h3;
  assign T80 = T60 | T16;
  assign T81 = cmdMul ^ 1'h1;
  assign T82 = isHi ? 3'h3 : 3'h5;
  assign T83 = T121 & T84;
  assign T84 = count == 7'h3f;
  assign T85 = isHi ? 3'h3 : T86;
  assign T86 = neg_out ? 3'h4 : 3'h5;
  assign T87 = T130 & T88;
  assign T88 = count == 7'h40;
  assign T89 = T90 | io_kill;
  assign T90 = io_resp_ready & io_resp_valid;
  assign T91 = T92 ? 3'h1 : 3'h2;
  assign T92 = lhs_sign | T93;
  assign T93 = rhs_sign & T94;
  assign T94 = cmdMul ^ 1'h1;
  assign T151 = {66'h0, negated_remainder};
  assign T96 = state == 3'h4;
  assign T152 = {66'h0, T97};
  assign T97 = remainder[8'h80:7'h41];
  assign T98 = state == 3'h3;
  assign T99 = {T120, T100};
  assign T100 = {1'h0, T101};
  assign T101 = T102[6'h3f:1'h0];
  assign T102 = {T119, T103};
  assign T103 = T104[6'h3f:1'h0];
  assign T104 = T105;
  assign T105 = {T111, T106};
  assign T106 = T107[6'h3f:1'h1];
  assign T107 = T108[6'h3f:1'h0];
  assign T108 = {T110, T109};
  assign T109 = remainder[6'h3f:1'h0];
  assign T110 = remainder[8'h81:7'h41];
  assign T111 = T114 + T153;
  assign T153 = {T154, T112};
  assign T112 = T113;
  assign T113 = T108[8'h80:7'h40];
  assign T154 = T112[7'h40:7'h40];
  assign T114 = $signed(T118) * $signed(T115);
  assign T115 = T116;
  assign T116 = {1'h0, T117};
  assign T117 = T107[1'h0:1'h0];
  assign T118 = divisor;
  assign T119 = T104[8'h80:7'h40];
  assign T120 = T102 >> 7'h40;
  assign T121 = T122 & isMul;
  assign T122 = state == 3'h2;
  assign T155 = {1'h0, T123};
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = less ^ 1'h1;
  assign T126 = remainder[6'h3f:1'h0];
  assign T127 = less ? T129 : T128;
  assign T128 = subtractor[6'h3f:1'h0];
  assign T129 = remainder[7'h7f:7'h40];
  assign T130 = T132 & T131;
  assign T131 = isMul ^ 1'h1;
  assign T132 = state == 3'h2;
  assign T156 = {66'h0, lhs_in};
  assign lhs_in = {T134, T133};
  assign T133 = io_req_bits_in1[5'h1f:1'h0];
  assign T134 = T137 ? T136 : T135;
  assign T135 = 32'h0 - T157;
  assign T157 = {31'h0, lhs_sign};
  assign T136 = io_req_bits_in1[6'h3f:6'h20];
  assign T137 = 1'h1 == T138;
  assign T138 = io_req_bits_dw & 1'h1;
  assign T139 = {T141, T140};
  assign T140 = remainder[5'h1f:1'h0];
  assign T141 = 32'h0 - T158;
  assign T158 = {31'h0, T142};
  assign T142 = remainder[5'h1f:5'h1f];
  assign T143 = 1'h0 == T144;
  assign T144 = req_dw & 1'h1;
  assign T145 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T146;
  assign T146 = state == 3'h5;
  assign io_req_ready = T147;
  assign T147 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T156;
    end else if(T130) begin
      remainder <= T155;
    end else if(T121) begin
      remainder <= T99;
    end else if(T98) begin
      remainder <= T152;
    end else if(T96) begin
      remainder <= T151;
    end else if(T10) begin
      remainder <= T148;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T91;
    end else if(T89) begin
      state <= 3'h0;
    end else if(T87) begin
      state <= T85;
    end else if(T83) begin
      state <= T82;
    end else if(T98) begin
      state <= T27;
    end else if(T96) begin
      state <= 3'h5;
    end else if(T19) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T69;
    end else if(T30) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T47;
    end else if(T44) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T130) begin
      count <= T68;
    end else if(T121) begin
      count <= T67;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module Rocket(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [11:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[39:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [39:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [38:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_btb_update_bits_pc,
    output[38:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output[38:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_bht_update_bits_prediction_bits_target,
    output[2:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[3:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output[38:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_ras_update_bits_prediction_bits_target,
    output[2:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[3:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    output io_imem_invalidate,
    input [39:0] io_imem_npc,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output[39:0] io_dmem_req_bits_addr,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_kill,
    output io_dmem_req_bits_phys,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [39:0] io_dmem_resp_bits_addr,
    input [7:0] io_dmem_resp_bits_tag,
    input [4:0] io_dmem_resp_bits_cmd,
    input [2:0] io_dmem_resp_bits_typ,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    output io_dmem_invalidate_lr,
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_status_sd,
    output[30:0] io_ptw_status_zero2,
    output io_ptw_status_sd_rv32,
    output[8:0] io_ptw_status_zero1,
    output[4:0] io_ptw_status_vm,
    output io_ptw_status_mprv,
    output[1:0] io_ptw_status_xs,
    output[1:0] io_ptw_status_fs,
    output[1:0] io_ptw_status_prv3,
    output io_ptw_status_ie3,
    output[1:0] io_ptw_status_prv2,
    output io_ptw_status_ie2,
    output[1:0] io_ptw_status_prv1,
    output io_ptw_status_ie1,
    output[1:0] io_ptw_status_prv,
    output io_ptw_status_ie,
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    output io_fpu_valid,
    //input  io_fpu_fcsr_rdy
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    //input [4:0] io_fpu_dec_cmd
    //input  io_fpu_dec_ldst
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    //input  io_fpu_dec_swap12
    //input  io_fpu_dec_swap23
    //input  io_fpu_dec_single
    //input  io_fpu_dec_fromint
    //input  io_fpu_dec_toint
    //input  io_fpu_dec_fastpipe
    //input  io_fpu_dec_fma
    //input  io_fpu_dec_div
    //input  io_fpu_dec_sqrt
    //input  io_fpu_dec_round
    //input  io_fpu_dec_wflags
    //input  io_fpu_sboard_set
    //input  io_fpu_sboard_clr
    //input [4:0] io_fpu_sboard_clra
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [25:0] io_rocc_imem_acquire_bits_addr_block,
    input  io_rocc_imem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_imem_acquire_bits_addr_beat,
    input [127:0] io_rocc_imem_acquire_bits_data,
    input  io_rocc_imem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_imem_acquire_bits_a_type,
    input [16:0] io_rocc_imem_acquire_bits_union,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_addr_beat
    //output[127:0] io_rocc_imem_grant_bits_data
    //output io_rocc_imem_grant_bits_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_manager_xact_id
    //output io_rocc_imem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_imem_grant_bits_g_type
    //output io_rocc_dmem_acquire_ready
    input  io_rocc_dmem_acquire_valid,
    input [25:0] io_rocc_dmem_acquire_bits_addr_block,
    input  io_rocc_dmem_acquire_bits_client_xact_id,
    input [1:0] io_rocc_dmem_acquire_bits_addr_beat,
    input [127:0] io_rocc_dmem_acquire_bits_data,
    input  io_rocc_dmem_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_dmem_acquire_bits_a_type,
    input [16:0] io_rocc_dmem_acquire_bits_union,
    input  io_rocc_dmem_grant_ready,
    //output io_rocc_dmem_grant_valid
    //output[1:0] io_rocc_dmem_grant_bits_addr_beat
    //output[127:0] io_rocc_dmem_grant_bits_data
    //output io_rocc_dmem_grant_bits_client_xact_id
    //output[2:0] io_rocc_dmem_grant_bits_manager_xact_id
    //output io_rocc_dmem_grant_bits_is_builtin_type
    //output[3:0] io_rocc_dmem_grant_bits_g_type
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  wire ctrl_killd;
  wire T7;
  wire T8;
  wire ctrl_stalld;
  wire T9;
  wire id_do_fence;
  wire T10;
  wire id_csr_en;
  wire[2:0] id_ctrl_csr;
  wire[2:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire[31:0] T16;
  wire T17;
  wire[31:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire id_ctrl_rocc;
  wire id_ctrl_mem;
  wire T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire[31:0] T38;
  reg  id_reg_fence;
  wire T916;
  wire T39;
  wire T40;
  wire id_fence_next;
  wire T41;
  wire id_amo_rl;
  wire id_ctrl_amo;
  wire T42;
  wire[31:0] T43;
  wire id_ctrl_fence;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire id_ctrl_fence_i;
  wire T47;
  wire[31:0] T48;
  wire T49;
  wire id_amo_aq;
  wire id_mem_busy;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire id_sboard_hazard;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[4:0] T59;
  wire[4:0] T60;
  wire[4:0] id_waddr_1;
  wire T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[4:0] ll_waddr;
  wire[4:0] T66;
  wire[4:0] dmem_resp_waddr;
  wire[7:0] T67;
  wire T68;
  wire dmem_resp_xpu;
  wire T69;
  wire T70;
  wire dmem_resp_replay;
  wire ll_wen;
  wire T71;
  wire T72;
  reg [31:0] R73;
  wire[31:0] T917;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[31:0] T76;
  wire[31:0] T77;
  wire[31:0] T78;
  wire[4:0] wb_waddr;
  wire T79;
  wire wb_wen;
  reg  wb_ctrl_wxd;
  wire T80;
  reg  mem_ctrl_wxd;
  wire T81;
  reg  ex_ctrl_wxd;
  wire T82;
  wire id_ctrl_wxd;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire[31:0] T91;
  wire T92;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire T96;
  wire[31:0] T97;
  wire T98;
  wire T99;
  wire[31:0] T100;
  wire T101;
  wire[31:0] T102;
  wire T103;
  wire wb_valid;
  wire T104;
  wire T105;
  wire T106;
  wire replay_wb;
  wire T107;
  wire T108;
  wire T109;
  reg  wb_ctrl_rocc;
  wire T110;
  reg  mem_ctrl_rocc;
  wire T111;
  reg  ex_ctrl_rocc;
  wire T112;
  wire replay_wb_common;
  wire T113;
  reg  wb_reg_replay;
  wire T114;
  wire T115;
  wire take_pc_wb;
  wire T116;
  wire T117;
  wire wb_xcpt;
  reg  wb_reg_xcpt;
  wire T118;
  wire T119;
  wire mem_xcpt;
  wire T120;
  wire T121;
  reg  mem_ctrl_mem;
  wire T122;
  reg  ex_ctrl_mem;
  wire T123;
  reg  mem_reg_valid;
  wire T124;
  wire ctrl_killx;
  wire T125;
  reg  ex_reg_valid;
  wire T126;
  wire T127;
  wire replay_ex;
  wire T128;
  wire replay_ex_load_use;
  reg  ex_reg_load_use;
  wire T129;
  wire id_load_use;
  wire T130;
  wire T131;
  wire data_hazard_mem;
  wire T132;
  wire T133;
  wire T134;
  wire[4:0] mem_waddr;
  wire T135;
  wire T136;
  wire T137;
  wire[4:0] id_raddr_1;
  wire T138;
  wire T139;
  wire id_ctrl_rxs2;
  wire T140;
  wire T141;
  wire[31:0] T142;
  wire T143;
  wire T144;
  wire[31:0] T145;
  wire T146;
  wire[31:0] T147;
  wire T148;
  wire T149;
  wire[4:0] id_raddr_0;
  wire T150;
  wire T151;
  wire id_ctrl_rxs1;
  wire T152;
  wire T153;
  wire[31:0] T154;
  wire T155;
  wire T156;
  wire[31:0] T157;
  wire T158;
  wire T159;
  wire[31:0] T160;
  wire T161;
  wire[31:0] T162;
  wire wb_dcache_miss;
  wire T163;
  reg  wb_ctrl_mem;
  wire T164;
  wire replay_ex_structural;
  wire T165;
  wire T166;
  reg  ex_ctrl_div;
  wire T167;
  wire id_ctrl_div;
  wire T168;
  wire[31:0] T169;
  wire T170;
  wire T171;
  wire take_pc;
  wire take_pc_mem;
  wire T172;
  wire T173;
  wire mem_npc_misaligned;
  wire[39:0] mem_npc;
  wire[39:0] T174;
  wire[39:0] T175;
  wire[39:0] mem_br_target;
  wire[39:0] T918;
  wire[21:0] T176;
  wire[21:0] T177;
  wire[21:0] T178;
  wire[21:0] T179;
  wire[11:0] T180;
  wire[4:0] T181;
  wire[3:0] T182;
  wire[6:0] T183;
  wire[5:0] T184;
  wire T185;
  wire T186;
  wire[9:0] T187;
  wire[8:0] T188;
  wire[7:0] T189;
  wire[7:0] T190;
  wire T191;
  wire T192;
  reg  mem_ctrl_jal;
  wire T193;
  reg  ex_ctrl_jal;
  wire T194;
  wire id_ctrl_jal;
  wire[21:0] T919;
  wire[14:0] T195;
  wire[14:0] T196;
  wire[11:0] T197;
  wire[4:0] T198;
  wire[3:0] T199;
  wire[6:0] T200;
  wire[5:0] T201;
  wire T202;
  wire T203;
  wire[2:0] T204;
  wire[1:0] T205;
  wire T206;
  wire T207;
  wire[6:0] T920;
  wire T921;
  wire T208;
  wire mem_br_taken;
  reg [63:0] bypass_mux_1;
  wire[63:0] T209;
  reg  mem_ctrl_branch;
  wire T210;
  reg  ex_ctrl_branch;
  wire T211;
  wire id_ctrl_branch;
  wire T212;
  wire[31:0] T213;
  wire[17:0] T922;
  wire T923;
  wire[39:0] T214;
  reg [39:0] mem_reg_pc;
  wire[39:0] T215;
  reg [39:0] ex_reg_pc;
  wire[39:0] T216;
  wire[39:0] T217;
  wire[39:0] T218;
  wire[38:0] T219;
  wire T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire T224;
  wire[1:0] T225;
  wire T226;
  wire T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire T230;
  wire[25:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  reg  mem_ctrl_jalr;
  wire T236;
  reg  ex_ctrl_jalr;
  wire T237;
  wire id_ctrl_jalr;
  wire T238;
  wire[31:0] T239;
  wire want_take_pc_mem;
  wire T240;
  reg  mem_reg_flush_pipe;
  wire T241;
  reg  ex_reg_flush_pipe;
  wire T242;
  wire T243;
  wire id_csr_flush;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  wire[11:0] id_csr_addr;
  wire T249;
  wire T250;
  wire id_csr_ren;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire id_system_insn;
  wire mem_misprediction;
  wire T255;
  wire T256;
  wire T257;
  wire mem_wrong_npc;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  reg  mem_reg_xcpt;
  wire T272;
  wire ex_xcpt;
  wire T273;
  reg  ex_ctrl_fp;
  wire T274;
  wire id_ctrl_fp;
  wire T275;
  reg  ex_reg_xcpt;
  wire T276;
  wire id_xcpt;
  wire id_illegal_insn;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire id_ctrl_legal;
  wire T285;
  wire T286;
  wire[31:0] T287;
  wire T288;
  wire T289;
  wire[31:0] T290;
  wire T291;
  wire T292;
  wire[31:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[31:0] T298;
  wire T299;
  wire T300;
  wire T301;
  wire[31:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire[31:0] T306;
  wire T307;
  wire T308;
  wire[31:0] T309;
  wire T310;
  wire T311;
  wire[31:0] T312;
  wire T313;
  wire T314;
  wire[31:0] T315;
  wire T316;
  wire T317;
  wire[31:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire[31:0] T322;
  wire T323;
  wire T324;
  wire[31:0] T325;
  wire T326;
  wire T327;
  wire[31:0] T328;
  wire T329;
  wire T330;
  wire[31:0] T331;
  wire T332;
  wire T333;
  wire[31:0] T334;
  wire T335;
  wire T336;
  wire[31:0] T337;
  wire T338;
  wire T339;
  wire[31:0] T340;
  wire T341;
  wire T342;
  wire[31:0] T343;
  wire T344;
  wire T345;
  wire[31:0] T346;
  wire T347;
  wire T348;
  wire[31:0] T349;
  wire T350;
  wire T351;
  wire[31:0] T352;
  wire T353;
  wire T354;
  wire[31:0] T355;
  wire T356;
  wire T357;
  wire T358;
  reg  ex_reg_xcpt_interrupt;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  reg  mem_reg_xcpt_interrupt;
  wire T363;
  wire T364;
  wire replay_mem;
  wire fpu_kill_mem;
  wire T365;
  reg  mem_ctrl_fp;
  wire T366;
  wire T367;
  reg  mem_reg_replay;
  wire T368;
  wire T369;
  wire dcache_kill_mem;
  wire T370;
  reg  wb_reg_valid;
  wire T371;
  wire ctrl_killm;
  wire T372;
  wire killm_common;
  wire T373;
  wire T374;
  wire T375;
  wire wb_set_sboard;
  wire T376;
  reg  wb_ctrl_div;
  wire T377;
  reg  mem_ctrl_div;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire[4:0] T394;
  wire[4:0] T395;
  wire T396;
  wire T397;
  wire id_wb_hazard;
  wire T398;
  wire fp_data_hazard_wb;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire[4:0] id_raddr3;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  reg  wb_ctrl_wfd;
  wire T410;
  reg  mem_ctrl_wfd;
  wire T411;
  reg  ex_ctrl_wfd;
  wire T412;
  wire id_ctrl_wfd;
  wire T413;
  wire data_hazard_wb;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire id_mem_hazard;
  wire T423;
  wire fp_data_hazard_mem;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire mem_cannot_bypass;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  reg  mem_mem_cmd_bh;
  wire T440;
  wire ex_slow_bypass;
  wire T441;
  wire T442;
  reg [2:0] ex_ctrl_mem_type;
  wire[2:0] T443;
  wire[2:0] id_ctrl_mem_type;
  wire[2:0] T444;
  wire[1:0] T445;
  wire T446;
  wire[31:0] T447;
  wire T448;
  wire[31:0] T449;
  wire T450;
  wire[31:0] T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  reg [4:0] ex_ctrl_mem_cmd;
  wire[4:0] T458;
  wire[4:0] id_ctrl_mem_cmd;
  wire[4:0] T459;
  wire[3:0] T460;
  wire[2:0] T461;
  wire[1:0] T462;
  wire T463;
  wire T464;
  wire[31:0] T465;
  wire T466;
  wire T467;
  wire[31:0] T468;
  wire T469;
  wire[31:0] T470;
  wire T471;
  wire T472;
  wire[31:0] T473;
  wire T474;
  wire[31:0] T475;
  wire T476;
  wire T477;
  wire[31:0] T478;
  wire T479;
  wire T480;
  wire[31:0] T481;
  wire T482;
  wire[31:0] T483;
  wire T484;
  reg [2:0] mem_ctrl_csr;
  wire[2:0] T485;
  reg [2:0] ex_ctrl_csr;
  wire[2:0] T486;
  wire[2:0] T487;
  wire[2:0] id_csr;
  wire id_ex_hazard;
  wire T488;
  wire fp_data_hazard_ex;
  wire T489;
  wire T490;
  wire T491;
  wire[4:0] ex_waddr;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire ex_cannot_bypass;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire data_hazard_ex;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire[31:0] T519;
  wire[63:0] T520;
  reg [63:0] R521;
  reg [63:0] R522;
  wire[63:0] ex_rs_1;
  wire[63:0] T523;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire[1:0] T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire[1:0] T538;
  wire[63:0] id_rs_1;
  wire[63:0] T539;
  wire[63:0] T540;
  reg [63:0] T541 [30:0];
  wire[63:0] T542;
  wire T543;
  wire T544;
  wire[4:0] T545;
  wire T546;
  wire T547;
  wire[4:0] rf_waddr;
  wire rf_wen;
  wire[4:0] T548;
  wire[4:0] T549;
  wire[63:0] rf_wdata;
  wire[63:0] T550;
  wire[63:0] T551;
  reg [63:0] bypass_mux_2;
  wire[63:0] T552;
  wire[63:0] T553;
  wire[63:0] mem_int_wdata;
  wire[63:0] T554;
  wire[63:0] T555;
  wire[63:0] T924;
  wire[23:0] T925;
  wire T926;
  wire T556;
  wire T557;
  reg [2:0] wb_ctrl_csr;
  wire[2:0] T558;
  wire[63:0] ll_wdata;
  wire T559;
  wire dmem_resp_valid;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T571;
  wire[61:0] T572;
  wire[63:0] T573;
  wire[63:0] T574;
  wire T575;
  wire[1:0] T576;
  wire[63:0] T577;
  wire T578;
  wire T579;
  reg  ex_reg_rs_bypass_1;
  wire T580;
  wire[4:0] T581;
  wire[4:0] T582;
  wire[63:0] T583;
  reg [63:0] R584;
  reg [63:0] R585;
  wire[63:0] ex_rs_0;
  wire[63:0] T586;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[1:0] T597;
  wire[63:0] id_rs_0;
  wire[63:0] T598;
  wire[63:0] T599;
  wire[4:0] T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T611;
  wire[61:0] T612;
  wire[63:0] T613;
  wire[63:0] T614;
  wire T615;
  wire[1:0] T616;
  wire[63:0] T617;
  wire T618;
  wire T619;
  reg  ex_reg_rs_bypass_0;
  wire T620;
  wire[4:0] T621;
  wire[4:0] T622;
  wire T623;
  wire[63:0] T624;
  wire[4:0] T625;
  wire[4:0] T626;
  wire[39:0] T627;
  reg [39:0] wb_reg_pc;
  wire[39:0] T628;
  wire T629;
  wire[32:0] T630;
  wire[32:0] T631;
  wire T632;
  wire[1127:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  reg  R638;
  wire T639;
  reg  ex_ctrl_alu_dw;
  wire T640;
  wire id_ctrl_alu_dw;
  wire T641;
  wire T642;
  wire[31:0] T643;
  wire T644;
  wire[31:0] T645;
  reg [3:0] ex_ctrl_alu_fn;
  wire[3:0] T646;
  wire[3:0] id_ctrl_alu_fn;
  wire[3:0] T647;
  wire[2:0] T648;
  wire[1:0] T649;
  wire T650;
  wire T651;
  wire[31:0] T652;
  wire T653;
  wire T654;
  wire[31:0] T655;
  wire T656;
  wire[31:0] T657;
  wire T658;
  wire T659;
  wire[31:0] T660;
  wire T661;
  wire T662;
  wire[31:0] T663;
  wire T664;
  wire T665;
  wire[31:0] T666;
  wire T667;
  wire T668;
  wire[31:0] T669;
  wire T670;
  wire[31:0] T671;
  wire T672;
  wire T673;
  wire[31:0] T674;
  wire T675;
  wire T676;
  wire[31:0] T677;
  wire T678;
  wire T679;
  wire[31:0] T680;
  wire T681;
  wire[31:0] T682;
  wire T683;
  wire T684;
  wire[31:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[31:0] T689;
  wire T690;
  wire[63:0] T691;
  wire[63:0] ex_op1;
  wire[63:0] T927;
  wire[39:0] T692;
  wire[39:0] T693;
  wire T694;
  reg [1:0] ex_ctrl_sel_alu1;
  wire[1:0] T695;
  wire[1:0] id_ctrl_sel_alu1;
  wire[1:0] T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire[31:0] T701;
  wire T702;
  wire T703;
  wire[31:0] T704;
  wire[23:0] T928;
  wire T929;
  wire[63:0] T705;
  wire T706;
  wire[63:0] T707;
  wire[63:0] ex_op2;
  wire[63:0] T930;
  wire[31:0] T708;
  wire[31:0] T931;
  wire[3:0] T709;
  wire T710;
  reg [1:0] ex_ctrl_sel_alu2;
  wire[1:0] T711;
  wire[1:0] id_ctrl_sel_alu2;
  wire[1:0] T712;
  wire T713;
  wire T714;
  wire[31:0] T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[31:0] T720;
  wire T721;
  wire[31:0] T722;
  wire T723;
  wire T724;
  wire[31:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[31:0] T729;
  wire[27:0] T932;
  wire T933;
  wire[31:0] ex_imm;
  wire[31:0] T730;
  wire[11:0] T731;
  wire[4:0] T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  reg [2:0] ex_ctrl_sel_imm;
  wire[2:0] T738;
  wire[2:0] id_ctrl_sel_imm;
  wire[2:0] T739;
  wire[1:0] T740;
  wire T741;
  wire T742;
  wire[31:0] T743;
  wire T744;
  wire[31:0] T745;
  wire T746;
  wire T747;
  wire[31:0] T748;
  wire T749;
  wire T750;
  wire[31:0] T751;
  wire T752;
  wire T753;
  wire[31:0] T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire[3:0] T759;
  wire[3:0] T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire T764;
  wire[3:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire[6:0] T770;
  wire[5:0] T771;
  wire[5:0] T772;
  wire T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire[19:0] T792;
  wire[18:0] T793;
  wire[7:0] T794;
  wire[7:0] T795;
  wire[7:0] T796;
  wire[7:0] T934;
  wire T797;
  wire T798;
  wire T799;
  wire[10:0] T800;
  wire[10:0] T935;
  wire[10:0] T801;
  wire[10:0] T802;
  wire T803;
  wire T804;
  wire[31:0] T936;
  wire T937;
  wire[63:0] T805;
  wire T806;
  reg [63:0] wb_reg_cause;
  wire[63:0] T807;
  wire[63:0] mem_cause;
  wire[63:0] T938;
  wire[2:0] T808;
  wire[2:0] T809;
  wire[2:0] T810;
  wire[2:0] T811;
  reg [63:0] mem_reg_cause;
  wire[63:0] T812;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T813;
  wire[63:0] id_cause;
  wire[63:0] T939;
  wire[1:0] T814;
  wire[2:0] T815;
  wire[11:0] T816;
  wire T817;
  wire T818;
  wire T819;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T820;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T821;
  wire T822;
  wire T823;
  wire T824;
  reg  ex_ctrl_rxs2;
  wire T825;
  wire T826;
  wire[6:0] T827;
  wire[4:0] T828;
  wire T829;
  wire T830;
  wire T831;
  wire[4:0] T832;
  wire[4:0] T833;
  wire[6:0] T834;
  wire wb_rocc_val;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire dmem_resp_fpu;
  wire T840;
  wire[63:0] T841;
  wire T842;
  wire[7:0] T940;
  wire[5:0] T843;
  wire[39:0] T844;
  wire[39:0] T845;
  wire[38:0] T846;
  wire T847;
  wire T848;
  wire T849;
  wire[1:0] T850;
  wire T851;
  wire[1:0] T852;
  wire T853;
  wire T854;
  wire[25:0] T855;
  wire[25:0] T856;
  wire T857;
  wire[25:0] T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  reg  wb_ctrl_fence_i;
  wire T865;
  reg  mem_ctrl_fence_i;
  wire T866;
  reg  ex_ctrl_fence_i;
  wire T867;
  wire[38:0] T941;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire[38:0] T942;
  wire T875;
  wire T876;
  wire T877;
  wire[38:0] T943;
  wire T878;
  wire T879;
  wire[4:0] T880;
  wire[4:0] T881;
  wire T882;
  wire[38:0] T944;
  wire[38:0] T945;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T883;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T884;
  wire T885;
  wire T886;
  reg  ex_reg_btb_hit;
  wire T887;
  reg [3:0] mem_reg_btb_resp_bht_history;
  wire[3:0] T888;
  reg [3:0] ex_reg_btb_resp_bht_history;
  wire[3:0] T889;
  reg [2:0] mem_reg_btb_resp_entry;
  wire[2:0] T890;
  reg [2:0] ex_reg_btb_resp_entry;
  wire[2:0] T891;
  reg [38:0] mem_reg_btb_resp_target;
  wire[38:0] T892;
  reg [38:0] ex_reg_btb_resp_target;
  wire[38:0] T893;
  reg  mem_reg_btb_resp_bridx;
  wire T894;
  reg  ex_reg_btb_resp_bridx;
  wire T895;
  reg  mem_reg_btb_resp_mask;
  wire T896;
  reg  ex_reg_btb_resp_mask;
  wire T897;
  reg  mem_reg_btb_resp_taken;
  wire T898;
  reg  ex_reg_btb_resp_taken;
  wire T899;
  reg  mem_reg_btb_hit;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire[39:0] T912;
  wire[39:0] T913;
  wire[39:0] T914;
  wire T915;
  wire csr_io_host_pcr_req_ready;
  wire csr_io_host_pcr_rep_valid;
  wire[63:0] csr_io_host_pcr_rep_bits;
  wire csr_io_host_ipi_req_valid;
  wire csr_io_host_ipi_req_bits;
  wire csr_io_host_ipi_rep_ready;
  wire csr_io_host_debug_stats_pcr;
  wire[63:0] csr_io_rw_rdata;
  wire csr_io_csr_replay;
  wire csr_io_csr_stall;
  wire csr_io_csr_xcpt;
  wire csr_io_eret;
  wire csr_io_status_sd;
  wire[30:0] csr_io_status_zero2;
  wire csr_io_status_sd_rv32;
  wire[8:0] csr_io_status_zero1;
  wire[4:0] csr_io_status_vm;
  wire csr_io_status_mprv;
  wire[1:0] csr_io_status_xs;
  wire[1:0] csr_io_status_fs;
  wire[1:0] csr_io_status_prv3;
  wire csr_io_status_ie3;
  wire[1:0] csr_io_status_prv2;
  wire csr_io_status_ie2;
  wire[1:0] csr_io_status_prv1;
  wire csr_io_status_ie1;
  wire[1:0] csr_io_status_prv;
  wire csr_io_status_ie;
  wire[31:0] csr_io_ptbr;
  wire[39:0] csr_io_evec;
  wire csr_io_fatc;
  wire[63:0] csr_io_time;
  wire[2:0] csr_io_fcsr_rm;
  wire csr_io_interrupt;
  wire[63:0] csr_io_interrupt_cause;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    id_reg_fence = {1{$random}};
    R73 = {1{$random}};
    wb_ctrl_wxd = {1{$random}};
    mem_ctrl_wxd = {1{$random}};
    ex_ctrl_wxd = {1{$random}};
    wb_ctrl_rocc = {1{$random}};
    mem_ctrl_rocc = {1{$random}};
    ex_ctrl_rocc = {1{$random}};
    wb_reg_replay = {1{$random}};
    wb_reg_xcpt = {1{$random}};
    mem_ctrl_mem = {1{$random}};
    ex_ctrl_mem = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    ex_reg_load_use = {1{$random}};
    wb_ctrl_mem = {1{$random}};
    ex_ctrl_div = {1{$random}};
    mem_ctrl_jal = {1{$random}};
    ex_ctrl_jal = {1{$random}};
    bypass_mux_1 = {2{$random}};
    mem_ctrl_branch = {1{$random}};
    ex_ctrl_branch = {1{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    mem_ctrl_jalr = {1{$random}};
    ex_ctrl_jalr = {1{$random}};
    mem_reg_flush_pipe = {1{$random}};
    ex_reg_flush_pipe = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_ctrl_fp = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    mem_ctrl_fp = {1{$random}};
    mem_reg_replay = {1{$random}};
    wb_reg_valid = {1{$random}};
    wb_ctrl_div = {1{$random}};
    mem_ctrl_div = {1{$random}};
    wb_ctrl_wfd = {1{$random}};
    mem_ctrl_wfd = {1{$random}};
    ex_ctrl_wfd = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_ctrl_mem_type = {1{$random}};
    ex_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_csr = {1{$random}};
    ex_ctrl_csr = {1{$random}};
    R521 = {2{$random}};
    R522 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T541[initvar] = {2{$random}};
    bypass_mux_2 = {2{$random}};
    wb_ctrl_csr = {1{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R584 = {2{$random}};
    R585 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    R638 = {1{$random}};
    ex_ctrl_alu_dw = {1{$random}};
    ex_ctrl_alu_fn = {1{$random}};
    ex_ctrl_sel_alu1 = {1{$random}};
    ex_ctrl_sel_alu2 = {1{$random}};
    ex_ctrl_sel_imm = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
    ex_ctrl_rxs2 = {1{$random}};
    wb_ctrl_fence_i = {1{$random}};
    mem_ctrl_fence_i = {1{$random}};
    ex_ctrl_fence_i = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_bridx = {1{$random}};
    ex_reg_btb_resp_bridx = {1{$random}};
    mem_reg_btb_resp_mask = {1{$random}};
    ex_reg_btb_resp_mask = {1{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_dmem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_dmem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dmem_grant_bits_data = {4{$random}};
//  assign io_rocc_dmem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_dmem_grant_valid = {1{$random}};
//  assign io_rocc_dmem_acquire_ready = {1{$random}};
//  assign io_rocc_imem_grant_bits_g_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_imem_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_imem_grant_bits_data = {4{$random}};
//  assign io_rocc_imem_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_imem_grant_valid = {1{$random}};
//  assign io_rocc_imem_acquire_ready = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_subword = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_imem_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T517 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T516 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign T5 = T6 | csr_io_interrupt;
  assign T6 = ctrl_killd ^ 1'h1;
  assign ctrl_killd = T7;
  assign T7 = T8 | csr_io_interrupt;
  assign T8 = T514 | ctrl_stalld;
  assign ctrl_stalld = T9 | csr_io_csr_stall;
  assign T9 = T51 | id_do_fence;
  assign id_do_fence = id_mem_busy & T10;
  assign T10 = T19 | id_csr_en;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_ctrl_csr = T11;
  assign T11 = {T17, T12};
  assign T12 = {T15, T13};
  assign T13 = T14 == 32'h1050;
  assign T14 = io_imem_resp_bits_data_0 & 32'h1050;
  assign T15 = T16 == 32'h2050;
  assign T16 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T17 = T18 == 32'h50;
  assign T18 = io_imem_resp_bits_data_0 & 32'h3050;
  assign T19 = T46 | T20;
  assign T20 = id_reg_fence & T21;
  assign T21 = id_ctrl_mem | id_ctrl_rocc;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_mem = T22;
  assign T22 = T25 | T23;
  assign T23 = T24 == 32'h1000202f;
  assign T24 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h800202f;
  assign T27 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h202f;
  assign T30 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h3;
  assign T33 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T34 = T37 | T35;
  assign T35 = T36 == 32'h3;
  assign T36 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T37 = T38 == 32'h3;
  assign T38 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T916 = reset ? 1'h0 : T39;
  assign T39 = id_fence_next | T40;
  assign T40 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_ctrl_fence | T41;
  assign T41 = id_ctrl_amo & id_amo_rl;
  assign id_amo_rl = io_imem_resp_bits_data_0[5'h19:5'h19];
  assign id_ctrl_amo = T42;
  assign T42 = T43 == 32'h2008;
  assign T43 = io_imem_resp_bits_data_0 & 32'h6048;
  assign id_ctrl_fence = T44;
  assign T44 = T45 == 32'h8;
  assign T45 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T46 = T49 | id_ctrl_fence_i;
  assign id_ctrl_fence_i = T47;
  assign T47 = T48 == 32'h1008;
  assign T48 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T49 = id_ctrl_amo & id_amo_aq;
  assign id_amo_aq = io_imem_resp_bits_data_0[5'h1a:5'h1a];
  assign id_mem_busy = T50 | io_dmem_req_valid;
  assign T50 = io_dmem_ordered ^ 1'h1;
  assign T51 = T54 | T52;
  assign T52 = id_ctrl_mem & T53;
  assign T53 = io_dmem_req_ready ^ 1'h1;
  assign T54 = T397 | id_sboard_hazard;
  assign id_sboard_hazard = T382 | T55;
  assign T55 = T380 & T56;
  assign T56 = T61 & T57;
  assign T57 = T58 - 1'h1;
  assign T58 = 1'h1 << T59;
  assign T59 = T60 + 5'h1;
  assign T60 = id_waddr_1 - id_waddr_1;
  assign id_waddr_1 = io_imem_resp_bits_data_0[4'hb:3'h7];
  assign T61 = T62 >> id_waddr_1;
  assign T62 = R73 & T63;
  assign T63 = ~ T64;
  assign T64 = ll_wen ? T65 : 32'h0;
  assign T65 = 1'h1 << ll_waddr;
  assign ll_waddr = T66;
  assign T66 = T68 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign dmem_resp_waddr = T67[3'h5:1'h1];
  assign T67 = io_dmem_resp_bits_tag;
  assign T68 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_xpu = T69 ^ 1'h1;
  assign T69 = T70;
  assign T70 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign ll_wen = T71;
  assign T71 = T68 ? 1'h1 : T72;
  assign T72 = T634 & div_io_resp_valid;
  assign T917 = reset ? 32'h0 : T74;
  assign T74 = T379 ? T76 : T75;
  assign T75 = ll_wen ? T62 : R73;
  assign T76 = T62 | T77;
  assign T77 = T79 ? T78 : 32'h0;
  assign T78 = 1'h1 << wb_waddr;
  assign wb_waddr = wb_reg_inst[4'hb:3'h7];
  assign T79 = wb_set_sboard & wb_wen;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign T80 = T517 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign T81 = T516 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign T82 = T103 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign id_ctrl_wxd = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h0;
  assign T85 = io_imem_resp_bits_data_0 & 32'h28;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h2010;
  assign T88 = io_imem_resp_bits_data_0 & 32'h2010;
  assign T89 = T92 | T90;
  assign T90 = T91 == 32'h2008;
  assign T91 = io_imem_resp_bits_data_0 & 32'h2008;
  assign T92 = T95 | T93;
  assign T93 = T94 == 32'h1010;
  assign T94 = io_imem_resp_bits_data_0 & 32'h1010;
  assign T95 = T98 | T96;
  assign T96 = T97 == 32'h48;
  assign T97 = io_imem_resp_bits_data_0 & 32'h48;
  assign T98 = T101 | T99;
  assign T99 = T100 == 32'h10;
  assign T100 = io_imem_resp_bits_data_0 & 32'h50;
  assign T101 = T102 == 32'h4;
  assign T102 = io_imem_resp_bits_data_0 & 32'hc;
  assign T103 = ctrl_killd ^ 1'h1;
  assign wb_valid = T105 & T104;
  assign T104 = csr_io_csr_xcpt ^ 1'h1;
  assign T105 = wb_reg_valid & T106;
  assign T106 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T107;
  assign T107 = T109 & T108;
  assign T108 = io_rocc_cmd_ready ^ 1'h1;
  assign T109 = wb_reg_valid & wb_ctrl_rocc;
  assign T110 = T517 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign T111 = T516 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign T112 = T103 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign replay_wb_common = T113 | csr_io_csr_replay;
  assign T113 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T114 = replay_mem & T115;
  assign T115 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T116;
  assign T116 = T117 | csr_io_eret;
  assign T117 = replay_wb | wb_xcpt;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T118 = mem_xcpt & T119;
  assign T119 = take_pc_wb ^ 1'h1;
  assign mem_xcpt = T260 | T120;
  assign T120 = T121 & io_dmem_xcpt_pf_ld;
  assign T121 = mem_reg_valid & mem_ctrl_mem;
  assign T122 = T516 ? ex_ctrl_mem : mem_ctrl_mem;
  assign T123 = T103 ? id_ctrl_mem : ex_ctrl_mem;
  assign T124 = ctrl_killx ^ 1'h1;
  assign ctrl_killx = T127 | T125;
  assign T125 = ex_reg_valid ^ 1'h1;
  assign T126 = ctrl_killd ^ 1'h1;
  assign T127 = take_pc | replay_ex;
  assign replay_ex = ex_reg_valid & T128;
  assign T128 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T129 = T103 ? id_load_use : ex_reg_load_use;
  assign id_load_use = T130;
  assign T130 = T131 & mem_ctrl_mem;
  assign T131 = mem_reg_valid & data_hazard_mem;
  assign data_hazard_mem = mem_ctrl_wxd & T132;
  assign T132 = T135 | T133;
  assign T133 = T380 & T134;
  assign T134 = id_waddr_1 == mem_waddr;
  assign mem_waddr = mem_reg_inst[4'hb:3'h7];
  assign T135 = T148 | T136;
  assign T136 = T138 & T137;
  assign T137 = id_raddr_1 == mem_waddr;
  assign id_raddr_1 = io_imem_resp_bits_data_0[5'h18:5'h14];
  assign T138 = id_ctrl_rxs2 & T139;
  assign T139 = id_raddr_1 != 5'h0;
  assign id_ctrl_rxs2 = T140;
  assign T140 = T143 | T141;
  assign T141 = T142 == 32'h20;
  assign T142 = io_imem_resp_bits_data_0 & 32'h34;
  assign T143 = T146 | T144;
  assign T144 = T145 == 32'h20;
  assign T145 = io_imem_resp_bits_data_0 & 32'h64;
  assign T146 = T147 == 32'h20;
  assign T147 = io_imem_resp_bits_data_0 & 32'h70;
  assign T148 = T150 & T149;
  assign T149 = id_raddr_0 == mem_waddr;
  assign id_raddr_0 = io_imem_resp_bits_data_0[5'h13:4'hf];
  assign T150 = id_ctrl_rxs1 & T151;
  assign T151 = id_raddr_0 != 5'h0;
  assign id_ctrl_rxs1 = T152;
  assign T152 = T155 | T153;
  assign T153 = T154 == 32'h2000;
  assign T154 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T155 = T158 | T156;
  assign T156 = T157 == 32'h0;
  assign T157 = io_imem_resp_bits_data_0 & 32'h18;
  assign T158 = T161 | T159;
  assign T159 = T160 == 32'h0;
  assign T160 = io_imem_resp_bits_data_0 & 32'h44;
  assign T161 = T162 == 32'h0;
  assign T162 = io_imem_resp_bits_data_0 & 32'h4004;
  assign wb_dcache_miss = wb_ctrl_mem & T163;
  assign T163 = io_dmem_resp_valid ^ 1'h1;
  assign T164 = T517 ? mem_ctrl_mem : wb_ctrl_mem;
  assign replay_ex_structural = T170 | T165;
  assign T165 = ex_ctrl_div & T166;
  assign T166 = div_io_req_ready ^ 1'h1;
  assign T167 = T103 ? id_ctrl_div : ex_ctrl_div;
  assign id_ctrl_div = T168;
  assign T168 = T169 == 32'h2000030;
  assign T169 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T170 = ex_ctrl_mem & T171;
  assign T171 = io_dmem_req_ready ^ 1'h1;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = T172;
  assign T172 = want_take_pc_mem & T173;
  assign T173 = mem_npc_misaligned ^ 1'h1;
  assign mem_npc_misaligned = mem_npc[1'h1:1'h1];
  assign mem_npc = T174;
  assign T174 = T175 & 40'hfffffffffe;
  assign T175 = mem_ctrl_jalr ? T217 : mem_br_target;
  assign mem_br_target = T214 + T918;
  assign T918 = {T922, T176};
  assign T176 = T208 ? T919 : T177;
  assign T177 = mem_ctrl_jal ? T178 : 22'h4;
  assign T178 = T179;
  assign T179 = {T187, T180};
  assign T180 = {T183, T181};
  assign T181 = {T182, 1'h0};
  assign T182 = mem_reg_inst[5'h18:5'h15];
  assign T183 = {T185, T184};
  assign T184 = mem_reg_inst[5'h1e:5'h19];
  assign T185 = T186;
  assign T186 = mem_reg_inst[5'h14:5'h14];
  assign T187 = {T191, T188};
  assign T188 = {T191, T189};
  assign T189 = T190;
  assign T190 = mem_reg_inst[5'h13:4'hc];
  assign T191 = T192;
  assign T192 = mem_reg_inst[5'h1f:5'h1f];
  assign T193 = T516 ? ex_ctrl_jal : mem_ctrl_jal;
  assign T194 = T103 ? id_ctrl_jal : ex_ctrl_jal;
  assign id_ctrl_jal = T96;
  assign T919 = {T920, T195};
  assign T195 = T196;
  assign T196 = {T204, T197};
  assign T197 = {T200, T198};
  assign T198 = {T199, 1'h0};
  assign T199 = mem_reg_inst[4'hb:4'h8];
  assign T200 = {T202, T201};
  assign T201 = mem_reg_inst[5'h1e:5'h19];
  assign T202 = T203;
  assign T203 = mem_reg_inst[3'h7:3'h7];
  assign T204 = {T206, T205};
  assign T205 = {T206, T206};
  assign T206 = T207;
  assign T207 = mem_reg_inst[5'h1f:5'h1f];
  assign T920 = T921 ? 7'h7f : 7'h0;
  assign T921 = T195[4'he:4'he];
  assign T208 = mem_ctrl_branch & mem_br_taken;
  assign mem_br_taken = bypass_mux_1[1'h0:1'h0];
  assign T209 = T516 ? alu_io_out : bypass_mux_1;
  assign T210 = T516 ? ex_ctrl_branch : mem_ctrl_branch;
  assign T211 = T103 ? id_ctrl_branch : ex_ctrl_branch;
  assign id_ctrl_branch = T212;
  assign T212 = T213 == 32'h40;
  assign T213 = io_imem_resp_bits_data_0 & 32'h54;
  assign T922 = T923 ? 18'h3ffff : 18'h0;
  assign T923 = T176[5'h15:5'h15];
  assign T214 = mem_reg_pc;
  assign T215 = T516 ? ex_reg_pc : mem_reg_pc;
  assign T216 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T217 = T218;
  assign T218 = {T220, T219};
  assign T219 = bypass_mux_1[6'h26:1'h0];
  assign T220 = T233 ? T232 : T221;
  assign T221 = T226 ? T224 : T222;
  assign T222 = T223[1'h0:1'h0];
  assign T223 = bypass_mux_1[6'h27:6'h26];
  assign T224 = T225 == 2'h3;
  assign T225 = T223;
  assign T226 = T230 | T227;
  assign T227 = T228 == 26'h3fffffe;
  assign T228 = T229;
  assign T229 = bypass_mux_1 >> 6'h26;
  assign T230 = T231 == 26'h3ffffff;
  assign T231 = T229;
  assign T232 = T223 != 2'h0;
  assign T233 = T235 | T234;
  assign T234 = T229 == 26'h1;
  assign T235 = T229 == 26'h0;
  assign T236 = T516 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign T237 = T103 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign id_ctrl_jalr = T238;
  assign T238 = T239 == 32'h4;
  assign T239 = io_imem_resp_bits_data_0 & 32'h1c;
  assign want_take_pc_mem = mem_reg_valid & T240;
  assign T240 = mem_misprediction | mem_reg_flush_pipe;
  assign T241 = T516 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign T242 = T103 ? T243 : ex_reg_flush_pipe;
  assign T243 = id_ctrl_fence_i | id_csr_flush;
  assign id_csr_flush = id_system_insn | T244;
  assign T244 = T249 & T245;
  assign T245 = T246 ^ 1'h1;
  assign T246 = T247;
  assign T247 = T248 == 12'h40;
  assign T248 = id_csr_addr & 12'h8c4;
  assign id_csr_addr = io_imem_resp_bits_data_0[5'h1f:5'h14];
  assign T249 = id_csr_en & T250;
  assign T250 = id_csr_ren ^ 1'h1;
  assign id_csr_ren = T252 & T251;
  assign T251 = id_raddr_0 == 5'h0;
  assign T252 = T254 | T253;
  assign T253 = id_ctrl_csr == 3'h3;
  assign T254 = id_ctrl_csr == 3'h2;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign mem_misprediction = T257 & T255;
  assign T255 = T256 | mem_ctrl_jal;
  assign T256 = mem_ctrl_branch | mem_ctrl_jalr;
  assign T257 = mem_wrong_npc & mem_reg_valid;
  assign mem_wrong_npc = T259 | T258;
  assign T258 = ex_reg_valid ^ 1'h1;
  assign T259 = mem_npc != ex_reg_pc;
  assign T260 = T263 | T261;
  assign T261 = T262 & io_dmem_xcpt_pf_st;
  assign T262 = mem_reg_valid & mem_ctrl_mem;
  assign T263 = T266 | T264;
  assign T264 = T265 & io_dmem_xcpt_ma_ld;
  assign T265 = mem_reg_valid & mem_ctrl_mem;
  assign T266 = T269 | T267;
  assign T267 = T268 & io_dmem_xcpt_ma_st;
  assign T268 = mem_reg_valid & mem_ctrl_mem;
  assign T269 = T271 | T270;
  assign T270 = want_take_pc_mem & mem_npc_misaligned;
  assign T271 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T272 = T362 & ex_xcpt;
  assign ex_xcpt = T275 | T273;
  assign T273 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign T274 = T103 ? id_ctrl_fp : ex_ctrl_fp;
  assign id_ctrl_fp = 1'h0;
  assign T275 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T276 = T358 & id_xcpt;
  assign id_xcpt = T357 | id_illegal_insn;
  assign id_illegal_insn = T280 | T277;
  assign T277 = id_ctrl_rocc & T278;
  assign T278 = T279 ^ 1'h1;
  assign T279 = csr_io_status_xs != 2'h0;
  assign T280 = T284 | T281;
  assign T281 = id_ctrl_fp & T282;
  assign T282 = T283 ^ 1'h1;
  assign T283 = csr_io_status_fs != 2'h0;
  assign T284 = id_ctrl_legal ^ 1'h1;
  assign id_ctrl_legal = T285;
  assign T285 = T288 | T286;
  assign T286 = T287 == 32'h33;
  assign T287 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T288 = T291 | T289;
  assign T289 = T290 == 32'h4063;
  assign T290 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T291 = T294 | T292;
  assign T292 = T293 == 32'h1063;
  assign T293 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T294 = T296 | T295;
  assign T295 = io_imem_resp_bits_data_0 == 32'h30500073;
  assign T296 = T299 | T297;
  assign T297 = T298 == 32'h10100073;
  assign T298 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T299 = T300 | T23;
  assign T300 = T303 | T301;
  assign T301 = T302 == 32'h10000073;
  assign T302 = io_imem_resp_bits_data_0 & 32'hffdfffff;
  assign T303 = T304 | T26;
  assign T304 = T307 | T305;
  assign T305 = T306 == 32'h2004033;
  assign T306 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T307 = T310 | T308;
  assign T308 = T309 == 32'h5033;
  assign T309 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T310 = T313 | T311;
  assign T311 = T312 == 32'h501b;
  assign T312 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T313 = T316 | T314;
  assign T314 = T315 == 32'h5013;
  assign T315 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T316 = T319 | T317;
  assign T317 = T318 == 32'h2073;
  assign T318 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T319 = T320 | T29;
  assign T320 = T323 | T321;
  assign T321 = T322 == 32'h2013;
  assign T322 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T323 = T326 | T324;
  assign T324 = T325 == 32'h101b;
  assign T325 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T326 = T329 | T327;
  assign T327 = T328 == 32'h1013;
  assign T328 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T329 = T332 | T330;
  assign T330 = T331 == 32'h73;
  assign T331 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T332 = T335 | T333;
  assign T333 = T334 == 32'h6f;
  assign T334 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T335 = T338 | T336;
  assign T336 = T337 == 32'h63;
  assign T337 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T338 = T341 | T339;
  assign T339 = T340 == 32'h33;
  assign T340 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T341 = T344 | T342;
  assign T342 = T343 == 32'h33;
  assign T343 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T344 = T347 | T345;
  assign T345 = T346 == 32'h17;
  assign T346 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T347 = T350 | T348;
  assign T348 = T349 == 32'h13;
  assign T349 = io_imem_resp_bits_data_0 & 32'h7077;
  assign T350 = T353 | T351;
  assign T351 = T352 == 32'hf;
  assign T352 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T353 = T356 | T354;
  assign T354 = T355 == 32'h3;
  assign T355 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T356 = T37 | T35;
  assign T357 = csr_io_interrupt | io_imem_resp_bits_xcpt_if;
  assign T358 = ctrl_killd ^ 1'h1;
  assign T359 = T360 & io_imem_resp_valid;
  assign T360 = csr_io_interrupt & T361;
  assign T361 = take_pc ^ 1'h1;
  assign T362 = ctrl_killx ^ 1'h1;
  assign T363 = T364 & ex_reg_xcpt_interrupt;
  assign T364 = take_pc ^ 1'h1;
  assign replay_mem = T367 | fpu_kill_mem;
  assign fpu_kill_mem = T365 & io_fpu_nack_mem;
  assign T365 = mem_reg_valid & mem_ctrl_fp;
  assign T366 = T516 ? ex_ctrl_fp : mem_ctrl_fp;
  assign T367 = dcache_kill_mem | mem_reg_replay;
  assign T368 = T369 & replay_ex;
  assign T369 = take_pc ^ 1'h1;
  assign dcache_kill_mem = T370 & io_dmem_replay_next_valid;
  assign T370 = mem_reg_valid & mem_ctrl_wxd;
  assign T371 = ctrl_killm ^ 1'h1;
  assign ctrl_killm = T372 | fpu_kill_mem;
  assign T372 = killm_common | mem_xcpt;
  assign killm_common = T374 | T373;
  assign T373 = mem_reg_valid ^ 1'h1;
  assign T374 = T375 | mem_reg_xcpt;
  assign T375 = dcache_kill_mem | take_pc_wb;
  assign wb_set_sboard = T376 | wb_ctrl_rocc;
  assign T376 = wb_ctrl_div | wb_dcache_miss;
  assign T377 = T517 ? mem_ctrl_div : wb_ctrl_div;
  assign T378 = T516 ? ex_ctrl_div : mem_ctrl_div;
  assign T379 = ll_wen | T79;
  assign T380 = id_ctrl_wxd & T381;
  assign T381 = id_waddr_1 != 5'h0;
  assign T382 = T390 | T383;
  assign T383 = T138 & T384;
  assign T384 = T389 & T385;
  assign T385 = T386 - 1'h1;
  assign T386 = 1'h1 << T387;
  assign T387 = T388 + 5'h1;
  assign T388 = id_raddr_1 - id_raddr_1;
  assign T389 = T62 >> id_raddr_1;
  assign T390 = T150 & T391;
  assign T391 = T396 & T392;
  assign T392 = T393 - 1'h1;
  assign T393 = 1'h1 << T394;
  assign T394 = T395 + 5'h1;
  assign T395 = id_raddr_0 - id_raddr_0;
  assign T396 = T62 >> id_raddr_0;
  assign T397 = T422 | id_wb_hazard;
  assign id_wb_hazard = wb_reg_valid & T398;
  assign T398 = T413 | fp_data_hazard_wb;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T399;
  assign T399 = T402 | T400;
  assign T400 = io_fpu_dec_wen & T401;
  assign T401 = id_waddr_1 == wb_waddr;
  assign T402 = T405 | T403;
  assign T403 = io_fpu_dec_ren3 & T404;
  assign T404 = id_raddr3 == wb_waddr;
  assign id_raddr3 = io_imem_resp_bits_data_0[5'h1f:5'h1b];
  assign T405 = T408 | T406;
  assign T406 = io_fpu_dec_ren2 & T407;
  assign T407 = id_raddr_1 == wb_waddr;
  assign T408 = io_fpu_dec_ren1 & T409;
  assign T409 = id_raddr_0 == wb_waddr;
  assign T410 = T517 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign T411 = T516 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign T412 = T103 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign id_ctrl_wfd = 1'h0;
  assign T413 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_ctrl_wxd & T414;
  assign T414 = T417 | T415;
  assign T415 = T380 & T416;
  assign T416 = id_waddr_1 == wb_waddr;
  assign T417 = T420 | T418;
  assign T418 = T138 & T419;
  assign T419 = id_raddr_1 == wb_waddr;
  assign T420 = T150 & T421;
  assign T421 = id_raddr_0 == wb_waddr;
  assign T422 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = mem_reg_valid & T423;
  assign T423 = T435 | fp_data_hazard_mem;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T424;
  assign T424 = T427 | T425;
  assign T425 = io_fpu_dec_wen & T426;
  assign T426 = id_waddr_1 == mem_waddr;
  assign T427 = T430 | T428;
  assign T428 = io_fpu_dec_ren3 & T429;
  assign T429 = id_raddr3 == mem_waddr;
  assign T430 = T433 | T431;
  assign T431 = io_fpu_dec_ren2 & T432;
  assign T432 = id_raddr_1 == mem_waddr;
  assign T433 = io_fpu_dec_ren1 & T434;
  assign T434 = id_raddr_0 == mem_waddr;
  assign T435 = data_hazard_mem & mem_cannot_bypass;
  assign mem_cannot_bypass = T436 | mem_ctrl_rocc;
  assign T436 = T437 | mem_ctrl_fp;
  assign T437 = T438 | mem_ctrl_div;
  assign T438 = T484 | T439;
  assign T439 = mem_ctrl_mem & mem_mem_cmd_bh;
  assign T440 = T516 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T457 | T441;
  assign T441 = T452 | T442;
  assign T442 = 3'h5 == ex_ctrl_mem_type;
  assign T443 = T103 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign id_ctrl_mem_type = T444;
  assign T444 = {T450, T445};
  assign T445 = {T448, T446};
  assign T446 = T447 == 32'h1000;
  assign T447 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T448 = T449 == 32'h2000;
  assign T449 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T450 = T451 == 32'h4000;
  assign T451 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T452 = T454 | T453;
  assign T453 = 3'h1 == ex_ctrl_mem_type;
  assign T454 = T456 | T455;
  assign T455 = 3'h4 == ex_ctrl_mem_type;
  assign T456 = 3'h0 == ex_ctrl_mem_type;
  assign T457 = ex_ctrl_mem_cmd == 5'h7;
  assign T458 = T103 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign id_ctrl_mem_cmd = T459;
  assign T459 = {1'h0, T460};
  assign T460 = {T482, T461};
  assign T461 = {T476, T462};
  assign T462 = {T471, T463};
  assign T463 = T466 | T464;
  assign T464 = T465 == 32'h20000020;
  assign T465 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T466 = T469 | T467;
  assign T467 = T468 == 32'h18000020;
  assign T468 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T469 = T470 == 32'h20;
  assign T470 = io_imem_resp_bits_data_0 & 32'h28;
  assign T471 = T474 | T472;
  assign T472 = T473 == 32'h40000008;
  assign T473 = io_imem_resp_bits_data_0 & 32'h40000008;
  assign T474 = T475 == 32'h10000008;
  assign T475 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T476 = T479 | T477;
  assign T477 = T478 == 32'h80000008;
  assign T478 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T479 = T480 | T474;
  assign T480 = T481 == 32'h8000008;
  assign T481 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T482 = T483 == 32'h8;
  assign T483 = io_imem_resp_bits_data_0 & 32'h18000008;
  assign T484 = mem_ctrl_csr != 3'h0;
  assign T485 = T516 ? ex_ctrl_csr : mem_ctrl_csr;
  assign T486 = T103 ? id_csr : T487;
  assign T487 = T103 ? id_ctrl_csr : ex_ctrl_csr;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_ex_hazard = ex_reg_valid & T488;
  assign T488 = T500 | fp_data_hazard_ex;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T489;
  assign T489 = T492 | T490;
  assign T490 = io_fpu_dec_wen & T491;
  assign T491 = id_waddr_1 == ex_waddr;
  assign ex_waddr = ex_reg_inst[4'hb:3'h7];
  assign T492 = T495 | T493;
  assign T493 = io_fpu_dec_ren3 & T494;
  assign T494 = id_raddr3 == ex_waddr;
  assign T495 = T498 | T496;
  assign T496 = io_fpu_dec_ren2 & T497;
  assign T497 = id_raddr_1 == ex_waddr;
  assign T498 = io_fpu_dec_ren1 & T499;
  assign T499 = id_raddr_0 == ex_waddr;
  assign T500 = data_hazard_ex & ex_cannot_bypass;
  assign ex_cannot_bypass = T501 | ex_ctrl_rocc;
  assign T501 = T502 | ex_ctrl_fp;
  assign T502 = T503 | ex_ctrl_div;
  assign T503 = T504 | ex_ctrl_mem;
  assign T504 = T505 | ex_ctrl_jalr;
  assign T505 = ex_ctrl_csr != 3'h0;
  assign data_hazard_ex = ex_ctrl_wxd & T506;
  assign T506 = T509 | T507;
  assign T507 = T380 & T508;
  assign T508 = id_waddr_1 == ex_waddr;
  assign T509 = T512 | T510;
  assign T510 = T138 & T511;
  assign T511 = id_raddr_1 == ex_waddr;
  assign T512 = T150 & T513;
  assign T513 = id_raddr_0 == ex_waddr;
  assign T514 = T515 | take_pc;
  assign T515 = io_imem_resp_valid ^ 1'h1;
  assign T516 = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T517 = T518 | mem_reg_xcpt_interrupt;
  assign T518 = mem_reg_valid | mem_reg_replay;
  assign T519 = wb_reg_inst;
  assign T520 = R521;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T573 : T523;
  assign T523 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T524 = T562 ? T538 : T525;
  assign T525 = T103 ? T526 : ex_reg_rs_lsb_1;
  assign T526 = T537 ? 2'h0 : T527;
  assign T527 = T534 ? 2'h1 : T528;
  assign T528 = T529 ? 2'h2 : 2'h3;
  assign T529 = T531 & T530;
  assign T530 = mem_waddr == id_raddr_1;
  assign T531 = T533 & T532;
  assign T532 = mem_ctrl_mem ^ 1'h1;
  assign T533 = mem_reg_valid & mem_ctrl_wxd;
  assign T534 = T536 & T535;
  assign T535 = ex_waddr == id_raddr_1;
  assign T536 = ex_reg_valid & ex_ctrl_wxd;
  assign T537 = 5'h0 == id_raddr_1;
  assign T538 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T539;
  assign T539 = T560 ? rf_wdata : T540;
  assign T540 = T541[T549];
  assign T543 = T546 & T544;
  assign T544 = T545 < 5'h1f;
  assign T545 = T548[3'h4:1'h0];
  assign T546 = rf_wen & T547;
  assign T547 = rf_waddr != 5'h0;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign rf_wen = wb_wen | ll_wen;
  assign T548 = ~ rf_waddr;
  assign T549 = ~ id_raddr_1;
  assign rf_wdata = T559 ? io_dmem_resp_bits_data_subword : T550;
  assign T550 = ll_wen ? ll_wdata : T551;
  assign T551 = T557 ? csr_io_rw_rdata : bypass_mux_2;
  assign T552 = T517 ? T553 : bypass_mux_2;
  assign T553 = T556 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = T554;
  assign T554 = mem_ctrl_jalr ? T924 : T555;
  assign T555 = bypass_mux_1;
  assign T924 = {T925, mem_br_target};
  assign T925 = T926 ? 24'hffffff : 24'h0;
  assign T926 = mem_br_target[6'h27:6'h27];
  assign T556 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T557 = wb_ctrl_csr != 3'h0;
  assign T558 = T517 ? mem_ctrl_csr : wb_ctrl_csr;
  assign ll_wdata = div_io_resp_bits_data;
  assign T559 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T560 = T546 & T561;
  assign T561 = rf_waddr == id_raddr_1;
  assign T562 = T103 & T563;
  assign T563 = id_ctrl_rxs2 & T564;
  assign T564 = T565 ^ 1'h1;
  assign T565 = T569 | T566;
  assign T566 = T568 & T567;
  assign T567 = mem_waddr == id_raddr_1;
  assign T568 = mem_reg_valid & mem_ctrl_wxd;
  assign T569 = T570 | T529;
  assign T570 = T537 | T534;
  assign T571 = T562 ? T572 : ex_reg_rs_msb_1;
  assign T572 = id_rs_1 >> 2'h2;
  assign T573 = T579 ? T577 : T574;
  assign T574 = T575 ? bypass_mux_1 : 64'h0;
  assign T575 = T576[1'h0:1'h0];
  assign T576 = ex_reg_rs_lsb_1;
  assign T577 = T578 ? io_dmem_resp_bits_data : bypass_mux_2;
  assign T578 = T576[1'h0:1'h0];
  assign T579 = T576[1'h1:1'h1];
  assign T580 = T103 ? T565 : ex_reg_rs_bypass_1;
  assign T581 = T582;
  assign T582 = wb_reg_inst[5'h18:5'h14];
  assign T583 = R584;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T613 : T586;
  assign T586 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T587 = T603 ? T597 : T588;
  assign T588 = T103 ? T589 : ex_reg_rs_lsb_0;
  assign T589 = T596 ? 2'h0 : T590;
  assign T590 = T594 ? 2'h1 : T591;
  assign T591 = T592 ? 2'h2 : 2'h3;
  assign T592 = T531 & T593;
  assign T593 = mem_waddr == id_raddr_0;
  assign T594 = T536 & T595;
  assign T595 = ex_waddr == id_raddr_0;
  assign T596 = 5'h0 == id_raddr_0;
  assign T597 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T598;
  assign T598 = T601 ? rf_wdata : T599;
  assign T599 = T541[T600];
  assign T600 = ~ id_raddr_0;
  assign T601 = T546 & T602;
  assign T602 = rf_waddr == id_raddr_0;
  assign T603 = T103 & T604;
  assign T604 = id_ctrl_rxs1 & T605;
  assign T605 = T606 ^ 1'h1;
  assign T606 = T609 | T607;
  assign T607 = T568 & T608;
  assign T608 = mem_waddr == id_raddr_0;
  assign T609 = T610 | T592;
  assign T610 = T596 | T594;
  assign T611 = T603 ? T612 : ex_reg_rs_msb_0;
  assign T612 = id_rs_0 >> 2'h2;
  assign T613 = T619 ? T617 : T614;
  assign T614 = T615 ? bypass_mux_1 : 64'h0;
  assign T615 = T616[1'h0:1'h0];
  assign T616 = ex_reg_rs_lsb_0;
  assign T617 = T618 ? io_dmem_resp_bits_data : bypass_mux_2;
  assign T618 = T616[1'h0:1'h0];
  assign T619 = T616[1'h1:1'h1];
  assign T620 = T103 ? T606 : ex_reg_rs_bypass_0;
  assign T621 = T622;
  assign T622 = wb_reg_inst[5'h13:4'hf];
  assign T623 = rf_wen;
  assign T624 = rf_wdata;
  assign T625 = T626;
  assign T626 = rf_wen ? rf_waddr : 5'h0;
  assign T627 = wb_reg_pc;
  assign T628 = T517 ? mem_reg_pc : wb_reg_pc;
  assign T629 = wb_valid;
  assign T630 = T631;
  assign T631 = csr_io_time[6'h20:1'h0];
  assign T632 = io_host_id;
  assign T634 = T68 ? 1'h0 : T635;
  assign T635 = T636 ^ 1'h1;
  assign T636 = wb_reg_valid & wb_ctrl_wxd;
  assign T637 = killm_common & R638;
  assign T639 = div_io_req_ready & T690;
  assign T640 = T103 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign id_ctrl_alu_dw = T641;
  assign T641 = T644 | T642;
  assign T642 = T643 == 32'h0;
  assign T643 = io_imem_resp_bits_data_0 & 32'h8;
  assign T644 = T645 == 32'h0;
  assign T645 = io_imem_resp_bits_data_0 & 32'h10;
  assign T646 = T103 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign id_ctrl_alu_fn = T647;
  assign T647 = {T683, T648};
  assign T648 = {T672, T649};
  assign T649 = {T658, T650};
  assign T650 = T653 | T651;
  assign T651 = T652 == 32'h7000;
  assign T652 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T653 = T656 | T654;
  assign T654 = T655 == 32'h1040;
  assign T655 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T656 = T657 == 32'h1010;
  assign T657 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T658 = T661 | T659;
  assign T659 = T660 == 32'h40001010;
  assign T660 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T661 = T664 | T662;
  assign T662 = T663 == 32'h40000030;
  assign T663 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T664 = T667 | T665;
  assign T665 = T666 == 32'h6010;
  assign T666 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T667 = T670 | T668;
  assign T668 = T669 == 32'h3010;
  assign T669 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T670 = T671 == 32'h2040;
  assign T671 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T672 = T675 | T673;
  assign T673 = T674 == 32'h4040;
  assign T674 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T675 = T678 | T676;
  assign T676 = T677 == 32'h4010;
  assign T677 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T678 = T681 | T679;
  assign T679 = T680 == 32'h4010;
  assign T680 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T681 = T682 == 32'h2010;
  assign T682 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T683 = T686 | T684;
  assign T684 = T685 == 32'h40001010;
  assign T685 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T686 = T687 | T662;
  assign T687 = T212 | T688;
  assign T688 = T689 == 32'h2010;
  assign T689 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T690 = ex_reg_valid & ex_ctrl_div;
  assign T691 = ex_op1;
  assign ex_op1 = T706 ? T705 : T927;
  assign T927 = {T928, T692};
  assign T692 = T694 ? T693 : 40'h0;
  assign T693 = ex_reg_pc;
  assign T694 = ex_ctrl_sel_alu1 == 2'h2;
  assign T695 = T103 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign id_ctrl_sel_alu1 = T696;
  assign T696 = {T702, T697};
  assign T697 = T698 | T156;
  assign T698 = T699 | T159;
  assign T699 = T161 | T700;
  assign T700 = T701 == 32'h0;
  assign T701 = io_imem_resp_bits_data_0 & 32'h50;
  assign T702 = T703 | T96;
  assign T703 = T704 == 32'h4;
  assign T704 = io_imem_resp_bits_data_0 & 32'h24;
  assign T928 = T929 ? 24'hffffff : 24'h0;
  assign T929 = T692[6'h27:6'h27];
  assign T705 = ex_rs_0;
  assign T706 = ex_ctrl_sel_alu1 == 2'h1;
  assign T707 = ex_op2;
  assign ex_op2 = T806 ? T805 : T930;
  assign T930 = {T936, T708};
  assign T708 = T804 ? ex_imm : T931;
  assign T931 = {T932, T709};
  assign T709 = T710 ? 4'h4 : 4'h0;
  assign T710 = ex_ctrl_sel_alu2 == 2'h1;
  assign T711 = T103 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign id_ctrl_sel_alu2 = T712;
  assign T712 = {T723, T713};
  assign T713 = T716 | T714;
  assign T714 = T715 == 32'h4050;
  assign T715 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T716 = T717 | T96;
  assign T717 = T718 | T101;
  assign T718 = T721 | T719;
  assign T719 = T720 == 32'h0;
  assign T720 = io_imem_resp_bits_data_0 & 32'h20;
  assign T721 = T722 == 32'h0;
  assign T722 = io_imem_resp_bits_data_0 & 32'h58;
  assign T723 = T726 | T724;
  assign T724 = T725 == 32'h4000;
  assign T725 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T726 = T727 | T156;
  assign T727 = T728 | T159;
  assign T728 = T729 == 32'h0;
  assign T729 = io_imem_resp_bits_data_0 & 32'h48;
  assign T932 = T933 ? 28'hfffffff : 28'h0;
  assign T933 = T709[2'h3:2'h3];
  assign ex_imm = T730;
  assign T730 = {T792, T731};
  assign T731 = {T770, T732};
  assign T732 = {T759, T733};
  assign T733 = T758 ? T757 : T734;
  assign T734 = T756 ? T755 : T735;
  assign T735 = T737 ? T736 : 1'h0;
  assign T736 = ex_reg_inst[4'hf:4'hf];
  assign T737 = ex_ctrl_sel_imm == 3'h5;
  assign T738 = T103 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign id_ctrl_sel_imm = T739;
  assign T739 = {T749, T740};
  assign T740 = {T746, T741};
  assign T741 = T744 | T742;
  assign T742 = T743 == 32'h40;
  assign T743 = io_imem_resp_bits_data_0 & 32'h44;
  assign T744 = T745 == 32'h8;
  assign T745 = io_imem_resp_bits_data_0 & 32'h18;
  assign T746 = T747 | T744;
  assign T747 = T748 == 32'h4;
  assign T748 = io_imem_resp_bits_data_0 & 32'h44;
  assign T749 = T752 | T750;
  assign T750 = T751 == 32'h10;
  assign T751 = io_imem_resp_bits_data_0 & 32'h14;
  assign T752 = T753 | T238;
  assign T753 = T754 == 32'h0;
  assign T754 = io_imem_resp_bits_data_0 & 32'h24;
  assign T755 = ex_reg_inst[5'h14:5'h14];
  assign T756 = ex_ctrl_sel_imm == 3'h4;
  assign T757 = ex_reg_inst[3'h7:3'h7];
  assign T758 = ex_ctrl_sel_imm == 3'h0;
  assign T759 = T769 ? 4'h0 : T760;
  assign T760 = T766 ? T765 : T761;
  assign T761 = T764 ? T763 : T762;
  assign T762 = ex_reg_inst[5'h18:5'h15];
  assign T763 = ex_reg_inst[5'h13:5'h10];
  assign T764 = ex_ctrl_sel_imm == 3'h5;
  assign T765 = ex_reg_inst[4'hb:4'h8];
  assign T766 = T768 | T767;
  assign T767 = ex_ctrl_sel_imm == 3'h1;
  assign T768 = ex_ctrl_sel_imm == 3'h0;
  assign T769 = ex_ctrl_sel_imm == 3'h2;
  assign T770 = {T776, T771};
  assign T771 = T773 ? 6'h0 : T772;
  assign T772 = ex_reg_inst[5'h1e:5'h19];
  assign T773 = T775 | T774;
  assign T774 = ex_ctrl_sel_imm == 3'h5;
  assign T775 = ex_ctrl_sel_imm == 3'h2;
  assign T776 = T789 ? 1'h0 : T777;
  assign T777 = T788 ? T786 : T778;
  assign T778 = T785 ? T783 : T779;
  assign T779 = T782 ? 1'h0 : T780;
  assign T780 = T781;
  assign T781 = ex_reg_inst[5'h1f:5'h1f];
  assign T782 = ex_ctrl_sel_imm == 3'h5;
  assign T783 = T784;
  assign T784 = ex_reg_inst[3'h7:3'h7];
  assign T785 = ex_ctrl_sel_imm == 3'h1;
  assign T786 = T787;
  assign T787 = ex_reg_inst[5'h14:5'h14];
  assign T788 = ex_ctrl_sel_imm == 3'h3;
  assign T789 = T791 | T790;
  assign T790 = ex_ctrl_sel_imm == 3'h5;
  assign T791 = ex_ctrl_sel_imm == 3'h2;
  assign T792 = {T779, T793};
  assign T793 = {T800, T794};
  assign T794 = T797 ? T934 : T795;
  assign T795 = T796;
  assign T796 = ex_reg_inst[5'h13:4'hc];
  assign T934 = T779 ? 8'hff : 8'h0;
  assign T797 = T799 & T798;
  assign T798 = ex_ctrl_sel_imm != 3'h3;
  assign T799 = ex_ctrl_sel_imm != 3'h2;
  assign T800 = T803 ? T801 : T935;
  assign T935 = T779 ? 11'h7ff : 11'h0;
  assign T801 = T802;
  assign T802 = ex_reg_inst[5'h1e:5'h14];
  assign T803 = ex_ctrl_sel_imm == 3'h2;
  assign T804 = ex_ctrl_sel_alu2 == 2'h3;
  assign T936 = T937 ? 32'hffffffff : 32'h0;
  assign T937 = T708[5'h1f:5'h1f];
  assign T805 = ex_rs_1;
  assign T806 = ex_ctrl_sel_alu2 == 2'h2;
  assign T807 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T271 ? mem_reg_cause : T938;
  assign T938 = {61'h0, T808};
  assign T808 = T270 ? 3'h0 : T809;
  assign T809 = T267 ? 3'h6 : T810;
  assign T810 = T264 ? 3'h4 : T811;
  assign T811 = T261 ? 3'h7 : 3'h5;
  assign T812 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T275 ? ex_reg_cause : 64'h2;
  assign T813 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : T939;
  assign T939 = {62'h0, T814};
  assign T814 = io_imem_resp_bits_xcpt_if ? 2'h1 : 2'h2;
  assign T815 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T816 = wb_reg_inst[5'h1f:5'h14];
  assign io_rocc_exception = T817;
  assign T817 = wb_xcpt & T818;
  assign T818 = csr_io_status_xs != 2'h0;
  assign io_rocc_s = T819;
  assign T819 = csr_io_status_prv != 2'h0;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T820 = T826 ? mem_reg_rs2 : wb_reg_rs2;
  assign T821 = T822 ? ex_rs_1 : mem_reg_rs2;
  assign T822 = T516 & T823;
  assign T823 = ex_ctrl_rxs2 & T824;
  assign T824 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T825 = T103 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign T826 = T517 & mem_ctrl_rocc;
  assign io_rocc_cmd_bits_rs1 = bypass_mux_2;
  assign io_rocc_cmd_bits_inst_opcode = T827;
  assign T827 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T828;
  assign T828 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T829;
  assign T829 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T830;
  assign T830 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T831;
  assign T831 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T832;
  assign T832 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T833;
  assign T833 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T834;
  assign T834 = wb_reg_inst[5'h1f:5'h19];
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = T836 & T835;
  assign T835 = replay_wb_common ^ 1'h1;
  assign T836 = wb_reg_valid & wb_ctrl_rocc;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T837;
  assign T837 = T838 & id_ctrl_fp;
  assign T838 = ctrl_killd ^ 1'h1;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T839;
  assign T839 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T840;
  assign T840 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_ptw_status_ie = csr_io_status_ie;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_ie1 = csr_io_status_ie1;
  assign io_ptw_status_prv1 = csr_io_status_prv1;
  assign io_ptw_status_ie2 = csr_io_status_ie2;
  assign io_ptw_status_prv2 = csr_io_status_prv2;
  assign io_ptw_status_ie3 = csr_io_status_ie3;
  assign io_ptw_status_prv3 = csr_io_status_prv3;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_ptbr = csr_io_ptbr;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_dmem_req_bits_data = T841;
  assign T841 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_kill = T842;
  assign T842 = killm_common | mem_xcpt;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_tag = T940;
  assign T940 = {2'h0, T843};
  assign T843 = {ex_waddr, ex_ctrl_fp};
  assign io_dmem_req_bits_addr = T844;
  assign T844 = T845;
  assign T845 = {T847, T846};
  assign T846 = alu_io_adder_out[6'h26:1'h0];
  assign T847 = T860 ? T859 : T848;
  assign T848 = T853 ? T851 : T849;
  assign T849 = T850[1'h0:1'h0];
  assign T850 = alu_io_adder_out[6'h27:6'h26];
  assign T851 = T852 == 2'h3;
  assign T852 = T850;
  assign T853 = T857 | T854;
  assign T854 = T855 == 26'h3fffffe;
  assign T855 = T856;
  assign T856 = ex_rs_0 >> 6'h26;
  assign T857 = T858 == 26'h3ffffff;
  assign T858 = T856;
  assign T859 = T850 != 2'h0;
  assign T860 = T862 | T861;
  assign T861 = T856 == 26'h1;
  assign T862 = T856 == 26'h0;
  assign io_dmem_req_valid = T863;
  assign T863 = ex_reg_valid & ex_ctrl_mem;
  assign io_imem_invalidate = T864;
  assign T864 = wb_reg_valid & wb_ctrl_fence_i;
  assign T865 = T517 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign T866 = T516 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign T867 = T103 ? id_ctrl_fence_i : ex_ctrl_fence_i;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_returnAddr = T941;
  assign T941 = mem_int_wdata[6'h26:1'h0];
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_isCall = T868;
  assign T868 = mem_ctrl_wxd & T869;
  assign T869 = mem_waddr[1'h0:1'h0];
  assign io_imem_ras_update_valid = T870;
  assign T870 = T872 & T871;
  assign T871 = take_pc_wb ^ 1'h1;
  assign T872 = T874 & T873;
  assign T873 = mem_npc_misaligned ^ 1'h1;
  assign T874 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_pc = T942;
  assign T942 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_valid = T875;
  assign T875 = T877 & T876;
  assign T876 = take_pc_wb ^ 1'h1;
  assign T877 = mem_reg_valid & mem_ctrl_branch;
  assign io_imem_btb_update_bits_br_pc = T943;
  assign T943 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_isReturn = T878;
  assign T878 = mem_ctrl_jalr & T879;
  assign T879 = 5'h1 == T880;
  assign T880 = T881 & 5'h19;
  assign T881 = mem_reg_inst[5'h13:4'hf];
  assign io_imem_btb_update_bits_isJump = T882;
  assign T882 = mem_ctrl_jal | mem_ctrl_jalr;
  assign io_imem_btb_update_bits_target = T944;
  assign T944 = io_imem_req_bits_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_pc = T945;
  assign T945 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T883 = T886 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T884 = T885 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T885 = T103 & io_imem_btb_resp_valid;
  assign T886 = T516 & ex_reg_btb_hit;
  assign T887 = T103 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T888 = T886 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T889 = T885 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T890 = T886 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T891 = T885 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T892 = T886 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T893 = T885 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign T894 = T886 ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign T895 = T885 ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign T896 = T886 ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign T897 = T885 ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T898 = T886 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T899 = T885 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T900 = T516 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T901;
  assign T901 = T903 & T902;
  assign T902 = take_pc_wb ^ 1'h1;
  assign T903 = T907 & T904;
  assign T904 = T905 | mem_ctrl_jal;
  assign T905 = T906 | mem_ctrl_jalr;
  assign T906 = mem_ctrl_branch & mem_br_taken;
  assign T907 = T908 & mem_wrong_npc;
  assign T908 = mem_reg_valid & T909;
  assign T909 = mem_npc_misaligned ^ 1'h1;
  assign io_imem_resp_ready = T910;
  assign T910 = T911 | csr_io_interrupt;
  assign T911 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_bits_pc = T912;
  assign T912 = T913;
  assign T913 = T915 ? csr_io_evec : T914;
  assign T914 = replay_wb ? wb_reg_pc : mem_npc;
  assign T915 = wb_xcpt | csr_io_eret;
  assign io_imem_req_valid = take_pc;
  assign io_host_debug_stats_pcr = csr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = csr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = csr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = csr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = csr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = csr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = csr_io_host_pcr_req_ready;
  CSRFile csr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( csr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( csr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( csr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( csr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( csr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( csr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( csr_io_host_debug_stats_pcr ),
       .io_rw_addr( T816 ),
       .io_rw_cmd( T815 ),
       .io_rw_rdata( csr_io_rw_rdata ),
       .io_rw_wdata( bypass_mux_2 ),
       .io_csr_replay( csr_io_csr_replay ),
       .io_csr_stall( csr_io_csr_stall ),
       .io_csr_xcpt( csr_io_csr_xcpt ),
       .io_eret( csr_io_eret ),
       .io_status_sd( csr_io_status_sd ),
       .io_status_zero2( csr_io_status_zero2 ),
       .io_status_sd_rv32( csr_io_status_sd_rv32 ),
       .io_status_zero1( csr_io_status_zero1 ),
       .io_status_vm( csr_io_status_vm ),
       .io_status_mprv( csr_io_status_mprv ),
       .io_status_xs( csr_io_status_xs ),
       .io_status_fs( csr_io_status_fs ),
       .io_status_prv3( csr_io_status_prv3 ),
       .io_status_ie3( csr_io_status_ie3 ),
       .io_status_prv2( csr_io_status_prv2 ),
       .io_status_ie2( csr_io_status_ie2 ),
       .io_status_prv1( csr_io_status_prv1 ),
       .io_status_ie1( csr_io_status_ie1 ),
       .io_status_prv( csr_io_status_prv ),
       .io_status_ie( csr_io_status_ie ),
       .io_ptbr( csr_io_ptbr ),
       .io_evec( csr_io_evec ),
       .io_exception( wb_reg_xcpt ),
       .io_retire( wb_valid ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( wb_reg_cause ),
       .io_pc( wb_reg_pc ),
       .io_fatc( csr_io_fatc ),
       .io_time( csr_io_time ),
       .io_fcsr_rm( csr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_invalidate_lr( io_rocc_mem_invalidate_lr ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_addr_block( io_rocc_imem_acquire_bits_addr_block ),
       .io_rocc_imem_acquire_bits_client_xact_id( io_rocc_imem_acquire_bits_client_xact_id ),
       .io_rocc_imem_acquire_bits_addr_beat( io_rocc_imem_acquire_bits_addr_beat ),
       .io_rocc_imem_acquire_bits_data( io_rocc_imem_acquire_bits_data ),
       .io_rocc_imem_acquire_bits_is_builtin_type( io_rocc_imem_acquire_bits_is_builtin_type ),
       .io_rocc_imem_acquire_bits_a_type( io_rocc_imem_acquire_bits_a_type ),
       .io_rocc_imem_acquire_bits_union( io_rocc_imem_acquire_bits_union ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_addr_beat(  )
       //.io_rocc_imem_grant_bits_data(  )
       //.io_rocc_imem_grant_bits_client_xact_id(  )
       //.io_rocc_imem_grant_bits_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_is_builtin_type(  )
       //.io_rocc_imem_grant_bits_g_type(  )
       //.io_rocc_dmem_acquire_ready(  )
       .io_rocc_dmem_acquire_valid( io_rocc_dmem_acquire_valid ),
       .io_rocc_dmem_acquire_bits_addr_block( io_rocc_dmem_acquire_bits_addr_block ),
       .io_rocc_dmem_acquire_bits_client_xact_id( io_rocc_dmem_acquire_bits_client_xact_id ),
       .io_rocc_dmem_acquire_bits_addr_beat( io_rocc_dmem_acquire_bits_addr_beat ),
       .io_rocc_dmem_acquire_bits_data( io_rocc_dmem_acquire_bits_data ),
       .io_rocc_dmem_acquire_bits_is_builtin_type( io_rocc_dmem_acquire_bits_is_builtin_type ),
       .io_rocc_dmem_acquire_bits_a_type( io_rocc_dmem_acquire_bits_a_type ),
       .io_rocc_dmem_acquire_bits_union( io_rocc_dmem_acquire_bits_union ),
       .io_rocc_dmem_grant_ready( io_rocc_dmem_grant_ready ),
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_addr_beat(  )
       //.io_rocc_dmem_grant_bits_data(  )
       //.io_rocc_dmem_grant_bits_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_is_builtin_type(  )
       //.io_rocc_dmem_grant_bits_g_type(  )
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits_addr( io_rocc_iptw_req_bits_addr ),
       .io_rocc_iptw_req_bits_prv( io_rocc_iptw_req_bits_prv ),
       .io_rocc_iptw_req_bits_store( io_rocc_iptw_req_bits_store ),
       .io_rocc_iptw_req_bits_fetch( io_rocc_iptw_req_bits_fetch ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits_addr( io_rocc_dptw_req_bits_addr ),
       .io_rocc_dptw_req_bits_prv( io_rocc_dptw_req_bits_prv ),
       .io_rocc_dptw_req_bits_store( io_rocc_dptw_req_bits_store ),
       .io_rocc_dptw_req_bits_fetch( io_rocc_dptw_req_bits_fetch ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits_addr( io_rocc_pptw_req_bits_addr ),
       .io_rocc_pptw_req_bits_prv( io_rocc_pptw_req_bits_prv ),
       .io_rocc_pptw_req_bits_store( io_rocc_pptw_req_bits_store ),
       .io_rocc_pptw_req_bits_fetch( io_rocc_pptw_req_bits_fetch ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_exception(  )
       .io_interrupt( csr_io_interrupt ),
       .io_interrupt_cause( csr_io_interrupt_cause )
  );
  ALU alu(
       .io_dw( ex_ctrl_alu_dw ),
       .io_fn( ex_ctrl_alu_fn ),
       .io_in2( T707 ),
       .io_in1( T691 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( T690 ),
       .io_req_bits_fn( ex_ctrl_alu_fn ),
       .io_req_bits_dw( ex_ctrl_alu_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( ex_waddr ),
       .io_kill( T637 ),
       .io_resp_ready( T634 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );

  always @(posedge clk) begin
    if(T517) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T516) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data_0;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T39;
    end
    if(reset) begin
      R73 <= 32'h0;
    end else if(T379) begin
      R73 <= T76;
    end else if(ll_wen) begin
      R73 <= T62;
    end
    if(T517) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if(T516) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if(T103) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if(T517) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if(T516) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if(T103) begin
      ex_ctrl_rocc <= id_ctrl_rocc;
    end
    wb_reg_replay <= T114;
    wb_reg_xcpt <= T118;
    if(T516) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    mem_reg_valid <= T124;
    ex_reg_valid <= T126;
    if(T103) begin
      ex_reg_load_use <= id_load_use;
    end
    if(T517) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if(T516) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if(T103) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if(T516) begin
      bypass_mux_1 <= alu_io_out;
    end
    if(T516) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if(T103) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if(T516) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T516) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if(T103) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if(T516) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if(T103) begin
      ex_reg_flush_pipe <= T243;
    end
    mem_reg_xcpt <= T272;
    if(T103) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    ex_reg_xcpt <= T276;
    ex_reg_xcpt_interrupt <= T359;
    mem_reg_xcpt_interrupt <= T363;
    if(T516) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    mem_reg_replay <= T368;
    wb_reg_valid <= T371;
    if(T517) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if(T516) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if(T517) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if(T516) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if(T103) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if(T516) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T103) begin
      ex_ctrl_mem_type <= id_ctrl_mem_type;
    end
    if(T103) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if(T516) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if(T103) begin
      ex_ctrl_csr <= id_csr;
    end else if(T103) begin
      ex_ctrl_csr <= id_ctrl_csr;
    end
    R521 <= R522;
    if(ex_reg_rs_bypass_1) begin
      R522 <= T573;
    end else begin
      R522 <= T523;
    end
    if(T562) begin
      ex_reg_rs_lsb_1 <= T538;
    end else if(T103) begin
      ex_reg_rs_lsb_1 <= T526;
    end
    if (T543)
      T541[T548] <= rf_wdata;
    if(T517) begin
      bypass_mux_2 <= T553;
    end
    if(T517) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if(T562) begin
      ex_reg_rs_msb_1 <= T572;
    end
    if(T103) begin
      ex_reg_rs_bypass_1 <= T565;
    end
    R584 <= R585;
    if(ex_reg_rs_bypass_0) begin
      R585 <= T613;
    end else begin
      R585 <= T586;
    end
    if(T603) begin
      ex_reg_rs_lsb_0 <= T597;
    end else if(T103) begin
      ex_reg_rs_lsb_0 <= T589;
    end
    if(T603) begin
      ex_reg_rs_msb_0 <= T612;
    end
    if(T103) begin
      ex_reg_rs_bypass_0 <= T606;
    end
    if(T517) begin
      wb_reg_pc <= mem_reg_pc;
    end
    R638 <= T639;
    if(T103) begin
      ex_ctrl_alu_dw <= id_ctrl_alu_dw;
    end
    if(T103) begin
      ex_ctrl_alu_fn <= id_ctrl_alu_fn;
    end
    if(T103) begin
      ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
    end
    if(T103) begin
      ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
    end
    if(T103) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(T826) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(T822) begin
      mem_reg_rs2 <= ex_rs_1;
    end
    if(T103) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if(T517) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if(T516) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if(T103) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if(T886) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T885) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(T103) begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T886) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T885) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T886) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T885) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T886) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T885) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T886) begin
      mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
    end
    if(T885) begin
      ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
    end
    if(T886) begin
      mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
    end
    if(T885) begin
      ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
    end
    if(T886) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T885) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T516) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T632, T630, T629, T627, T625, T624, T623, T621, T583, T581, T520, T519, T1);
// synthesis translate_on
`endif
  end
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [39:0] io_requestor_1_req_bits_addr,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_kill,
    input  io_requestor_1_req_bits_phys,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[39:0] io_requestor_1_resp_bits_addr,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[4:0] io_requestor_1_resp_bits_cmd,
    output[2:0] io_requestor_1_resp_bits_typ,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    input  io_requestor_1_invalidate_lr,
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [39:0] io_requestor_0_req_bits_addr,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_kill,
    input  io_requestor_0_req_bits_phys,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[39:0] io_requestor_0_resp_bits_addr,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[4:0] io_requestor_0_resp_bits_cmd,
    output[2:0] io_requestor_0_resp_bits_typ,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_invalidate_lr
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [7:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered
);

  wire[63:0] T0;
  reg  r_valid_0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[4:0] T4;
  wire[7:0] T32;
  wire[8:0] T5;
  wire[8:0] T6;
  wire[8:0] T7;
  wire[39:0] T8;
  wire T9;
  wire[7:0] T33;
  wire[6:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T34;
  wire[6:0] T18;
  wire T19;
  wire[7:0] T35;
  wire[6:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[7:0] T36;
  wire[6:0] T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_phys = T1;
  assign T1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_kill = T2;
  assign T2 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_bits_typ = T3;
  assign T3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_cmd = T4;
  assign T4 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T5[3'h7:1'h0];
  assign T5 = io_requestor_0_req_valid ? T7 : T6;
  assign T6 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T7 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_addr = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_replay = T14;
  assign T14 = io_mem_resp_bits_replay & T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T17;
  assign T17 = io_mem_resp_bits_nack & T15;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T18};
  assign T18 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T15;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_replay = T24;
  assign T24 = io_mem_resp_bits_replay & T25;
  assign T25 = T26 == 1'h1;
  assign T26 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T27;
  assign T27 = io_mem_resp_bits_nack & T25;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T28};
  assign T28 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T25;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RocketTile(input clk, input reset,
    input  io_cached_acquire_ready,
    output io_cached_acquire_valid,
    output[25:0] io_cached_acquire_bits_addr_block,
    output io_cached_acquire_bits_client_xact_id,
    output[1:0] io_cached_acquire_bits_addr_beat,
    output[127:0] io_cached_acquire_bits_data,
    output io_cached_acquire_bits_is_builtin_type,
    output[2:0] io_cached_acquire_bits_a_type,
    output[16:0] io_cached_acquire_bits_union,
    output io_cached_grant_ready,
    input  io_cached_grant_valid,
    input [1:0] io_cached_grant_bits_addr_beat,
    input [127:0] io_cached_grant_bits_data,
    input  io_cached_grant_bits_client_xact_id,
    input [2:0] io_cached_grant_bits_manager_xact_id,
    input  io_cached_grant_bits_is_builtin_type,
    input [3:0] io_cached_grant_bits_g_type,
    output io_cached_probe_ready,
    input  io_cached_probe_valid,
    input [25:0] io_cached_probe_bits_addr_block,
    input [1:0] io_cached_probe_bits_p_type,
    input  io_cached_release_ready,
    output io_cached_release_valid,
    output[25:0] io_cached_release_bits_addr_block,
    output io_cached_release_bits_client_xact_id,
    output[1:0] io_cached_release_bits_addr_beat,
    output[127:0] io_cached_release_bits_data,
    output[2:0] io_cached_release_bits_r_type,
    output io_cached_release_bits_voluntary,
    input  io_uncached_acquire_ready,
    output io_uncached_acquire_valid,
    output[25:0] io_uncached_acquire_bits_addr_block,
    output io_uncached_acquire_bits_client_xact_id,
    output[1:0] io_uncached_acquire_bits_addr_beat,
    output[127:0] io_uncached_acquire_bits_data,
    output io_uncached_acquire_bits_is_builtin_type,
    output[2:0] io_uncached_acquire_bits_a_type,
    output[16:0] io_uncached_acquire_bits_union,
    output io_uncached_grant_ready,
    input  io_uncached_grant_valid,
    input [1:0] io_uncached_grant_bits_addr_beat,
    input [127:0] io_uncached_grant_bits_data,
    input  io_uncached_grant_bits_client_xact_id,
    input [2:0] io_uncached_grant_bits_manager_xact_id,
    input  io_uncached_grant_bits_is_builtin_type,
    input [3:0] io_uncached_grant_bits_g_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [11:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr
);

  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[7:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[7:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[7:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[7:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire[39:0] dcArb_io_mem_req_bits_addr;
  wire[7:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_kill;
  wire dcArb_io_mem_req_bits_phys;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[19:0] ptw_io_requestor_1_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_1_resp_bits_pte_d;
  wire ptw_io_requestor_1_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_1_resp_bits_pte_typ;
  wire ptw_io_requestor_1_resp_bits_pte_v;
  wire ptw_io_requestor_1_status_sd;
  wire[30:0] ptw_io_requestor_1_status_zero2;
  wire ptw_io_requestor_1_status_sd_rv32;
  wire[8:0] ptw_io_requestor_1_status_zero1;
  wire[4:0] ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_mprv;
  wire[1:0] ptw_io_requestor_1_status_xs;
  wire[1:0] ptw_io_requestor_1_status_fs;
  wire[1:0] ptw_io_requestor_1_status_prv3;
  wire ptw_io_requestor_1_status_ie3;
  wire[1:0] ptw_io_requestor_1_status_prv2;
  wire ptw_io_requestor_1_status_ie2;
  wire[1:0] ptw_io_requestor_1_status_prv1;
  wire ptw_io_requestor_1_status_ie1;
  wire[1:0] ptw_io_requestor_1_status_prv;
  wire ptw_io_requestor_1_status_ie;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[19:0] ptw_io_requestor_0_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_0_resp_bits_pte_d;
  wire ptw_io_requestor_0_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_0_resp_bits_pte_typ;
  wire ptw_io_requestor_0_resp_bits_pte_v;
  wire ptw_io_requestor_0_status_sd;
  wire[30:0] ptw_io_requestor_0_status_zero2;
  wire ptw_io_requestor_0_status_sd_rv32;
  wire[8:0] ptw_io_requestor_0_status_zero1;
  wire[4:0] ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_mprv;
  wire[1:0] ptw_io_requestor_0_status_xs;
  wire[1:0] ptw_io_requestor_0_status_fs;
  wire[1:0] ptw_io_requestor_0_status_prv3;
  wire ptw_io_requestor_0_status_ie3;
  wire[1:0] ptw_io_requestor_0_status_prv2;
  wire ptw_io_requestor_0_status_ie2;
  wire[1:0] ptw_io_requestor_0_status_prv1;
  wire ptw_io_requestor_0_status_ie1;
  wire[1:0] ptw_io_requestor_0_status_prv;
  wire ptw_io_requestor_0_status_ie;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_mem_req_valid;
  wire[39:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_bits_phys;
  wire[63:0] ptw_io_mem_req_bits_data;
  wire core_io_host_pcr_req_ready;
  wire core_io_host_pcr_rep_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_ipi_req_valid;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_debug_stats_pcr;
  wire core_io_imem_req_valid;
  wire[39:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_bits_mask;
  wire core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_btb_update_bits_pc;
  wire[38:0] core_io_imem_btb_update_bits_target;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isReturn;
  wire[38:0] core_io_imem_btb_update_bits_br_pc;
  wire core_io_imem_bht_update_valid;
  wire core_io_imem_bht_update_bits_prediction_valid;
  wire core_io_imem_bht_update_bits_prediction_bits_taken;
  wire core_io_imem_bht_update_bits_prediction_bits_mask;
  wire core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_bht_update_bits_pc;
  wire core_io_imem_bht_update_bits_taken;
  wire core_io_imem_bht_update_bits_mispredict;
  wire core_io_imem_ras_update_valid;
  wire core_io_imem_ras_update_bits_isCall;
  wire core_io_imem_ras_update_bits_isReturn;
  wire[38:0] core_io_imem_ras_update_bits_returnAddr;
  wire core_io_imem_ras_update_bits_prediction_valid;
  wire core_io_imem_ras_update_bits_prediction_bits_taken;
  wire core_io_imem_ras_update_bits_prediction_bits_mask;
  wire core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire[39:0] core_io_dmem_req_bits_addr;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_bits_phys;
  wire[63:0] core_io_dmem_req_bits_data;
  wire core_io_dmem_invalidate_lr;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_status_sd;
  wire[30:0] core_io_ptw_status_zero2;
  wire core_io_ptw_status_sd_rv32;
  wire[8:0] core_io_ptw_status_zero1;
  wire[4:0] core_io_ptw_status_vm;
  wire core_io_ptw_status_mprv;
  wire[1:0] core_io_ptw_status_xs;
  wire[1:0] core_io_ptw_status_fs;
  wire[1:0] core_io_ptw_status_prv3;
  wire core_io_ptw_status_ie3;
  wire[1:0] core_io_ptw_status_prv2;
  wire core_io_ptw_status_ie2;
  wire[1:0] core_io_ptw_status_prv1;
  wire core_io_ptw_status_ie1;
  wire[1:0] core_io_ptw_status_prv;
  wire core_io_ptw_status_ie;
  wire icache_io_cpu_resp_valid;
  wire[39:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data_0;
  wire icache_io_cpu_resp_bits_mask;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_bits_mask;
  wire icache_io_cpu_btb_resp_bits_bridx;
  wire[38:0] icache_io_cpu_btb_resp_bits_target;
  wire[2:0] icache_io_cpu_btb_resp_bits_entry;
  wire[3:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[39:0] icache_io_cpu_npc;
  wire icache_io_ptw_req_valid;
  wire[26:0] icache_io_ptw_req_bits_addr;
  wire[1:0] icache_io_ptw_req_bits_prv;
  wire icache_io_ptw_req_bits_store;
  wire icache_io_ptw_req_bits_fetch;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire icache_io_mem_grant_ready;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[39:0] dcache_io_cpu_resp_bits_addr;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[4:0] dcache_io_cpu_resp_bits_cmd;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ordered;
  wire dcache_io_ptw_req_valid;
  wire[26:0] dcache_io_ptw_req_bits_addr;
  wire[1:0] dcache_io_ptw_req_bits_prv;
  wire dcache_io_ptw_req_bits_store;
  wire dcache_io_ptw_req_bits_fetch;
  wire dcache_io_mem_acquire_valid;
  wire[25:0] dcache_io_mem_acquire_bits_addr_block;
  wire dcache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] dcache_io_mem_acquire_bits_addr_beat;
  wire[127:0] dcache_io_mem_acquire_bits_data;
  wire dcache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] dcache_io_mem_acquire_bits_a_type;
  wire[16:0] dcache_io_mem_acquire_bits_union;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[25:0] dcache_io_mem_release_bits_addr_block;
  wire dcache_io_mem_release_bits_client_xact_id;
  wire[1:0] dcache_io_mem_release_bits_addr_beat;
  wire[127:0] dcache_io_mem_release_bits_data;
  wire[2:0] dcache_io_mem_release_bits_r_type;
  wire dcache_io_mem_release_bits_voluntary;


  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_uncached_grant_ready = icache_io_mem_grant_ready;
  assign io_uncached_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_uncached_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_uncached_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_uncached_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_uncached_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_uncached_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_uncached_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_uncached_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cached_release_bits_voluntary = dcache_io_mem_release_bits_voluntary;
  assign io_cached_release_bits_r_type = dcache_io_mem_release_bits_r_type;
  assign io_cached_release_bits_data = dcache_io_mem_release_bits_data;
  assign io_cached_release_bits_addr_beat = dcache_io_mem_release_bits_addr_beat;
  assign io_cached_release_bits_client_xact_id = dcache_io_mem_release_bits_client_xact_id;
  assign io_cached_release_bits_addr_block = dcache_io_mem_release_bits_addr_block;
  assign io_cached_release_valid = dcache_io_mem_release_valid;
  assign io_cached_probe_ready = dcache_io_mem_probe_ready;
  assign io_cached_grant_ready = dcache_io_mem_grant_ready;
  assign io_cached_acquire_bits_union = dcache_io_mem_acquire_bits_union;
  assign io_cached_acquire_bits_a_type = dcache_io_mem_acquire_bits_a_type;
  assign io_cached_acquire_bits_is_builtin_type = dcache_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_acquire_bits_data = dcache_io_mem_acquire_bits_data;
  assign io_cached_acquire_bits_addr_beat = dcache_io_mem_acquire_bits_addr_beat;
  assign io_cached_acquire_bits_client_xact_id = dcache_io_mem_acquire_bits_client_xact_id;
  assign io_cached_acquire_bits_addr_block = dcache_io_mem_acquire_bits_addr_block;
  assign io_cached_acquire_valid = dcache_io_mem_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_cpu_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_cpu_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_cpu_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_cpu_btb_update_bits_taken(  )
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_cpu_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_cpu_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_cpu_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_cpu_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_cpu_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_cpu_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_cpu_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_cpu_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_cpu_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_cpu_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_cpu_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_cpu_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_cpu_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_cpu_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_cpu_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_cpu_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_cpu_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_cpu_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_cpu_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_cpu_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_cpu_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_cpu_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_cpu_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_cpu_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_cpu_npc( icache_io_cpu_npc ),
       .io_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_ptw_req_valid( icache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_0_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_0_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_0_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_0_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_0_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_acquire_ready( io_uncached_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_uncached_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_uncached_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( io_uncached_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( io_uncached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_uncached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_uncached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_uncached_grant_bits_g_type )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign icache.io_cpu_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_ptw_req_valid( dcache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_1_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_1_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_1_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_1_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_1_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_mem_acquire_ready( io_cached_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( dcache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( dcache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( dcache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_data( dcache_io_mem_acquire_bits_data ),
       .io_mem_acquire_bits_is_builtin_type( dcache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( dcache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( dcache_io_mem_acquire_bits_union ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_cached_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_cached_grant_bits_addr_beat ),
       .io_mem_grant_bits_data( io_cached_grant_bits_data ),
       .io_mem_grant_bits_client_xact_id( io_cached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_cached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_cached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_cached_grant_bits_g_type ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_cached_probe_valid ),
       .io_mem_probe_bits_addr_block( io_cached_probe_bits_addr_block ),
       .io_mem_probe_bits_p_type( io_cached_probe_bits_p_type ),
       .io_mem_release_ready( io_cached_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_addr_block( dcache_io_mem_release_bits_addr_block ),
       .io_mem_release_bits_client_xact_id( dcache_io_mem_release_bits_client_xact_id ),
       .io_mem_release_bits_addr_beat( dcache_io_mem_release_bits_addr_beat ),
       .io_mem_release_bits_data( dcache_io_mem_release_bits_data ),
       .io_mem_release_bits_r_type( dcache_io_mem_release_bits_r_type ),
       .io_mem_release_bits_voluntary( dcache_io_mem_release_bits_voluntary )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_ptw_req_valid ),
       .io_requestor_1_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_requestor_1_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_requestor_1_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_requestor_1_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_requestor_1_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_requestor_1_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_requestor_1_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_requestor_1_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_requestor_1_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_requestor_1_status_sd( ptw_io_requestor_1_status_sd ),
       .io_requestor_1_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_requestor_1_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_requestor_1_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_requestor_1_status_xs( ptw_io_requestor_1_status_xs ),
       .io_requestor_1_status_fs( ptw_io_requestor_1_status_fs ),
       .io_requestor_1_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_requestor_1_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_requestor_1_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_requestor_1_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_requestor_1_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_requestor_1_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_requestor_1_status_prv( ptw_io_requestor_1_status_prv ),
       .io_requestor_1_status_ie( ptw_io_requestor_1_status_ie ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_ptw_req_valid ),
       .io_requestor_0_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_requestor_0_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_requestor_0_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_requestor_0_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_requestor_0_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_requestor_0_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_requestor_0_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_requestor_0_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_requestor_0_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_requestor_0_status_sd( ptw_io_requestor_0_status_sd ),
       .io_requestor_0_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_requestor_0_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_requestor_0_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_requestor_0_status_xs( ptw_io_requestor_0_status_xs ),
       .io_requestor_0_status_fs( ptw_io_requestor_0_status_fs ),
       .io_requestor_0_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_requestor_0_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_requestor_0_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_requestor_0_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_requestor_0_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_requestor_0_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_requestor_0_status_prv( ptw_io_requestor_0_status_prv ),
       .io_requestor_0_status_ie( ptw_io_requestor_0_status_ie ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_status_sd( core_io_ptw_status_sd ),
       .io_dpath_status_zero2( core_io_ptw_status_zero2 ),
       .io_dpath_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_dpath_status_zero1( core_io_ptw_status_zero1 ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_mprv( core_io_ptw_status_mprv ),
       .io_dpath_status_xs( core_io_ptw_status_xs ),
       .io_dpath_status_fs( core_io_ptw_status_fs ),
       .io_dpath_status_prv3( core_io_ptw_status_prv3 ),
       .io_dpath_status_ie3( core_io_ptw_status_ie3 ),
       .io_dpath_status_prv2( core_io_ptw_status_prv2 ),
       .io_dpath_status_ie2( core_io_ptw_status_ie2 ),
       .io_dpath_status_prv1( core_io_ptw_status_prv1 ),
       .io_dpath_status_ie1( core_io_ptw_status_ie1 ),
       .io_dpath_status_prv( core_io_ptw_status_prv ),
       .io_dpath_status_ie( core_io_ptw_status_ie )
  );
  Rocket core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_imem_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_imem_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_imem_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_imem_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_imem_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_imem_npc( icache_io_cpu_npc ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_dmem_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_status_sd( core_io_ptw_status_sd ),
       .io_ptw_status_zero2( core_io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( core_io_ptw_status_zero1 ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_mprv( core_io_ptw_status_mprv ),
       .io_ptw_status_xs( core_io_ptw_status_xs ),
       .io_ptw_status_fs( core_io_ptw_status_fs ),
       .io_ptw_status_prv3( core_io_ptw_status_prv3 ),
       .io_ptw_status_ie3( core_io_ptw_status_ie3 ),
       .io_ptw_status_prv2( core_io_ptw_status_prv2 ),
       .io_ptw_status_ie2( core_io_ptw_status_ie2 ),
       .io_ptw_status_prv1( core_io_ptw_status_prv1 ),
       .io_ptw_status_ie1( core_io_ptw_status_ie1 ),
       .io_ptw_status_prv( core_io_ptw_status_prv ),
       .io_ptw_status_ie( core_io_ptw_status_ie )
       //.io_fpu_inst(  )
       //.io_fpu_fromint_data(  )
       //.io_fpu_fcsr_rm(  )
       //.io_fpu_fcsr_flags_valid(  )
       //.io_fpu_fcsr_flags_bits(  )
       //.io_fpu_store_data(  )
       //.io_fpu_toint_data(  )
       //.io_fpu_dmem_resp_val(  )
       //.io_fpu_dmem_resp_type(  )
       //.io_fpu_dmem_resp_tag(  )
       //.io_fpu_dmem_resp_data(  )
       //.io_fpu_valid(  )
       //.io_fpu_fcsr_rdy(  )
       //.io_fpu_nack_mem(  )
       //.io_fpu_illegal_rm(  )
       //.io_fpu_killx(  )
       //.io_fpu_killm(  )
       //.io_fpu_dec_cmd(  )
       //.io_fpu_dec_ldst(  )
       //.io_fpu_dec_wen(  )
       //.io_fpu_dec_ren1(  )
       //.io_fpu_dec_ren2(  )
       //.io_fpu_dec_ren3(  )
       //.io_fpu_dec_swap12(  )
       //.io_fpu_dec_swap23(  )
       //.io_fpu_dec_single(  )
       //.io_fpu_dec_fromint(  )
       //.io_fpu_dec_toint(  )
       //.io_fpu_dec_fastpipe(  )
       //.io_fpu_dec_fma(  )
       //.io_fpu_dec_div(  )
       //.io_fpu_dec_sqrt(  )
       //.io_fpu_dec_round(  )
       //.io_fpu_dec_wflags(  )
       //.io_fpu_sboard_set(  )
       //.io_fpu_sboard_clr(  )
       //.io_fpu_sboard_clra(  )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_invalidate_lr(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_addr_block(  )
       //.io_rocc_imem_acquire_bits_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_addr_beat(  )
       //.io_rocc_imem_acquire_bits_data(  )
       //.io_rocc_imem_acquire_bits_is_builtin_type(  )
       //.io_rocc_imem_acquire_bits_a_type(  )
       //.io_rocc_imem_acquire_bits_union(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_addr_beat(  )
       //.io_rocc_imem_grant_bits_data(  )
       //.io_rocc_imem_grant_bits_client_xact_id(  )
       //.io_rocc_imem_grant_bits_manager_xact_id(  )
       //.io_rocc_imem_grant_bits_is_builtin_type(  )
       //.io_rocc_imem_grant_bits_g_type(  )
       //.io_rocc_dmem_acquire_ready(  )
       //.io_rocc_dmem_acquire_valid(  )
       //.io_rocc_dmem_acquire_bits_addr_block(  )
       //.io_rocc_dmem_acquire_bits_client_xact_id(  )
       //.io_rocc_dmem_acquire_bits_addr_beat(  )
       //.io_rocc_dmem_acquire_bits_data(  )
       //.io_rocc_dmem_acquire_bits_is_builtin_type(  )
       //.io_rocc_dmem_acquire_bits_a_type(  )
       //.io_rocc_dmem_acquire_bits_union(  )
       //.io_rocc_dmem_grant_ready(  )
       //.io_rocc_dmem_grant_valid(  )
       //.io_rocc_dmem_grant_bits_addr_beat(  )
       //.io_rocc_dmem_grant_bits_data(  )
       //.io_rocc_dmem_grant_bits_client_xact_id(  )
       //.io_rocc_dmem_grant_bits_manager_xact_id(  )
       //.io_rocc_dmem_grant_bits_is_builtin_type(  )
       //.io_rocc_dmem_grant_bits_g_type(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits_addr(  )
       //.io_rocc_iptw_req_bits_prv(  )
       //.io_rocc_iptw_req_bits_store(  )
       //.io_rocc_iptw_req_bits_fetch(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits_addr(  )
       //.io_rocc_dptw_req_bits_prv(  )
       //.io_rocc_dptw_req_bits_store(  )
       //.io_rocc_dptw_req_bits_fetch(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits_addr(  )
       //.io_rocc_pptw_req_bits_prv(  )
       //.io_rocc_pptw_req_bits_store(  )
       //.io_rocc_pptw_req_bits_fetch(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_exception(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign core.io_fpu_fcsr_flags_valid = {1{$random}};
    assign core.io_fpu_fcsr_flags_bits = {1{$random}};
    assign core.io_fpu_store_data = {2{$random}};
    assign core.io_fpu_toint_data = {2{$random}};
    assign core.io_fpu_nack_mem = {1{$random}};
    assign core.io_fpu_illegal_rm = {1{$random}};
    assign core.io_fpu_dec_wen = {1{$random}};
    assign core.io_fpu_dec_ren1 = {1{$random}};
    assign core.io_fpu_dec_ren2 = {1{$random}};
    assign core.io_fpu_dec_ren3 = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_invalidate_lr = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_data = {4{$random}};
    assign core.io_rocc_imem_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_union = {1{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_dmem_acquire_valid = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_data = {4{$random}};
    assign core.io_rocc_dmem_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_dmem_acquire_bits_union = {1{$random}};
    assign core.io_rocc_dmem_grant_ready = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_iptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_iptw_req_bits_store = {1{$random}};
    assign core.io_rocc_iptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_dptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_dptw_req_bits_store = {1{$random}};
    assign core.io_rocc_dptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_pptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_pptw_req_bits_store = {1{$random}};
    assign core.io_rocc_pptw_req_bits_fetch = {1{$random}};
// synthesis translate_on
`endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_requestor_1_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_invalidate_lr(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [11:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[11:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[76:0] T11;
  reg [76:0] ram [1:0];
  wire[76:0] T12;
  wire[76:0] T13;
  wire[76:0] T14;
  wire[75:0] T15;
  wire[11:0] T16;
  wire T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rw, T15};
  assign T15 = {io_enq_bits_addr, io_enq_bits_data};
  assign io_deq_bits_addr = T16;
  assign T16 = T11[7'h4b:7'h40];
  assign io_deq_bits_rw = T17;
  assign T17 = T11[7'h4c:7'h4c];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[63:0] T10;
  reg [63:0] ram [1:0];
  wire[63:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire T10;
  reg [0:0] ram [1:0];
  wire T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module MultiChannelTop(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    //output io_mem_backup_ctrl_out_valid
    input  io_mem_0_req_cmd_ready,
    output io_mem_0_req_cmd_valid,
    output[25:0] io_mem_0_req_cmd_bits_addr,
    output[5:0] io_mem_0_req_cmd_bits_tag,
    output io_mem_0_req_cmd_bits_rw,
    input  io_mem_0_req_data_ready,
    output io_mem_0_req_data_valid,
    output[127:0] io_mem_0_req_data_bits_data,
    output io_mem_0_resp_ready,
    input  io_mem_0_resp_valid,
    input [127:0] io_mem_0_resp_bits_data,
    input [5:0] io_mem_0_resp_bits_tag
);

  reg  R0;
  reg  R1;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire Queue_io_deq_bits_rw;
  wire[11:0] Queue_io_deq_bits_addr;
  wire[63:0] Queue_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire Queue_2_io_deq_bits;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire Queue_3_io_deq_bits;
  wire RocketTile_io_cached_acquire_valid;
  wire[25:0] RocketTile_io_cached_acquire_bits_addr_block;
  wire RocketTile_io_cached_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_cached_acquire_bits_addr_beat;
  wire[127:0] RocketTile_io_cached_acquire_bits_data;
  wire RocketTile_io_cached_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_cached_acquire_bits_a_type;
  wire[16:0] RocketTile_io_cached_acquire_bits_union;
  wire RocketTile_io_cached_grant_ready;
  wire RocketTile_io_cached_probe_ready;
  wire RocketTile_io_cached_release_valid;
  wire[25:0] RocketTile_io_cached_release_bits_addr_block;
  wire RocketTile_io_cached_release_bits_client_xact_id;
  wire[1:0] RocketTile_io_cached_release_bits_addr_beat;
  wire[127:0] RocketTile_io_cached_release_bits_data;
  wire[2:0] RocketTile_io_cached_release_bits_r_type;
  wire RocketTile_io_cached_release_bits_voluntary;
  wire RocketTile_io_uncached_acquire_valid;
  wire[25:0] RocketTile_io_uncached_acquire_bits_addr_block;
  wire RocketTile_io_uncached_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_uncached_acquire_bits_addr_beat;
  wire[127:0] RocketTile_io_uncached_acquire_bits_data;
  wire RocketTile_io_uncached_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_uncached_acquire_bits_a_type;
  wire[16:0] RocketTile_io_uncached_acquire_bits_union;
  wire RocketTile_io_uncached_grant_ready;
  wire RocketTile_io_host_pcr_req_ready;
  wire RocketTile_io_host_pcr_rep_valid;
  wire[63:0] RocketTile_io_host_pcr_rep_bits;
  wire RocketTile_io_host_ipi_req_valid;
  wire RocketTile_io_host_ipi_req_bits;
  wire RocketTile_io_host_ipi_rep_ready;
  wire RocketTile_io_host_debug_stats_pcr;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_pcr;
  wire uncore_io_mem_0_req_cmd_valid;
  wire[25:0] uncore_io_mem_0_req_cmd_bits_addr;
  wire[5:0] uncore_io_mem_0_req_cmd_bits_tag;
  wire uncore_io_mem_0_req_cmd_bits_rw;
  wire uncore_io_mem_0_req_data_valid;
  wire[127:0] uncore_io_mem_0_req_data_bits_data;
  wire uncore_io_mem_0_resp_ready;
  wire uncore_io_tiles_cached_0_acquire_ready;
  wire uncore_io_tiles_cached_0_grant_valid;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire[127:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[2:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire uncore_io_tiles_cached_0_probe_valid;
  wire[25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire uncore_io_tiles_cached_0_release_ready;
  wire uncore_io_tiles_uncached_0_acquire_ready;
  wire uncore_io_tiles_uncached_0_grant_valid;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[127:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[2:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_pcr_req_valid;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire[11:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire uncore_io_htif_0_ipi_req_ready;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_rep_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_0_resp_ready = uncore_io_mem_0_resp_ready;
  assign io_mem_0_req_data_bits_data = uncore_io_mem_0_req_data_bits_data;
  assign io_mem_0_req_data_valid = uncore_io_mem_0_req_data_valid;
  assign io_mem_0_req_cmd_bits_rw = uncore_io_mem_0_req_cmd_bits_rw;
  assign io_mem_0_req_cmd_bits_tag = uncore_io_mem_0_req_cmd_bits_tag;
  assign io_mem_0_req_cmd_bits_addr = uncore_io_mem_0_req_cmd_bits_addr;
  assign io_mem_0_req_cmd_valid = uncore_io_mem_0_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_0_req_cmd_ready( io_mem_0_req_cmd_ready ),
       .io_mem_0_req_cmd_valid( uncore_io_mem_0_req_cmd_valid ),
       .io_mem_0_req_cmd_bits_addr( uncore_io_mem_0_req_cmd_bits_addr ),
       .io_mem_0_req_cmd_bits_tag( uncore_io_mem_0_req_cmd_bits_tag ),
       .io_mem_0_req_cmd_bits_rw( uncore_io_mem_0_req_cmd_bits_rw ),
       .io_mem_0_req_data_ready( io_mem_0_req_data_ready ),
       .io_mem_0_req_data_valid( uncore_io_mem_0_req_data_valid ),
       .io_mem_0_req_data_bits_data( uncore_io_mem_0_req_data_bits_data ),
       .io_mem_0_resp_ready( uncore_io_mem_0_resp_ready ),
       .io_mem_0_resp_valid( io_mem_0_resp_valid ),
       .io_mem_0_resp_bits_data( io_mem_0_resp_bits_data ),
       .io_mem_0_resp_bits_tag( io_mem_0_resp_bits_tag ),
       .io_tiles_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( RocketTile_io_cached_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( RocketTile_io_cached_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_data( RocketTile_io_cached_acquire_bits_data ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( RocketTile_io_cached_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( RocketTile_io_cached_acquire_bits_union ),
       .io_tiles_cached_0_grant_ready( RocketTile_io_cached_grant_ready ),
       .io_tiles_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_probe_ready( RocketTile_io_cached_probe_ready ),
       .io_tiles_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( RocketTile_io_cached_release_valid ),
       .io_tiles_cached_0_release_bits_addr_block( RocketTile_io_cached_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( RocketTile_io_cached_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_addr_beat( RocketTile_io_cached_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_data( RocketTile_io_cached_release_bits_data ),
       .io_tiles_cached_0_release_bits_r_type( RocketTile_io_cached_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_voluntary( RocketTile_io_cached_release_bits_voluntary ),
       .io_tiles_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( RocketTile_io_uncached_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_data( RocketTile_io_uncached_acquire_bits_data ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( RocketTile_io_uncached_acquire_bits_union ),
       .io_tiles_uncached_0_grant_ready( RocketTile_io_uncached_grant_ready ),
       .io_tiles_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr )
       //.io_mem_backup_ctrl_en(  )
       //.io_mem_backup_ctrl_in_valid(  )
       //.io_mem_backup_ctrl_out_ready(  )
       //.io_mem_backup_ctrl_out_valid(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
// synthesis translate_on
`endif
  RocketTile RocketTile(.clk(clk), .reset(uncore_io_htif_0_reset),
       .io_cached_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_cached_acquire_valid( RocketTile_io_cached_acquire_valid ),
       .io_cached_acquire_bits_addr_block( RocketTile_io_cached_acquire_bits_addr_block ),
       .io_cached_acquire_bits_client_xact_id( RocketTile_io_cached_acquire_bits_client_xact_id ),
       .io_cached_acquire_bits_addr_beat( RocketTile_io_cached_acquire_bits_addr_beat ),
       .io_cached_acquire_bits_data( RocketTile_io_cached_acquire_bits_data ),
       .io_cached_acquire_bits_is_builtin_type( RocketTile_io_cached_acquire_bits_is_builtin_type ),
       .io_cached_acquire_bits_a_type( RocketTile_io_cached_acquire_bits_a_type ),
       .io_cached_acquire_bits_union( RocketTile_io_cached_acquire_bits_union ),
       .io_cached_grant_ready( RocketTile_io_cached_grant_ready ),
       .io_cached_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_cached_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_cached_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_cached_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_cached_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_cached_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_cached_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_cached_probe_ready( RocketTile_io_cached_probe_ready ),
       .io_cached_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_cached_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_cached_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_cached_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_cached_release_valid( RocketTile_io_cached_release_valid ),
       .io_cached_release_bits_addr_block( RocketTile_io_cached_release_bits_addr_block ),
       .io_cached_release_bits_client_xact_id( RocketTile_io_cached_release_bits_client_xact_id ),
       .io_cached_release_bits_addr_beat( RocketTile_io_cached_release_bits_addr_beat ),
       .io_cached_release_bits_data( RocketTile_io_cached_release_bits_data ),
       .io_cached_release_bits_r_type( RocketTile_io_cached_release_bits_r_type ),
       .io_cached_release_bits_voluntary( RocketTile_io_cached_release_bits_voluntary ),
       .io_uncached_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_uncached_acquire_valid( RocketTile_io_uncached_acquire_valid ),
       .io_uncached_acquire_bits_addr_block( RocketTile_io_uncached_acquire_bits_addr_block ),
       .io_uncached_acquire_bits_client_xact_id( RocketTile_io_uncached_acquire_bits_client_xact_id ),
       .io_uncached_acquire_bits_addr_beat( RocketTile_io_uncached_acquire_bits_addr_beat ),
       .io_uncached_acquire_bits_data( RocketTile_io_uncached_acquire_bits_data ),
       .io_uncached_acquire_bits_is_builtin_type( RocketTile_io_uncached_acquire_bits_is_builtin_type ),
       .io_uncached_acquire_bits_a_type( RocketTile_io_uncached_acquire_bits_a_type ),
       .io_uncached_acquire_bits_union( RocketTile_io_uncached_acquire_bits_union ),
       .io_uncached_grant_ready( RocketTile_io_uncached_grant_ready ),
       .io_uncached_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_uncached_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_uncached_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_uncached_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_uncached_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_uncached_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_uncached_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( RocketTile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( RocketTile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( RocketTile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( RocketTile_io_host_debug_stats_pcr )
  );
  Queue_0 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_rw( Queue_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_pcr_rep_valid ),
       .io_enq_bits( RocketTile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_ipi_req_valid ),
       .io_enq_bits( RocketTile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( RocketTile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module MemIOArbiter(
    output io_inner_0_req_cmd_ready,
    input  io_inner_0_req_cmd_valid,
    input [25:0] io_inner_0_req_cmd_bits_addr,
    input [5:0] io_inner_0_req_cmd_bits_tag,
    input  io_inner_0_req_cmd_bits_rw,
    output io_inner_0_req_data_ready,
    input  io_inner_0_req_data_valid,
    input [127:0] io_inner_0_req_data_bits_data,
    input  io_inner_0_resp_ready,
    output io_inner_0_resp_valid,
    output[127:0] io_inner_0_resp_bits_data,
    output[5:0] io_inner_0_resp_bits_tag,
    input  io_outer_req_cmd_ready,
    output io_outer_req_cmd_valid,
    output[25:0] io_outer_req_cmd_bits_addr,
    output[5:0] io_outer_req_cmd_bits_tag,
    output io_outer_req_cmd_bits_rw,
    input  io_outer_req_data_ready,
    output io_outer_req_data_valid,
    output[127:0] io_outer_req_data_bits_data,
    output io_outer_resp_ready,
    input  io_outer_resp_valid,
    input [127:0] io_outer_resp_bits_data,
    input [5:0] io_outer_resp_bits_tag
);



  assign io_outer_resp_ready = io_inner_0_resp_ready;
  assign io_outer_req_data_bits_data = io_inner_0_req_data_bits_data;
  assign io_outer_req_data_valid = io_inner_0_req_data_valid;
  assign io_outer_req_cmd_bits_rw = io_inner_0_req_cmd_bits_rw;
  assign io_outer_req_cmd_bits_tag = io_inner_0_req_cmd_bits_tag;
  assign io_outer_req_cmd_bits_addr = io_inner_0_req_cmd_bits_addr;
  assign io_outer_req_cmd_valid = io_inner_0_req_cmd_valid;
  assign io_inner_0_resp_bits_tag = io_outer_resp_bits_tag;
  assign io_inner_0_resp_bits_data = io_outer_resp_bits_data;
  assign io_inner_0_resp_valid = io_outer_resp_valid;
  assign io_inner_0_req_data_ready = io_outer_req_data_ready;
  assign io_inner_0_req_cmd_ready = io_outer_req_cmd_ready;
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    output io_mem_backup_ctrl_out_valid,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[5:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [5:0] io_mem_resp_bits_tag
);

  wire MemIOArbiter_io_inner_0_req_cmd_ready;
  wire MemIOArbiter_io_inner_0_req_data_ready;
  wire MemIOArbiter_io_inner_0_resp_valid;
  wire[127:0] MemIOArbiter_io_inner_0_resp_bits_data;
  wire[5:0] MemIOArbiter_io_inner_0_resp_bits_tag;
  wire MemIOArbiter_io_outer_req_cmd_valid;
  wire[25:0] MemIOArbiter_io_outer_req_cmd_bits_addr;
  wire[5:0] MemIOArbiter_io_outer_req_cmd_bits_tag;
  wire MemIOArbiter_io_outer_req_cmd_bits_rw;
  wire MemIOArbiter_io_outer_req_data_valid;
  wire[127:0] MemIOArbiter_io_outer_req_data_bits_data;
  wire MemIOArbiter_io_outer_resp_ready;
  wire MultiChannelTop_io_host_in_ready;
  wire MultiChannelTop_io_host_out_valid;
  wire[15:0] MultiChannelTop_io_host_out_bits;
  wire MultiChannelTop_io_host_debug_stats_pcr;
  wire MultiChannelTop_io_mem_0_req_cmd_valid;
  wire[25:0] MultiChannelTop_io_mem_0_req_cmd_bits_addr;
  wire[5:0] MultiChannelTop_io_mem_0_req_cmd_bits_tag;
  wire MultiChannelTop_io_mem_0_req_cmd_bits_rw;
  wire MultiChannelTop_io_mem_0_req_data_valid;
  wire[127:0] MultiChannelTop_io_mem_0_req_data_bits_data;
  wire MultiChannelTop_io_mem_0_resp_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_resp_ready = MemIOArbiter_io_outer_resp_ready;
  assign io_mem_req_data_bits_data = MemIOArbiter_io_outer_req_data_bits_data;
  assign io_mem_req_data_valid = MemIOArbiter_io_outer_req_data_valid;
  assign io_mem_req_cmd_bits_rw = MemIOArbiter_io_outer_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = MemIOArbiter_io_outer_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = MemIOArbiter_io_outer_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = MemIOArbiter_io_outer_req_cmd_valid;
  assign io_host_debug_stats_pcr = MultiChannelTop_io_host_debug_stats_pcr;
  assign io_host_out_bits = MultiChannelTop_io_host_out_bits;
  assign io_host_out_valid = MultiChannelTop_io_host_out_valid;
  assign io_host_in_ready = MultiChannelTop_io_host_in_ready;
  MultiChannelTop MultiChannelTop(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( MultiChannelTop_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( MultiChannelTop_io_host_out_valid ),
       .io_host_out_bits( MultiChannelTop_io_host_out_bits ),
       .io_host_debug_stats_pcr( MultiChannelTop_io_host_debug_stats_pcr ),
       .io_mem_backup_ctrl_en( io_mem_backup_ctrl_en ),
       .io_mem_backup_ctrl_in_valid( io_mem_backup_ctrl_in_valid ),
       .io_mem_backup_ctrl_out_ready( io_mem_backup_ctrl_out_ready ),
       //.io_mem_backup_ctrl_out_valid(  )
       .io_mem_0_req_cmd_ready( MemIOArbiter_io_inner_0_req_cmd_ready ),
       .io_mem_0_req_cmd_valid( MultiChannelTop_io_mem_0_req_cmd_valid ),
       .io_mem_0_req_cmd_bits_addr( MultiChannelTop_io_mem_0_req_cmd_bits_addr ),
       .io_mem_0_req_cmd_bits_tag( MultiChannelTop_io_mem_0_req_cmd_bits_tag ),
       .io_mem_0_req_cmd_bits_rw( MultiChannelTop_io_mem_0_req_cmd_bits_rw ),
       .io_mem_0_req_data_ready( MemIOArbiter_io_inner_0_req_data_ready ),
       .io_mem_0_req_data_valid( MultiChannelTop_io_mem_0_req_data_valid ),
       .io_mem_0_req_data_bits_data( MultiChannelTop_io_mem_0_req_data_bits_data ),
       .io_mem_0_resp_ready( MultiChannelTop_io_mem_0_resp_ready ),
       .io_mem_0_resp_valid( MemIOArbiter_io_inner_0_resp_valid ),
       .io_mem_0_resp_bits_data( MemIOArbiter_io_inner_0_resp_bits_data ),
       .io_mem_0_resp_bits_tag( MemIOArbiter_io_inner_0_resp_bits_tag )
  );
  MemIOArbiter MemIOArbiter(
       .io_inner_0_req_cmd_ready( MemIOArbiter_io_inner_0_req_cmd_ready ),
       .io_inner_0_req_cmd_valid( MultiChannelTop_io_mem_0_req_cmd_valid ),
       .io_inner_0_req_cmd_bits_addr( MultiChannelTop_io_mem_0_req_cmd_bits_addr ),
       .io_inner_0_req_cmd_bits_tag( MultiChannelTop_io_mem_0_req_cmd_bits_tag ),
       .io_inner_0_req_cmd_bits_rw( MultiChannelTop_io_mem_0_req_cmd_bits_rw ),
       .io_inner_0_req_data_ready( MemIOArbiter_io_inner_0_req_data_ready ),
       .io_inner_0_req_data_valid( MultiChannelTop_io_mem_0_req_data_valid ),
       .io_inner_0_req_data_bits_data( MultiChannelTop_io_mem_0_req_data_bits_data ),
       .io_inner_0_resp_ready( MultiChannelTop_io_mem_0_resp_ready ),
       .io_inner_0_resp_valid( MemIOArbiter_io_inner_0_resp_valid ),
       .io_inner_0_resp_bits_data( MemIOArbiter_io_inner_0_resp_bits_data ),
       .io_inner_0_resp_bits_tag( MemIOArbiter_io_inner_0_resp_bits_tag ),
       .io_outer_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_outer_req_cmd_valid( MemIOArbiter_io_outer_req_cmd_valid ),
       .io_outer_req_cmd_bits_addr( MemIOArbiter_io_outer_req_cmd_bits_addr ),
       .io_outer_req_cmd_bits_tag( MemIOArbiter_io_outer_req_cmd_bits_tag ),
       .io_outer_req_cmd_bits_rw( MemIOArbiter_io_outer_req_cmd_bits_rw ),
       .io_outer_req_data_ready( io_mem_req_data_ready ),
       .io_outer_req_data_valid( MemIOArbiter_io_outer_req_data_valid ),
       .io_outer_req_data_bits_data( MemIOArbiter_io_outer_req_data_bits_data ),
       .io_outer_resp_ready( MemIOArbiter_io_outer_resp_ready ),
       .io_outer_resp_valid( io_mem_resp_valid ),
       .io_outer_resp_bits_data( io_mem_resp_bits_data ),
       .io_outer_resp_bits_tag( io_mem_resp_bits_tag )
  );
endmodule

module DataArray_T1(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_T1(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [21:0] W0I,
  input [21:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [21:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+22) begin
    for (j=1; j<22; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [21:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][21:0] <= W0I[21:0];
end
assign R1O = ram[reg_R1A];

endmodule


module HellaFlowQueue_T3_1(
  input CLK,
  input RST,
  input init,
  input [4:0] W0A,
  input W0E,
  input [5:0] W0I,
  input [4:0] R1A,
  input R1E,
  output [5:0] R1O
);

reg [5:0] ram [23:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 24; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [4:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_T86(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [19:0] RW0M,
  input [19:0] RW0I,
  output [19:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+20) begin
    for (j=1; j<20; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [19:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][19:0] <= RW0I[19:0];
end
assign RW0O = ram[reg_RW0A];

endmodule


module ICache_T109(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


module HellaFlowQueue_T3(
  input CLK,
  input RST,
  input init,
  input [4:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [4:0] R1A,
  input R1E,
  output [127:0] R1O
);

reg [127:0] ram [23:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 24; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [4:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E) ram[W0A] <= W0I;
end
assign R1O = ram[reg_R1A];

endmodule


