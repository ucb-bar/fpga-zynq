module Htif(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    output io_cpu_0_reset,
    output io_cpu_0_id,
    input  io_cpu_0_csr_req_ready,
    output io_cpu_0_csr_req_valid,
    output io_cpu_0_csr_req_bits_rw,
    output[11:0] io_cpu_0_csr_req_bits_addr,
    output[63:0] io_cpu_0_csr_req_bits_data,
    output io_cpu_0_csr_resp_ready,
    input  io_cpu_0_csr_resp_valid,
    input [63:0] io_cpu_0_csr_resp_bits,
    input  io_cpu_0_debug_stats_csr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits
);

  wire[63:0] csr_wdata;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire T3;
  reg [2:0] state;
  wire[2:0] T210;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[3:0] rx_cmd;
  reg [3:0] cmd;
  wire[3:0] T20;
  wire T21;
  wire T22;
  reg [14:0] rx_count;
  wire[14:0] T211;
  wire[14:0] T23;
  wire[14:0] T24;
  wire[14:0] T25;
  wire T26;
  wire T27;
  wire[12:0] T212;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T28;
  wire[11:0] T29;
  wire[63:0] rx_shifter_in;
  wire[47:0] T30;
  reg [63:0] rx_shifter;
  wire[63:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire nack;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire bad_mem_packet;
  wire T44;
  wire[2:0] T45;
  reg [39:0] addr;
  wire[39:0] T46;
  wire[39:0] T47;
  wire[39:0] T48;
  wire[39:0] T49;
  wire[39:0] T50;
  wire[39:0] T51;
  wire T52;
  wire[2:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[12:0] tx_word_count;
  reg [14:0] tx_count;
  wire[14:0] T213;
  wire[14:0] T57;
  wire[14:0] T58;
  wire[14:0] T59;
  wire T60;
  wire T61;
  wire[3:0] next_cmd;
  wire T62;
  wire[12:0] rx_word_count;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire rx_done;
  wire T67;
  wire T68;
  wire T69;
  wire[2:0] T70;
  wire T71;
  wire[12:0] T214;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire rx_word_done;
  wire T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire cnt_done;
  wire T80;
  reg [1:0] cnt;
  wire[1:0] T215;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  reg [8:0] pos;
  wire[8:0] T94;
  wire[8:0] T95;
  wire[8:0] T96;
  wire[8:0] T97;
  wire[8:0] T98;
  wire[8:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[2:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[2:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire tx_done;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T117;
  wire T118;
  wire T119;
  wire[12:0] T216;
  wire T120;
  wire T121;
  wire[1:0] tx_subword_count;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire[11:0] csr_addr;
  wire T126;
  wire T127;
  wire[1:0] csr_coreid;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[2:0] T134;
  wire[63:0] T135;
  wire[63:0] T136;
  wire T137;
  wire T138;
  wire[2:0] T139;
  wire[63:0] T140;
  wire T141;
  wire[2:0] T142;
  wire[2:0] T143;
  wire[5:0] T144;
  wire[5:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[127:0] T150;
  wire[127:0] T151;
  wire[127:0] T152;
  wire[127:0] mem_req_data;
  wire[63:0] T153;
  wire[2:0] T154;
  wire[63:0] T155;
  wire[2:0] T156;
  wire T157;
  wire[16:0] T158;
  wire[16:0] T159;
  wire[16:0] T160;
  wire[16:0] T161;
  wire[15:0] T162;
  wire[2:0] T163;
  wire[2:0] T164;
  wire[2:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] T169;
  wire[1:0] T170;
  wire[1:0] T171;
  wire[1:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[25:0] T175;
  wire[25:0] T176;
  wire[25:0] T217;
  wire[36:0] init_addr;
  wire[39:0] T177;
  wire[25:0] T178;
  wire[25:0] T218;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg  R187;
  wire T219;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire[15:0] T220;
  wire[63:0] T192;
  wire[5:0] T193;
  wire[1:0] T194;
  wire[63:0] tx_data;
  wire[63:0] T195;
  wire[63:0] T196;
  reg [63:0] csrReadData;
  wire[63:0] T197;
  wire[63:0] T198;
  wire[63:0] T199;
  wire[63:0] T221;
  wire T200;
  wire T201;
  wire T202;
  wire[63:0] tx_header;
  wire[15:0] T203;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T204;
  reg [7:0] seqno;
  wire[7:0] T205;
  wire[7:0] T206;
  wire T207;
  wire T208;
  wire T209;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    state = {1{$random}};
    cmd = {1{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    rx_shifter = {2{$random}};
    addr = {2{$random}};
    tx_count = {1{$random}};
    cnt = {1{$random}};
    pos = {1{$random}};
    R187 = {1{$random}};
    csrReadData = {2{$random}};
    seqno = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
  assign io_cpu_0_id = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_scr_resp_ready = 1'h1;
  assign io_scr_req_bits_data = csr_wdata;
  assign csr_wdata = packet_ram[3'h0];
  assign T1 = io_mem_grant_bits_data[7'h7f:7'h40];
  assign T2 = T3 & io_mem_grant_valid;
  assign T3 = state == 3'h5;
  assign T210 = reset ? 3'h0 : T4;
  assign T4 = T132 ? 3'h7 : T5;
  assign T5 = T131 ? 3'h2 : T6;
  assign T6 = T129 ? 3'h7 : T7;
  assign T7 = T124 ? 3'h7 : T8;
  assign T8 = T123 ? 3'h2 : T9;
  assign T9 = T113 ? T109 : T10;
  assign T10 = T107 ? T103 : T11;
  assign T11 = T101 ? T91 : T12;
  assign T12 = T89 ? 3'h5 : T13;
  assign T13 = T79 ? 3'h6 : T14;
  assign T14 = T66 ? T15 : state;
  assign T15 = T65 ? 3'h3 : T16;
  assign T16 = T64 ? 3'h4 : T17;
  assign T17 = T18 ? 3'h1 : 3'h7;
  assign T18 = T63 | T19;
  assign T19 = rx_cmd == 4'h3;
  assign rx_cmd = T62 ? next_cmd : cmd;
  assign T20 = T21 ? next_cmd : cmd;
  assign T21 = T61 & T22;
  assign T22 = rx_count == 15'h3;
  assign T211 = reset ? 15'h0 : T23;
  assign T23 = T26 ? 15'h0 : T24;
  assign T24 = T61 ? T25 : rx_count;
  assign T25 = rx_count + 15'h1;
  assign T26 = T113 & T27;
  assign T27 = tx_word_count == T212;
  assign T212 = {1'h0, tx_size};
  assign tx_size = T32 ? size : 12'h0;
  assign T28 = T21 ? T29 : size;
  assign T29 = rx_shifter_in[4'hf:3'h4];
  assign rx_shifter_in = {io_host_in_bits, T30};
  assign T30 = rx_shifter[6'h3f:5'h10];
  assign T31 = T61 ? rx_shifter_in : rx_shifter;
  assign T32 = T38 & T33;
  assign T33 = T35 | T34;
  assign T34 = cmd == 4'h3;
  assign T35 = T37 | T36;
  assign T36 = cmd == 4'h2;
  assign T37 = cmd == 4'h0;
  assign T38 = nack ^ 1'h1;
  assign nack = T54 ? bad_mem_packet : T39;
  assign T39 = T41 ? T40 : 1'h1;
  assign T40 = size != 12'h1;
  assign T41 = T43 | T42;
  assign T42 = cmd == 4'h3;
  assign T43 = cmd == 4'h2;
  assign bad_mem_packet = T52 | T44;
  assign T44 = T45 != 3'h0;
  assign T45 = addr[2'h2:1'h0];
  assign T46 = T107 ? T51 : T47;
  assign T47 = T101 ? T50 : T48;
  assign T48 = T21 ? T49 : addr;
  assign T49 = rx_shifter_in[6'h3f:5'h18];
  assign T50 = addr + 40'h8;
  assign T51 = addr + 40'h8;
  assign T52 = T53 != 3'h0;
  assign T53 = size[2'h2:1'h0];
  assign T54 = T56 | T55;
  assign T55 = cmd == 4'h1;
  assign T56 = cmd == 4'h0;
  assign tx_word_count = tx_count[4'he:2'h2];
  assign T213 = reset ? 15'h0 : T57;
  assign T57 = T26 ? 15'h0 : T58;
  assign T58 = T60 ? T59 : tx_count;
  assign T59 = tx_count + 15'h1;
  assign T60 = io_host_out_valid & io_host_out_ready;
  assign T61 = io_host_in_valid & io_host_in_ready;
  assign next_cmd = rx_shifter_in[2'h3:1'h0];
  assign T62 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T63 = rx_cmd == 4'h2;
  assign T64 = rx_cmd == 4'h1;
  assign T65 = rx_cmd == 4'h0;
  assign T66 = T78 & rx_done;
  assign rx_done = rx_word_done & T67;
  assign T67 = T75 ? T72 : T68;
  assign T68 = T71 | T69;
  assign T69 = T70 == 3'h0;
  assign T70 = rx_word_count[2'h2:1'h0];
  assign T71 = rx_word_count == T214;
  assign T214 = {1'h0, size};
  assign T72 = T74 & T73;
  assign T73 = next_cmd != 4'h3;
  assign T74 = next_cmd != 4'h1;
  assign T75 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T76;
  assign T76 = T77 == 2'h3;
  assign T77 = rx_count[1'h1:1'h0];
  assign T78 = state == 3'h0;
  assign T79 = T88 & cnt_done;
  assign cnt_done = T83 & T80;
  assign T80 = cnt == 2'h3;
  assign T215 = reset ? 2'h0 : T81;
  assign T81 = T83 ? T82 : cnt;
  assign T82 = cnt + 2'h1;
  assign T83 = T86 | T84;
  assign T84 = T85 & io_mem_grant_valid;
  assign T85 = state == 3'h5;
  assign T86 = T87 & io_mem_acquire_ready;
  assign T87 = state == 3'h4;
  assign T88 = state == 3'h4;
  assign T89 = T90 & io_mem_acquire_ready;
  assign T90 = state == 3'h3;
  assign T91 = T92 ? 3'h7 : 3'h0;
  assign T92 = T100 | T93;
  assign T93 = pos == 9'h1;
  assign T94 = T107 ? T99 : T95;
  assign T95 = T101 ? T98 : T96;
  assign T96 = T21 ? T97 : pos;
  assign T97 = rx_shifter_in[4'hf:3'h7];
  assign T98 = pos - 9'h1;
  assign T99 = pos - 9'h1;
  assign T100 = cmd == 4'h0;
  assign T101 = T102 & io_mem_grant_valid;
  assign T102 = state == 3'h6;
  assign T103 = T104 ? 3'h7 : 3'h0;
  assign T104 = T106 | T105;
  assign T105 = pos == 9'h1;
  assign T106 = cmd == 4'h0;
  assign T107 = T108 & cnt_done;
  assign T108 = state == 3'h5;
  assign T109 = T110 ? 3'h3 : 3'h0;
  assign T110 = T112 & T111;
  assign T111 = pos != 9'h0;
  assign T112 = cmd == 4'h0;
  assign T113 = T122 & tx_done;
  assign tx_done = T120 & T114;
  assign T114 = T119 | T115;
  assign T115 = T118 & T116;
  assign T116 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T117 - 3'h1;
  assign T117 = tx_word_count[2'h2:1'h0];
  assign T118 = 13'h0 < tx_word_count;
  assign T119 = tx_word_count == T216;
  assign T216 = {1'h0, tx_size};
  assign T120 = io_host_out_ready & T121;
  assign T121 = tx_subword_count == 2'h3;
  assign tx_subword_count = tx_count[1'h1:1'h0];
  assign T122 = state == 3'h7;
  assign T123 = io_cpu_0_csr_req_ready & io_cpu_0_csr_req_valid;
  assign T124 = T126 & T125;
  assign T125 = csr_addr == 12'h782;
  assign csr_addr = addr[4'hb:1'h0];
  assign T126 = T128 & T127;
  assign T127 = csr_coreid == 2'h0;
  assign csr_coreid = addr[5'h15:5'h14];
  assign T128 = state == 3'h1;
  assign T129 = T130 & io_cpu_0_csr_resp_valid;
  assign T130 = state == 3'h2;
  assign T131 = io_scr_req_ready & io_scr_req_valid;
  assign T132 = T133 & io_scr_resp_valid;
  assign T133 = state == 3'h2;
  assign T134 = {io_mem_grant_bits_addr_beat, 1'h1};
  assign T136 = io_mem_grant_bits_data[6'h3f:1'h0];
  assign T137 = T138 & io_mem_grant_valid;
  assign T138 = state == 3'h5;
  assign T139 = {io_mem_grant_bits_addr_beat, 1'h0};
  assign T141 = rx_word_done & io_host_in_ready;
  assign T142 = T143 - 3'h1;
  assign T143 = rx_word_count[2'h2:1'h0];
  assign io_scr_req_bits_addr = T144;
  assign T144 = T145;
  assign T145 = addr[3'h5:1'h0];
  assign io_scr_req_bits_rw = T146;
  assign T146 = cmd == 4'h3;
  assign io_scr_req_valid = T147;
  assign T147 = T149 & T148;
  assign T148 = csr_coreid == 2'h3;
  assign T149 = state == 3'h1;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_data = T150;
  assign T150 = T157 ? T152 : T151;
  assign T151 = 128'h0;
  assign T152 = mem_req_data;
  assign mem_req_data = {T155, T153};
  assign T153 = packet_ram[T154];
  assign T154 = {cnt, 1'h0};
  assign T155 = packet_ram[T156];
  assign T156 = {cnt, 1'h1};
  assign T157 = cmd == 4'h1;
  assign io_mem_acquire_bits_union = T158;
  assign T158 = T157 ? T160 : T159;
  assign T159 = 17'h1c1;
  assign T160 = T161;
  assign T161 = {T162, 1'h1};
  assign T162 = 16'hffff;
  assign io_mem_acquire_bits_a_type = T163;
  assign T163 = T157 ? T165 : T164;
  assign T164 = 3'h1;
  assign T165 = 3'h3;
  assign io_mem_acquire_bits_is_builtin_type = T166;
  assign T166 = T157 ? T168 : T167;
  assign T167 = 1'h1;
  assign T168 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T169;
  assign T169 = T157 ? T171 : T170;
  assign T170 = 2'h0;
  assign T171 = cnt;
  assign io_mem_acquire_bits_client_xact_id = T172;
  assign T172 = T157 ? T174 : T173;
  assign T173 = 2'h0;
  assign T174 = 2'h0;
  assign io_mem_acquire_bits_addr_block = T175;
  assign T175 = T157 ? T178 : T176;
  assign T176 = T217;
  assign T217 = init_addr[5'h19:1'h0];
  assign init_addr = T177 >> 2'h3;
  assign T177 = addr;
  assign T178 = T218;
  assign T218 = init_addr[5'h19:1'h0];
  assign io_mem_acquire_valid = T179;
  assign T179 = T181 | T180;
  assign T180 = state == 3'h4;
  assign T181 = state == 3'h3;
  assign io_cpu_0_csr_resp_ready = 1'h1;
  assign io_cpu_0_csr_req_bits_data = csr_wdata;
  assign io_cpu_0_csr_req_bits_addr = csr_addr;
  assign io_cpu_0_csr_req_bits_rw = T182;
  assign T182 = cmd == 4'h3;
  assign io_cpu_0_csr_req_valid = T183;
  assign T183 = T185 & T184;
  assign T184 = csr_addr != 12'h782;
  assign T185 = T186 & T127;
  assign T186 = state == 3'h1;
  assign io_cpu_0_reset = R187;
  assign T219 = reset ? 1'h1 : T188;
  assign T188 = T190 ? T189 : R187;
  assign T189 = csr_wdata[1'h0:1'h0];
  assign T190 = T124 & T191;
  assign T191 = cmd == 4'h3;
  assign io_host_debug_stats_csr = io_cpu_0_debug_stats_csr;
  assign io_host_out_bits = T220;
  assign T220 = T192[4'hf:1'h0];
  assign T192 = tx_data >> T193;
  assign T193 = {T194, 4'h0};
  assign T194 = tx_count[1'h1:1'h0];
  assign tx_data = T207 ? tx_header : T195;
  assign T195 = T200 ? csrReadData : T196;
  assign T196 = packet_ram[packet_ram_raddr];
  assign T197 = T132 ? io_scr_resp_bits : T198;
  assign T198 = T129 ? io_cpu_0_csr_resp_bits : T199;
  assign T199 = T124 ? T221 : csrReadData;
  assign T221 = {63'h0, R187};
  assign T200 = T202 | T201;
  assign T201 = cmd == 4'h3;
  assign T202 = cmd == 4'h2;
  assign tx_header = {T204, T203};
  assign T203 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T204 = {addr, seqno};
  assign T205 = T21 ? T206 : seqno;
  assign T206 = rx_shifter_in[5'h17:5'h10];
  assign T207 = tx_word_count == 13'h0;
  assign io_host_out_valid = T208;
  assign T208 = state == 3'h7;
  assign io_host_in_ready = T209;
  assign T209 = state == 3'h0;

  always @(posedge clk) begin
    if (T2)
      packet_ram[T134] <= T1;
    if(reset) begin
      state <= 3'h0;
    end else if(T132) begin
      state <= 3'h7;
    end else if(T131) begin
      state <= 3'h2;
    end else if(T129) begin
      state <= 3'h7;
    end else if(T124) begin
      state <= 3'h7;
    end else if(T123) begin
      state <= 3'h2;
    end else if(T113) begin
      state <= T109;
    end else if(T107) begin
      state <= T103;
    end else if(T101) begin
      state <= T91;
    end else if(T89) begin
      state <= 3'h5;
    end else if(T79) begin
      state <= 3'h6;
    end else if(T66) begin
      state <= T15;
    end
    if(T21) begin
      cmd <= next_cmd;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T26) begin
      rx_count <= 15'h0;
    end else if(T61) begin
      rx_count <= T25;
    end
    if(T21) begin
      size <= T29;
    end
    if(T61) begin
      rx_shifter <= rx_shifter_in;
    end
    if(T107) begin
      addr <= T51;
    end else if(T101) begin
      addr <= T50;
    end else if(T21) begin
      addr <= T49;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T26) begin
      tx_count <= 15'h0;
    end else if(T60) begin
      tx_count <= T59;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T83) begin
      cnt <= T82;
    end
    if(T107) begin
      pos <= T99;
    end else if(T101) begin
      pos <= T98;
    end else if(T21) begin
      pos <= T97;
    end
    if (T137)
      packet_ram[T139] <= T136;
    if (T141)
      packet_ram[T142] <= rx_shifter_in;
    if(reset) begin
      R187 <= 1'h1;
    end else if(T190) begin
      R187 <= T189;
    end
    if(T132) begin
      csrReadData <= io_scr_resp_bits;
    end else if(T129) begin
      csrReadData <= io_cpu_0_csr_resp_bits;
    end else if(T124) begin
      csrReadData <= T221;
    end
    if(T21) begin
      seqno <= T206;
    end
  end
endmodule

module ClientTileLinkIOWrapper_0(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [1:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[1:0] io_in_grant_bits_client_xact_id,
    output[2:0] io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[1:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [1:0] io_out_grant_bits_client_xact_id,
    input [2:0] io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[1:0] io_out_release_bits_client_xact_id
    //output io_out_release_bits_voluntary
    //output[2:0] io_out_release_bits_r_type
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module FinishQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_fin_manager_xact_id,
    input [1:0] io_enq_bits_dst,
    input  io_deq_ready,
    output io_deq_valid,
    output[2:0] io_deq_bits_fin_manager_xact_id,
    output[1:0] io_deq_bits_dst,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T19;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T20;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T21;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[4:0] T11;
  reg [4:0] ram [1:0];
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[2:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T19 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T20 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T21 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_dst = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_fin_manager_xact_id, io_enq_bits_dst};
  assign io_deq_bits_fin_manager_xact_id = T15;
  assign T15 = T11[3'h4:2'h2];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module FinishUnit_0(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h0;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h0;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h0;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_0 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [1:0] io_enq_bits_payload_addr_beat,
    input  io_enq_bits_payload_is_builtin_type,
    input [2:0] io_enq_bits_payload_a_type,
    input [16:0] io_enq_bits_payload_union,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[1:0] io_deq_bits_payload_addr_beat,
    output io_deq_bits_payload_is_builtin_type,
    output[2:0] io_deq_bits_payload_a_type,
    output[16:0] io_deq_bits_payload_union,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T33;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T34;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T35;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[182:0] T11;
  reg [182:0] ram [1:0];
  wire[182:0] T12;
  wire[182:0] T13;
  wire[182:0] T14;
  wire[150:0] T15;
  wire[147:0] T16;
  wire[144:0] T17;
  wire[2:0] T18;
  wire[31:0] T19;
  wire[27:0] T20;
  wire[3:0] T21;
  wire[16:0] T22;
  wire[2:0] T23;
  wire T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[25:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire empty;
  wire T31;
  wire T32;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T33 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T34 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T35 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T19, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_payload_a_type, T17};
  assign T17 = {io_enq_bits_payload_union, io_enq_bits_payload_data};
  assign T18 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_is_builtin_type};
  assign T19 = {T21, T20};
  assign T20 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_client_xact_id};
  assign T21 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_union = T22;
  assign T22 = T11[8'h90:8'h80];
  assign io_deq_bits_payload_a_type = T23;
  assign T23 = T11[8'h93:8'h91];
  assign io_deq_bits_payload_is_builtin_type = T24;
  assign T24 = T11[8'h94:8'h94];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h96:8'h95];
  assign io_deq_bits_payload_client_xact_id = T26;
  assign T26 = T11[8'h98:8'h97];
  assign io_deq_bits_payload_addr_block = T27;
  assign T27 = T11[8'hb2:8'h99];
  assign io_deq_bits_header_dst = T28;
  assign T28 = T11[8'hb4:8'hb3];
  assign io_deq_bits_header_src = T29;
  assign T29 = T11[8'hb6:8'hb5];
  assign io_deq_valid = T30;
  assign T30 = empty ^ 1'h1;
  assign empty = ptr_match & T31;
  assign T31 = maybe_full ^ 1'h1;
  assign io_enq_ready = T32;
  assign T32 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_p_type,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T23;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T24;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire[31:0] T11;
  reg [31:0] ram [1:0];
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[27:0] T15;
  wire[3:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_p_type = T10;
  assign T10 = T11[1'h1:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_payload_addr_block, io_enq_bits_payload_p_type};
  assign T16 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T11[5'h1b:2'h2];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T11[5'h1d:5'h1c];
  assign io_deq_bits_header_src = T19;
  assign T19 = T11[5'h1f:5'h1e];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input  io_enq_bits_payload_voluntary,
    input [2:0] io_enq_bits_payload_r_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output io_deq_bits_payload_voluntary,
    output[2:0] io_deq_bits_payload_r_type,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[165:0] T11;
  reg [165:0] ram [1:0];
  wire[165:0] T12;
  wire[165:0] T13;
  wire[165:0] T14;
  wire[133:0] T15;
  wire[130:0] T16;
  wire[2:0] T17;
  wire[31:0] T18;
  wire[27:0] T19;
  wire[3:0] T20;
  wire[2:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[25:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_r_type, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_voluntary};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T21;
  assign T21 = T11[8'h82:8'h80];
  assign io_deq_bits_payload_voluntary = T22;
  assign T22 = T11[8'h83:8'h83];
  assign io_deq_bits_payload_client_xact_id = T23;
  assign T23 = T11[8'h85:8'h84];
  assign io_deq_bits_payload_addr_block = T24;
  assign T24 = T11[8'h9f:8'h86];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'ha1:8'ha0];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'ha3:8'ha2];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'ha5:8'ha4];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_manager_xact_id,
    input  io_enq_bits_payload_is_builtin_type,
    input [3:0] io_enq_bits_payload_g_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_manager_xact_id,
    output io_deq_bits_payload_is_builtin_type,
    output[3:0] io_deq_bits_payload_g_type,
    output[127:0] io_deq_bits_payload_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T31;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T32;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T33;
  wire T8;
  wire T9;
  wire[127:0] T10;
  wire[143:0] T11;
  reg [143:0] ram [1:0];
  wire[143:0] T12;
  wire[143:0] T13;
  wire[143:0] T14;
  wire[135:0] T15;
  wire[131:0] T16;
  wire[3:0] T17;
  wire[7:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[2:0] T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  wire T30;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T31 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T32 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T33 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_data = T10;
  assign T10 = T11[7'h7f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_payload_g_type, io_enq_bits_payload_data};
  assign T17 = {io_enq_bits_payload_manager_xact_id, io_enq_bits_payload_is_builtin_type};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_client_xact_id};
  assign T20 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_g_type = T21;
  assign T21 = T11[8'h83:8'h80];
  assign io_deq_bits_payload_is_builtin_type = T22;
  assign T22 = T11[8'h84:8'h84];
  assign io_deq_bits_payload_manager_xact_id = T23;
  assign T23 = T11[8'h87:8'h85];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T11[8'h89:8'h88];
  assign io_deq_bits_payload_addr_beat = T25;
  assign T25 = T11[8'h8b:8'h8a];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T11[8'h8d:8'h8c];
  assign io_deq_bits_header_src = T27;
  assign T27 = T11[8'h8f:8'h8e];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign io_enq_ready = T30;
  assign T30 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_manager_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_manager_xact_id,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[2:0] T10;
  wire[6:0] T11;
  reg [6:0] ram [1:0];
  wire[6:0] T12;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[4:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_payload_manager_xact_id = T10;
  assign T10 = T11[2'h2:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_header_src, T15};
  assign T15 = {io_enq_bits_header_dst, io_enq_bits_payload_manager_xact_id};
  assign io_deq_bits_header_dst = T16;
  assign T16 = T11[3'h4:2'h3];
  assign io_deq_bits_header_src = T17;
  assign T17 = T11[3'h6:3'h5];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module TileLinkEnqueuer_0(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [1:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[1:0] io_client_grant_bits_payload_client_xact_id,
    output[2:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [2:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [1:0] io_client_release_bits_payload_client_xact_id,
    input  io_client_release_bits_payload_voluntary,
    input [2:0] io_client_release_bits_payload_r_type,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[1:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [1:0] io_manager_grant_bits_payload_client_xact_id,
    input [2:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[2:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[1:0] io_manager_release_bits_payload_client_xact_id,
    output io_manager_release_bits_payload_voluntary,
    output[2:0] io_manager_release_bits_payload_r_type,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_io_deq_bits_payload_client_xact_id;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire Queue_io_deq_bits_payload_is_builtin_type;
  wire[2:0] Queue_io_deq_bits_payload_a_type;
  wire[16:0] Queue_io_deq_bits_payload_union;
  wire[127:0] Queue_io_deq_bits_payload_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[1:0] Queue_1_io_deq_bits_header_src;
  wire[1:0] Queue_1_io_deq_bits_header_dst;
  wire[25:0] Queue_1_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_1_io_deq_bits_payload_p_type;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[1:0] Queue_2_io_deq_bits_header_src;
  wire[1:0] Queue_2_io_deq_bits_header_dst;
  wire[1:0] Queue_2_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_2_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_2_io_deq_bits_payload_client_xact_id;
  wire Queue_2_io_deq_bits_payload_voluntary;
  wire[2:0] Queue_2_io_deq_bits_payload_r_type;
  wire[127:0] Queue_2_io_deq_bits_payload_data;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_header_src;
  wire[1:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_payload_addr_beat;
  wire[1:0] Queue_3_io_deq_bits_payload_client_xact_id;
  wire[2:0] Queue_3_io_deq_bits_payload_manager_xact_id;
  wire Queue_3_io_deq_bits_payload_is_builtin_type;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire[127:0] Queue_3_io_deq_bits_payload_data;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[2:0] Queue_4_io_deq_bits_payload_manager_xact_id;


  assign io_manager_release_bits_payload_data = Queue_2_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_r_type = Queue_2_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_voluntary = Queue_2_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_2_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_2_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_2_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_2_io_deq_valid;
  assign io_manager_probe_ready = Queue_1_io_enq_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = Queue_4_io_deq_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_finish_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_finish_valid = Queue_4_io_deq_valid;
  assign io_manager_grant_ready = Queue_3_io_enq_ready;
  assign io_manager_acquire_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = Queue_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = Queue_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_acquire_valid = Queue_io_deq_valid;
  assign io_client_release_ready = Queue_2_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = Queue_1_io_deq_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = Queue_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = Queue_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_header_src = Queue_1_io_deq_bits_header_src;
  assign io_client_probe_valid = Queue_1_io_deq_valid;
  assign io_client_finish_ready = Queue_4_io_enq_ready;
  assign io_client_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_client_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_client_grant_valid = Queue_3_io_deq_valid;
  assign io_client_acquire_ready = Queue_io_enq_ready;
  Queue_9 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_acquire_valid ),
       .io_enq_bits_header_src( io_client_acquire_bits_header_src ),
       .io_enq_bits_header_dst( io_client_acquire_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_client_acquire_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_acquire_bits_payload_client_xact_id ),
       .io_enq_bits_payload_addr_beat( io_client_acquire_bits_payload_addr_beat ),
       .io_enq_bits_payload_is_builtin_type( io_client_acquire_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_a_type( io_client_acquire_bits_payload_a_type ),
       .io_enq_bits_payload_union( io_client_acquire_bits_payload_union ),
       .io_enq_bits_payload_data( io_client_acquire_bits_payload_data ),
       .io_deq_ready( io_manager_acquire_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_is_builtin_type( Queue_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_a_type( Queue_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_union( Queue_io_deq_bits_payload_union ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_10 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( io_manager_probe_valid ),
       .io_enq_bits_header_src( io_manager_probe_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_probe_bits_header_dst ),
       .io_enq_bits_payload_addr_block( io_manager_probe_bits_payload_addr_block ),
       .io_enq_bits_payload_p_type( io_manager_probe_bits_payload_p_type ),
       .io_deq_ready( io_client_probe_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_block( Queue_1_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_p_type( Queue_1_io_deq_bits_payload_p_type )
       //.io_count(  )
  );
  Queue_11 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_2_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_2_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_2_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_voluntary( Queue_2_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_r_type( Queue_2_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_data( Queue_2_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_12 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( io_manager_grant_valid ),
       .io_enq_bits_header_src( io_manager_grant_bits_header_src ),
       .io_enq_bits_header_dst( io_manager_grant_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_manager_grant_bits_payload_addr_beat ),
       .io_enq_bits_payload_client_xact_id( io_manager_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_manager_xact_id( io_manager_grant_bits_payload_manager_xact_id ),
       .io_enq_bits_payload_is_builtin_type( io_manager_grant_bits_payload_is_builtin_type ),
       .io_enq_bits_payload_g_type( io_manager_grant_bits_payload_g_type ),
       .io_enq_bits_payload_data( io_manager_grant_bits_payload_data ),
       .io_deq_ready( io_client_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_3_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_manager_xact_id( Queue_3_io_deq_bits_payload_manager_xact_id ),
       .io_deq_bits_payload_is_builtin_type( Queue_3_io_deq_bits_payload_is_builtin_type ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data )
       //.io_count(  )
  );
  Queue_13 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( io_client_finish_valid ),
       .io_enq_bits_header_src( io_client_finish_bits_header_src ),
       .io_enq_bits_header_dst( io_client_finish_bits_header_dst ),
       .io_enq_bits_payload_manager_xact_id( io_client_finish_bits_payload_manager_xact_id ),
       .io_deq_ready( io_manager_finish_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_manager_xact_id( Queue_4_io_deq_bits_payload_manager_xact_id )
       //.io_count(  )
  );
endmodule

module FinishUnit_1(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h1;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h1;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_1 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module FinishUnit_2(input clk, input reset,
    output io_grant_ready,
    input  io_grant_valid,
    input [1:0] io_grant_bits_header_src,
    input [1:0] io_grant_bits_header_dst,
    input [1:0] io_grant_bits_payload_addr_beat,
    input [1:0] io_grant_bits_payload_client_xact_id,
    input [2:0] io_grant_bits_payload_manager_xact_id,
    input  io_grant_bits_payload_is_builtin_type,
    input [3:0] io_grant_bits_payload_g_type,
    input [127:0] io_grant_bits_payload_data,
    input  io_refill_ready,
    output io_refill_valid,
    output[1:0] io_refill_bits_addr_beat,
    output[1:0] io_refill_bits_client_xact_id,
    output[2:0] io_refill_bits_manager_xact_id,
    output io_refill_bits_is_builtin_type,
    output[3:0] io_refill_bits_g_type,
    output[127:0] io_refill_bits_data,
    input  io_finish_ready,
    output io_finish_valid,
    output[1:0] io_finish_bits_header_src,
    output[1:0] io_finish_bits_header_dst,
    output[2:0] io_finish_bits_payload_manager_xact_id,
    output io_ready
);

  wire[2:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  reg [1:0] R7;
  wire[1:0] T39;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire FinishQueue_io_enq_ready;
  wire FinishQueue_io_deq_valid;
  wire[2:0] FinishQueue_io_deq_bits_fin_manager_xact_id;
  wire[1:0] FinishQueue_io_deq_bits_dst;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R7 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_grant_bits_payload_manager_xact_id;
  assign T1 = T22 & T2;
  assign T2 = T16 | T3;
  assign T3 = T11 ? T5 : T4;
  assign T4 = io_grant_ready & io_grant_valid;
  assign T5 = T10 & T6;
  assign T6 = R7 == 2'h3;
  assign T39 = reset ? 2'h0 : T8;
  assign T8 = T10 ? T9 : R7;
  assign T9 = R7 + 2'h1;
  assign T10 = T4 & T11;
  assign T11 = io_grant_bits_payload_is_builtin_type ? T15 : T12;
  assign T12 = T14 | T13;
  assign T13 = 4'h1 == io_grant_bits_payload_g_type;
  assign T14 = 4'h0 == io_grant_bits_payload_g_type;
  assign T15 = 4'h5 == io_grant_bits_payload_g_type;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_grant_bits_payload_is_builtin_type ? T21 : T18;
  assign T18 = T20 | T19;
  assign T19 = 4'h1 == io_grant_bits_payload_g_type;
  assign T20 = 4'h0 == io_grant_bits_payload_g_type;
  assign T21 = 4'h5 == io_grant_bits_payload_g_type;
  assign T22 = T26 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_grant_bits_payload_is_builtin_type & T25;
  assign T25 = io_grant_bits_payload_g_type == 4'h0;
  assign T26 = io_grant_ready & io_grant_valid;
  assign io_ready = FinishQueue_io_enq_ready;
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_io_deq_bits_fin_manager_xact_id;
  assign io_finish_bits_header_dst = FinishQueue_io_deq_bits_dst;
  assign io_finish_bits_header_src = 2'h2;
  assign io_finish_valid = FinishQueue_io_deq_valid;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_valid = T27;
  assign T27 = T28 & io_grant_valid;
  assign T28 = FinishQueue_io_enq_ready | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 ^ 1'h1;
  assign T31 = io_grant_bits_payload_is_builtin_type & T32;
  assign T32 = io_grant_bits_payload_g_type == 4'h0;
  assign io_grant_ready = T33;
  assign T33 = T34 & io_refill_ready;
  assign T34 = FinishQueue_io_enq_ready | T35;
  assign T35 = T36 ^ 1'h1;
  assign T36 = T37 ^ 1'h1;
  assign T37 = io_grant_bits_payload_is_builtin_type & T38;
  assign T38 = io_grant_bits_payload_g_type == 4'h0;
  FinishQueue FinishQueue(.clk(clk), .reset(reset),
       .io_enq_ready( FinishQueue_io_enq_ready ),
       .io_enq_valid( T1 ),
       .io_enq_bits_fin_manager_xact_id( T0 ),
       .io_enq_bits_dst( io_grant_bits_header_src ),
       .io_deq_ready( io_finish_ready ),
       .io_deq_valid( FinishQueue_io_deq_valid ),
       .io_deq_bits_fin_manager_xact_id( FinishQueue_io_deq_bits_fin_manager_xact_id ),
       .io_deq_bits_dst( FinishQueue_io_deq_bits_dst )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      R7 <= 2'h0;
    end else if(T10) begin
      R7 <= T9;
    end
  end
endmodule

module ClientTileLinkNetworkPort_2(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [25:0] io_client_acquire_bits_addr_block,
    input [1:0] io_client_acquire_bits_client_xact_id,
    input [1:0] io_client_acquire_bits_addr_beat,
    input  io_client_acquire_bits_is_builtin_type,
    input [2:0] io_client_acquire_bits_a_type,
    input [16:0] io_client_acquire_bits_union,
    input [127:0] io_client_acquire_bits_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_addr_beat,
    output[1:0] io_client_grant_bits_client_xact_id,
    output[2:0] io_client_grant_bits_manager_xact_id,
    output io_client_grant_bits_is_builtin_type,
    output[3:0] io_client_grant_bits_g_type,
    output[127:0] io_client_grant_bits_data,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[25:0] io_client_probe_bits_addr_block,
    output[1:0] io_client_probe_bits_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_addr_beat,
    input [25:0] io_client_release_bits_addr_block,
    input [1:0] io_client_release_bits_client_xact_id,
    input  io_client_release_bits_voluntary,
    input [2:0] io_client_release_bits_r_type,
    input [127:0] io_client_release_bits_data,
    input  io_network_acquire_ready,
    output io_network_acquire_valid,
    output[1:0] io_network_acquire_bits_header_src,
    output[1:0] io_network_acquire_bits_header_dst,
    output[25:0] io_network_acquire_bits_payload_addr_block,
    output[1:0] io_network_acquire_bits_payload_client_xact_id,
    output[1:0] io_network_acquire_bits_payload_addr_beat,
    output io_network_acquire_bits_payload_is_builtin_type,
    output[2:0] io_network_acquire_bits_payload_a_type,
    output[16:0] io_network_acquire_bits_payload_union,
    output[127:0] io_network_acquire_bits_payload_data,
    output io_network_grant_ready,
    input  io_network_grant_valid,
    input [1:0] io_network_grant_bits_header_src,
    input [1:0] io_network_grant_bits_header_dst,
    input [1:0] io_network_grant_bits_payload_addr_beat,
    input [1:0] io_network_grant_bits_payload_client_xact_id,
    input [2:0] io_network_grant_bits_payload_manager_xact_id,
    input  io_network_grant_bits_payload_is_builtin_type,
    input [3:0] io_network_grant_bits_payload_g_type,
    input [127:0] io_network_grant_bits_payload_data,
    input  io_network_finish_ready,
    output io_network_finish_valid,
    output[1:0] io_network_finish_bits_header_src,
    output[1:0] io_network_finish_bits_header_dst,
    output[2:0] io_network_finish_bits_payload_manager_xact_id,
    output io_network_probe_ready,
    input  io_network_probe_valid,
    input [1:0] io_network_probe_bits_header_src,
    input [1:0] io_network_probe_bits_header_dst,
    input [25:0] io_network_probe_bits_payload_addr_block,
    input [1:0] io_network_probe_bits_payload_p_type,
    input  io_network_release_ready,
    output io_network_release_valid,
    output[1:0] io_network_release_bits_header_src,
    output[1:0] io_network_release_bits_header_dst,
    output[1:0] io_network_release_bits_payload_addr_beat,
    output[25:0] io_network_release_bits_payload_addr_block,
    output[1:0] io_network_release_bits_payload_client_xact_id,
    output io_network_release_bits_payload_voluntary,
    output[2:0] io_network_release_bits_payload_r_type,
    output[127:0] io_network_release_bits_payload_data
);

  wire[127:0] rel_with_header_bits_payload_data;
  wire[2:0] rel_with_header_bits_payload_r_type;
  wire rel_with_header_bits_payload_voluntary;
  wire[1:0] rel_with_header_bits_payload_client_xact_id;
  wire[25:0] rel_with_header_bits_payload_addr_block;
  wire[1:0] rel_with_header_bits_payload_addr_beat;
  wire[1:0] rel_with_header_bits_header_dst;
  wire[1:0] rel_with_header_bits_header_src;
  wire rel_with_header_valid;
  wire prb_without_header_ready;
  wire[127:0] acq_with_header_bits_payload_data;
  wire[16:0] acq_with_header_bits_payload_union;
  wire[2:0] acq_with_header_bits_payload_a_type;
  wire acq_with_header_bits_payload_is_builtin_type;
  wire[1:0] acq_with_header_bits_payload_addr_beat;
  wire[1:0] acq_with_header_bits_payload_client_xact_id;
  wire[25:0] acq_with_header_bits_payload_addr_block;
  wire[1:0] acq_with_header_bits_header_dst;
  wire[1:0] acq_with_header_bits_header_src;
  wire T0;
  wire acq_with_header_valid;
  wire rel_with_header_ready;
  wire[1:0] prb_without_header_bits_p_type;
  wire[25:0] prb_without_header_bits_addr_block;
  wire prb_without_header_valid;
  wire acq_with_header_ready;
  wire T1;
  wire finisher_io_grant_ready;
  wire finisher_io_refill_valid;
  wire[1:0] finisher_io_refill_bits_addr_beat;
  wire[1:0] finisher_io_refill_bits_client_xact_id;
  wire[2:0] finisher_io_refill_bits_manager_xact_id;
  wire finisher_io_refill_bits_is_builtin_type;
  wire[3:0] finisher_io_refill_bits_g_type;
  wire[127:0] finisher_io_refill_bits_data;
  wire finisher_io_finish_valid;
  wire[1:0] finisher_io_finish_bits_header_src;
  wire[1:0] finisher_io_finish_bits_header_dst;
  wire[2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire finisher_io_ready;


  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign rel_with_header_bits_header_dst = 2'h0;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign rel_with_header_bits_header_src = 2'h2;
  assign io_network_release_valid = rel_with_header_valid;
  assign rel_with_header_valid = io_client_release_valid;
  assign io_network_probe_ready = prb_without_header_ready;
  assign prb_without_header_ready = io_client_probe_ready;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign acq_with_header_bits_header_dst = 2'h0;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign acq_with_header_bits_header_src = 2'h2;
  assign io_network_acquire_valid = T0;
  assign T0 = acq_with_header_valid & finisher_io_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign io_client_release_ready = rel_with_header_ready;
  assign rel_with_header_ready = io_network_release_ready;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign io_client_probe_valid = prb_without_header_valid;
  assign prb_without_header_valid = io_network_probe_valid;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign acq_with_header_ready = T1;
  assign T1 = io_network_acquire_ready & finisher_io_ready;
  FinishUnit_2 finisher(.clk(clk), .reset(reset),
       .io_grant_ready( finisher_io_grant_ready ),
       .io_grant_valid( io_network_grant_valid ),
       .io_grant_bits_header_src( io_network_grant_bits_header_src ),
       .io_grant_bits_header_dst( io_network_grant_bits_header_dst ),
       .io_grant_bits_payload_addr_beat( io_network_grant_bits_payload_addr_beat ),
       .io_grant_bits_payload_client_xact_id( io_network_grant_bits_payload_client_xact_id ),
       .io_grant_bits_payload_manager_xact_id( io_network_grant_bits_payload_manager_xact_id ),
       .io_grant_bits_payload_is_builtin_type( io_network_grant_bits_payload_is_builtin_type ),
       .io_grant_bits_payload_g_type( io_network_grant_bits_payload_g_type ),
       .io_grant_bits_payload_data( io_network_grant_bits_payload_data ),
       .io_refill_ready( io_client_grant_ready ),
       .io_refill_valid( finisher_io_refill_valid ),
       .io_refill_bits_addr_beat( finisher_io_refill_bits_addr_beat ),
       .io_refill_bits_client_xact_id( finisher_io_refill_bits_client_xact_id ),
       .io_refill_bits_manager_xact_id( finisher_io_refill_bits_manager_xact_id ),
       .io_refill_bits_is_builtin_type( finisher_io_refill_bits_is_builtin_type ),
       .io_refill_bits_g_type( finisher_io_refill_bits_g_type ),
       .io_refill_bits_data( finisher_io_refill_bits_data ),
       .io_finish_ready( io_network_finish_ready ),
       .io_finish_valid( finisher_io_finish_valid ),
       .io_finish_bits_header_src( finisher_io_finish_bits_header_src ),
       .io_finish_bits_header_dst( finisher_io_finish_bits_header_dst ),
       .io_finish_bits_payload_manager_xact_id( finisher_io_finish_bits_payload_manager_xact_id ),
       .io_ready( finisher_io_ready )
  );
endmodule

module ManagerTileLinkNetworkPort(
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[25:0] io_manager_acquire_bits_addr_block,
    output[1:0] io_manager_acquire_bits_client_xact_id,
    output[1:0] io_manager_acquire_bits_addr_beat,
    output io_manager_acquire_bits_is_builtin_type,
    output[2:0] io_manager_acquire_bits_a_type,
    output[16:0] io_manager_acquire_bits_union,
    output[127:0] io_manager_acquire_bits_data,
    output[1:0] io_manager_acquire_bits_client_id,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_addr_beat,
    input [1:0] io_manager_grant_bits_client_xact_id,
    input [2:0] io_manager_grant_bits_manager_xact_id,
    input  io_manager_grant_bits_is_builtin_type,
    input [3:0] io_manager_grant_bits_g_type,
    input [127:0] io_manager_grant_bits_data,
    input [1:0] io_manager_grant_bits_client_id,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[2:0] io_manager_finish_bits_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [25:0] io_manager_probe_bits_addr_block,
    input [1:0] io_manager_probe_bits_p_type,
    input [1:0] io_manager_probe_bits_client_id,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_addr_beat,
    output[25:0] io_manager_release_bits_addr_block,
    output[1:0] io_manager_release_bits_client_xact_id,
    output io_manager_release_bits_voluntary,
    output[2:0] io_manager_release_bits_r_type,
    output[127:0] io_manager_release_bits_data,
    output[1:0] io_manager_release_bits_client_id,
    output io_network_acquire_ready,
    input  io_network_acquire_valid,
    input [1:0] io_network_acquire_bits_header_src,
    input [1:0] io_network_acquire_bits_header_dst,
    input [25:0] io_network_acquire_bits_payload_addr_block,
    input [1:0] io_network_acquire_bits_payload_client_xact_id,
    input [1:0] io_network_acquire_bits_payload_addr_beat,
    input  io_network_acquire_bits_payload_is_builtin_type,
    input [2:0] io_network_acquire_bits_payload_a_type,
    input [16:0] io_network_acquire_bits_payload_union,
    input [127:0] io_network_acquire_bits_payload_data,
    input  io_network_grant_ready,
    output io_network_grant_valid,
    output[1:0] io_network_grant_bits_header_src,
    output[1:0] io_network_grant_bits_header_dst,
    output[1:0] io_network_grant_bits_payload_addr_beat,
    output[1:0] io_network_grant_bits_payload_client_xact_id,
    output[2:0] io_network_grant_bits_payload_manager_xact_id,
    output io_network_grant_bits_payload_is_builtin_type,
    output[3:0] io_network_grant_bits_payload_g_type,
    output[127:0] io_network_grant_bits_payload_data,
    output io_network_finish_ready,
    input  io_network_finish_valid,
    input [1:0] io_network_finish_bits_header_src,
    input [1:0] io_network_finish_bits_header_dst,
    input [2:0] io_network_finish_bits_payload_manager_xact_id,
    input  io_network_probe_ready,
    output io_network_probe_valid,
    output[1:0] io_network_probe_bits_header_src,
    output[1:0] io_network_probe_bits_header_dst,
    output[25:0] io_network_probe_bits_payload_addr_block,
    output[1:0] io_network_probe_bits_payload_p_type,
    output io_network_release_ready,
    input  io_network_release_valid,
    input [1:0] io_network_release_bits_header_src,
    input [1:0] io_network_release_bits_header_dst,
    input [1:0] io_network_release_bits_payload_addr_beat,
    input [25:0] io_network_release_bits_payload_addr_block,
    input [1:0] io_network_release_bits_payload_client_xact_id,
    input  io_network_release_bits_payload_voluntary,
    input [2:0] io_network_release_bits_payload_r_type,
    input [127:0] io_network_release_bits_payload_data
);

  wire T0;
  wire[1:0] T1;
  wire[25:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire[127:0] T7;
  wire[3:0] T8;
  wire T9;
  wire[2:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire[1:0] T14;
  wire T15;
  wire T16;
  wire[127:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire[127:0] T28;
  wire[16:0] T29;
  wire[2:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[25:0] T34;
  wire T35;


  assign io_network_release_ready = T0;
  assign T0 = io_manager_release_ready;
  assign io_network_probe_bits_payload_p_type = T1;
  assign T1 = io_manager_probe_bits_p_type;
  assign io_network_probe_bits_payload_addr_block = T2;
  assign T2 = io_manager_probe_bits_addr_block;
  assign io_network_probe_bits_header_dst = T3;
  assign T3 = io_manager_probe_bits_client_id;
  assign io_network_probe_bits_header_src = T4;
  assign T4 = 2'h0;
  assign io_network_probe_valid = T5;
  assign T5 = io_manager_probe_valid;
  assign io_network_finish_ready = T6;
  assign T6 = io_manager_finish_ready;
  assign io_network_grant_bits_payload_data = T7;
  assign T7 = io_manager_grant_bits_data;
  assign io_network_grant_bits_payload_g_type = T8;
  assign T8 = io_manager_grant_bits_g_type;
  assign io_network_grant_bits_payload_is_builtin_type = T9;
  assign T9 = io_manager_grant_bits_is_builtin_type;
  assign io_network_grant_bits_payload_manager_xact_id = T10;
  assign T10 = io_manager_grant_bits_manager_xact_id;
  assign io_network_grant_bits_payload_client_xact_id = T11;
  assign T11 = io_manager_grant_bits_client_xact_id;
  assign io_network_grant_bits_payload_addr_beat = T12;
  assign T12 = io_manager_grant_bits_addr_beat;
  assign io_network_grant_bits_header_dst = T13;
  assign T13 = io_manager_grant_bits_client_id;
  assign io_network_grant_bits_header_src = T14;
  assign T14 = 2'h0;
  assign io_network_grant_valid = T15;
  assign T15 = io_manager_grant_valid;
  assign io_network_acquire_ready = T16;
  assign T16 = io_manager_acquire_ready;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src;
  assign io_manager_release_bits_data = T17;
  assign T17 = io_network_release_bits_payload_data;
  assign io_manager_release_bits_r_type = T18;
  assign T18 = io_network_release_bits_payload_r_type;
  assign io_manager_release_bits_voluntary = T19;
  assign T19 = io_network_release_bits_payload_voluntary;
  assign io_manager_release_bits_client_xact_id = T20;
  assign T20 = io_network_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_addr_block = T21;
  assign T21 = io_network_release_bits_payload_addr_block;
  assign io_manager_release_bits_addr_beat = T22;
  assign T22 = io_network_release_bits_payload_addr_beat;
  assign io_manager_release_valid = T23;
  assign T23 = io_network_release_valid;
  assign io_manager_probe_ready = T24;
  assign T24 = io_network_probe_ready;
  assign io_manager_finish_bits_manager_xact_id = T25;
  assign T25 = io_network_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_valid = T26;
  assign T26 = io_network_finish_valid;
  assign io_manager_grant_ready = T27;
  assign T27 = io_network_grant_ready;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src;
  assign io_manager_acquire_bits_data = T28;
  assign T28 = io_network_acquire_bits_payload_data;
  assign io_manager_acquire_bits_union = T29;
  assign T29 = io_network_acquire_bits_payload_union;
  assign io_manager_acquire_bits_a_type = T30;
  assign T30 = io_network_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_is_builtin_type = T31;
  assign T31 = io_network_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_addr_beat = T32;
  assign T32 = io_network_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_client_xact_id = T33;
  assign T33 = io_network_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_addr_block = T34;
  assign T34 = io_network_acquire_bits_payload_addr_block;
  assign io_manager_acquire_valid = T35;
  assign T35 = io_network_acquire_valid;
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [1:0] io_enq_bits_payload_addr_beat,
    input [25:0] io_enq_bits_payload_addr_block,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input  io_enq_bits_payload_voluntary,
    input [2:0] io_enq_bits_payload_r_type,
    input [127:0] io_enq_bits_payload_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[1:0] io_deq_bits_payload_addr_beat,
    output[25:0] io_deq_bits_payload_addr_block,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output io_deq_bits_payload_voluntary,
    output[2:0] io_deq_bits_payload_r_type,
    output[127:0] io_deq_bits_payload_data,
    output io_count
);

  wire T23;
  wire[1:0] T0;
  reg  full;
  wire T24;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[165:0] T4;
  reg [165:0] ram [0:0];
  wire[165:0] T5;
  wire[165:0] T6;
  wire[165:0] T7;
  wire[133:0] T8;
  wire[130:0] T9;
  wire[2:0] T10;
  wire[31:0] T11;
  wire[27:0] T12;
  wire[3:0] T13;
  wire[2:0] T14;
  wire T15;
  wire[1:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire empty;
  wire T22;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {6{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T23;
  assign T23 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T24 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {io_enq_bits_payload_r_type, io_enq_bits_payload_data};
  assign T10 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_voluntary};
  assign T11 = {T13, T12};
  assign T12 = {io_enq_bits_payload_addr_beat, io_enq_bits_payload_addr_block};
  assign T13 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign io_deq_bits_payload_r_type = T14;
  assign T14 = T4[8'h82:8'h80];
  assign io_deq_bits_payload_voluntary = T15;
  assign T15 = T4[8'h83:8'h83];
  assign io_deq_bits_payload_client_xact_id = T16;
  assign T16 = T4[8'h85:8'h84];
  assign io_deq_bits_payload_addr_block = T17;
  assign T17 = T4[8'h9f:8'h86];
  assign io_deq_bits_payload_addr_beat = T18;
  assign T18 = T4[8'ha1:8'ha0];
  assign io_deq_bits_header_dst = T19;
  assign T19 = T4[8'ha3:8'ha2];
  assign io_deq_bits_header_src = T20;
  assign T20 = T4[8'ha5:8'ha4];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module TileLinkEnqueuer_1(input clk, input reset,
    output io_client_acquire_ready,
    input  io_client_acquire_valid,
    input [1:0] io_client_acquire_bits_header_src,
    input [1:0] io_client_acquire_bits_header_dst,
    input [25:0] io_client_acquire_bits_payload_addr_block,
    input [1:0] io_client_acquire_bits_payload_client_xact_id,
    input [1:0] io_client_acquire_bits_payload_addr_beat,
    input  io_client_acquire_bits_payload_is_builtin_type,
    input [2:0] io_client_acquire_bits_payload_a_type,
    input [16:0] io_client_acquire_bits_payload_union,
    input [127:0] io_client_acquire_bits_payload_data,
    input  io_client_grant_ready,
    output io_client_grant_valid,
    output[1:0] io_client_grant_bits_header_src,
    output[1:0] io_client_grant_bits_header_dst,
    output[1:0] io_client_grant_bits_payload_addr_beat,
    output[1:0] io_client_grant_bits_payload_client_xact_id,
    output[2:0] io_client_grant_bits_payload_manager_xact_id,
    output io_client_grant_bits_payload_is_builtin_type,
    output[3:0] io_client_grant_bits_payload_g_type,
    output[127:0] io_client_grant_bits_payload_data,
    output io_client_finish_ready,
    input  io_client_finish_valid,
    input [1:0] io_client_finish_bits_header_src,
    input [1:0] io_client_finish_bits_header_dst,
    input [2:0] io_client_finish_bits_payload_manager_xact_id,
    input  io_client_probe_ready,
    output io_client_probe_valid,
    output[1:0] io_client_probe_bits_header_src,
    output[1:0] io_client_probe_bits_header_dst,
    output[25:0] io_client_probe_bits_payload_addr_block,
    output[1:0] io_client_probe_bits_payload_p_type,
    output io_client_release_ready,
    input  io_client_release_valid,
    input [1:0] io_client_release_bits_header_src,
    input [1:0] io_client_release_bits_header_dst,
    input [1:0] io_client_release_bits_payload_addr_beat,
    input [25:0] io_client_release_bits_payload_addr_block,
    input [1:0] io_client_release_bits_payload_client_xact_id,
    input  io_client_release_bits_payload_voluntary,
    input [2:0] io_client_release_bits_payload_r_type,
    input [127:0] io_client_release_bits_payload_data,
    input  io_manager_acquire_ready,
    output io_manager_acquire_valid,
    output[1:0] io_manager_acquire_bits_header_src,
    output[1:0] io_manager_acquire_bits_header_dst,
    output[25:0] io_manager_acquire_bits_payload_addr_block,
    output[1:0] io_manager_acquire_bits_payload_client_xact_id,
    output[1:0] io_manager_acquire_bits_payload_addr_beat,
    output io_manager_acquire_bits_payload_is_builtin_type,
    output[2:0] io_manager_acquire_bits_payload_a_type,
    output[16:0] io_manager_acquire_bits_payload_union,
    output[127:0] io_manager_acquire_bits_payload_data,
    output io_manager_grant_ready,
    input  io_manager_grant_valid,
    input [1:0] io_manager_grant_bits_header_src,
    input [1:0] io_manager_grant_bits_header_dst,
    input [1:0] io_manager_grant_bits_payload_addr_beat,
    input [1:0] io_manager_grant_bits_payload_client_xact_id,
    input [2:0] io_manager_grant_bits_payload_manager_xact_id,
    input  io_manager_grant_bits_payload_is_builtin_type,
    input [3:0] io_manager_grant_bits_payload_g_type,
    input [127:0] io_manager_grant_bits_payload_data,
    input  io_manager_finish_ready,
    output io_manager_finish_valid,
    output[1:0] io_manager_finish_bits_header_src,
    output[1:0] io_manager_finish_bits_header_dst,
    output[2:0] io_manager_finish_bits_payload_manager_xact_id,
    output io_manager_probe_ready,
    input  io_manager_probe_valid,
    input [1:0] io_manager_probe_bits_header_src,
    input [1:0] io_manager_probe_bits_header_dst,
    input [25:0] io_manager_probe_bits_payload_addr_block,
    input [1:0] io_manager_probe_bits_payload_p_type,
    input  io_manager_release_ready,
    output io_manager_release_valid,
    output[1:0] io_manager_release_bits_header_src,
    output[1:0] io_manager_release_bits_header_dst,
    output[1:0] io_manager_release_bits_payload_addr_beat,
    output[25:0] io_manager_release_bits_payload_addr_block,
    output[1:0] io_manager_release_bits_payload_client_xact_id,
    output io_manager_release_bits_payload_voluntary,
    output[2:0] io_manager_release_bits_payload_r_type,
    output[127:0] io_manager_release_bits_payload_data
);

  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[1:0] Queue_io_deq_bits_header_src;
  wire[1:0] Queue_io_deq_bits_header_dst;
  wire[1:0] Queue_io_deq_bits_payload_addr_beat;
  wire[25:0] Queue_io_deq_bits_payload_addr_block;
  wire[1:0] Queue_io_deq_bits_payload_client_xact_id;
  wire Queue_io_deq_bits_payload_voluntary;
  wire[2:0] Queue_io_deq_bits_payload_r_type;
  wire[127:0] Queue_io_deq_bits_payload_data;


  assign io_manager_release_bits_payload_data = Queue_io_deq_bits_payload_data;
  assign io_manager_release_bits_payload_r_type = Queue_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_voluntary = Queue_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_client_xact_id = Queue_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_addr_block = Queue_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_addr_beat = Queue_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_header_dst = Queue_io_deq_bits_header_dst;
  assign io_manager_release_bits_header_src = Queue_io_deq_bits_header_src;
  assign io_manager_release_valid = Queue_io_deq_valid;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_client_release_ready = Queue_io_enq_ready;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_acquire_ready = io_manager_acquire_ready;
  Queue_14 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_client_release_valid ),
       .io_enq_bits_header_src( io_client_release_bits_header_src ),
       .io_enq_bits_header_dst( io_client_release_bits_header_dst ),
       .io_enq_bits_payload_addr_beat( io_client_release_bits_payload_addr_beat ),
       .io_enq_bits_payload_addr_block( io_client_release_bits_payload_addr_block ),
       .io_enq_bits_payload_client_xact_id( io_client_release_bits_payload_client_xact_id ),
       .io_enq_bits_payload_voluntary( io_client_release_bits_payload_voluntary ),
       .io_enq_bits_payload_r_type( io_client_release_bits_payload_r_type ),
       .io_enq_bits_payload_data( io_client_release_bits_payload_data ),
       .io_deq_ready( io_manager_release_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_header_src( Queue_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr_beat( Queue_io_deq_bits_payload_addr_beat ),
       .io_deq_bits_payload_addr_block( Queue_io_deq_bits_payload_addr_block ),
       .io_deq_bits_payload_client_xact_id( Queue_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_voluntary( Queue_io_deq_bits_payload_voluntary ),
       .io_deq_bits_payload_r_type( Queue_io_deq_bits_payload_r_type ),
       .io_deq_bits_payload_data( Queue_io_deq_bits_payload_data )
       //.io_count(  )
  );
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input  io_in_2_bits_payload_is_builtin_type,
    input [2:0] io_in_2_bits_payload_a_type,
    input [16:0] io_in_2_bits_payload_union,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input  io_in_1_bits_payload_is_builtin_type,
    input [2:0] io_in_1_bits_payload_a_type,
    input [16:0] io_in_1_bits_payload_union,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input  io_in_0_bits_payload_is_builtin_type,
    input [2:0] io_in_0_bits_payload_a_type,
    input [16:0] io_in_0_bits_payload_union,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr_block,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[1:0] io_out_bits_payload_addr_beat,
    output io_out_bits_payload_is_builtin_type,
    output[2:0] io_out_bits_payload_a_type,
    output[16:0] io_out_bits_payload_union,
    output[127:0] io_out_bits_payload_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T107;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T108;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg  locked;
  wire T109;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  reg [1:0] R26;
  wire[1:0] T110;
  wire[1:0] T27;
  wire[127:0] T28;
  wire[127:0] T29;
  wire T30;
  wire[1:0] T31;
  wire T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire T35;
  wire T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire[25:0] T53;
  wire[25:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R26 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T107 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T108 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T20 & T18;
  assign T18 = io_out_bits_payload_is_builtin_type & T19;
  assign T19 = 3'h3 == io_out_bits_payload_a_type;
  assign T20 = io_out_ready & io_out_valid;
  assign T109 = reset ? 1'h0 : T21;
  assign T21 = T23 ? 1'h0 : T22;
  assign T22 = T15 ? 1'h1 : locked;
  assign T23 = T20 & T24;
  assign T24 = T25 == 2'h0;
  assign T25 = R26 + 2'h1;
  assign T110 = reset ? 2'h0 : T27;
  assign T27 = T17 ? T25 : R26;
  assign io_out_bits_payload_data = T28;
  assign T28 = T32 ? io_in_2_bits_payload_data : T29;
  assign T29 = T30 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T30 = T31[1'h0:1'h0];
  assign T31 = chosen;
  assign T32 = T31[1'h1:1'h1];
  assign io_out_bits_payload_union = T33;
  assign T33 = T36 ? io_in_2_bits_payload_union : T34;
  assign T34 = T35 ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign T35 = T31[1'h0:1'h0];
  assign T36 = T31[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T37;
  assign T37 = T40 ? io_in_2_bits_payload_a_type : T38;
  assign T38 = T39 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T39 = T31[1'h0:1'h0];
  assign T40 = T31[1'h1:1'h1];
  assign io_out_bits_payload_is_builtin_type = T41;
  assign T41 = T44 ? io_in_2_bits_payload_is_builtin_type : T42;
  assign T42 = T43 ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign T43 = T31[1'h0:1'h0];
  assign T44 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T45;
  assign T45 = T48 ? io_in_2_bits_payload_addr_beat : T46;
  assign T46 = T47 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T47 = T31[1'h0:1'h0];
  assign T48 = T31[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T49;
  assign T49 = T52 ? io_in_2_bits_payload_client_xact_id : T50;
  assign T50 = T51 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T51 = T31[1'h0:1'h0];
  assign T52 = T31[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T53;
  assign T53 = T56 ? io_in_2_bits_payload_addr_block : T54;
  assign T54 = T55 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T55 = T31[1'h0:1'h0];
  assign T56 = T31[1'h1:1'h1];
  assign io_out_bits_header_dst = T57;
  assign T57 = T60 ? io_in_2_bits_header_dst : T58;
  assign T58 = T59 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T59 = T31[1'h0:1'h0];
  assign T60 = T31[1'h1:1'h1];
  assign io_out_bits_header_src = T61;
  assign T61 = T64 ? io_in_2_bits_header_src : T62;
  assign T62 = T63 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T63 = T31[1'h0:1'h0];
  assign T64 = T31[1'h1:1'h1];
  assign io_out_valid = T65;
  assign T65 = T68 ? io_in_2_valid : T66;
  assign T66 = T67 ? io_in_1_valid : io_in_0_valid;
  assign T67 = T31[1'h0:1'h0];
  assign T68 = T31[1'h1:1'h1];
  assign io_in_0_ready = T69;
  assign T69 = T70 & io_out_ready;
  assign T70 = locked ? T82 : T71;
  assign T71 = T81 | T72;
  assign T72 = T73 ^ 1'h1;
  assign T73 = T76 | T74;
  assign T74 = io_in_2_valid & T75;
  assign T75 = last_grant < 2'h2;
  assign T76 = T79 | T77;
  assign T77 = io_in_1_valid & T78;
  assign T78 = last_grant < 2'h1;
  assign T79 = io_in_0_valid & T80;
  assign T80 = last_grant < 2'h0;
  assign T81 = last_grant < 2'h0;
  assign T82 = lockIdx == 2'h0;
  assign io_in_1_ready = T83;
  assign T83 = T84 & io_out_ready;
  assign T84 = locked ? T93 : T85;
  assign T85 = T90 | T86;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | io_in_0_valid;
  assign T88 = T89 | T74;
  assign T89 = T79 | T77;
  assign T90 = T92 & T91;
  assign T91 = last_grant < 2'h1;
  assign T92 = T79 ^ 1'h1;
  assign T93 = lockIdx == 2'h1;
  assign io_in_2_ready = T94;
  assign T94 = T95 & io_out_ready;
  assign T95 = locked ? T106 : T96;
  assign T96 = T102 | T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T99 | io_in_1_valid;
  assign T99 = T100 | io_in_0_valid;
  assign T100 = T101 | T74;
  assign T101 = T79 | T77;
  assign T102 = T104 & T103;
  assign T103 = last_grant < 2'h2;
  assign T104 = T105 ^ 1'h1;
  assign T105 = T79 | T77;
  assign T106 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T23) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R26 <= 2'h0;
    end else if(T17) begin
      R26 <= T25;
    end
  end
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [1:0] io_in_2_bits_payload_addr_beat,
    input [25:0] io_in_2_bits_payload_addr_block,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input  io_in_2_bits_payload_voluntary,
    input [2:0] io_in_2_bits_payload_r_type,
    input [127:0] io_in_2_bits_payload_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [1:0] io_in_1_bits_payload_addr_beat,
    input [25:0] io_in_1_bits_payload_addr_block,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input  io_in_1_bits_payload_voluntary,
    input [2:0] io_in_1_bits_payload_r_type,
    input [127:0] io_in_1_bits_payload_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [1:0] io_in_0_bits_payload_addr_beat,
    input [25:0] io_in_0_bits_payload_addr_block,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input  io_in_0_bits_payload_voluntary,
    input [2:0] io_in_0_bits_payload_r_type,
    input [127:0] io_in_0_bits_payload_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[1:0] io_out_bits_payload_addr_beat,
    output[25:0] io_out_bits_payload_addr_block,
    output[1:0] io_out_bits_payload_client_xact_id,
    output io_out_bits_payload_voluntary,
    output[2:0] io_out_bits_payload_r_type,
    output[127:0] io_out_bits_payload_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T106;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  reg [1:0] lockIdx;
  wire[1:0] T107;
  wire[1:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  reg  locked;
  wire T108;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  reg [1:0] R29;
  wire[1:0] T109;
  wire[1:0] T30;
  wire[127:0] T31;
  wire[127:0] T32;
  wire T33;
  wire[1:0] T34;
  wire T35;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire[25:0] T48;
  wire[25:0] T49;
  wire T50;
  wire T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R29 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T8 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T106 = reset ? 2'h0 : T6;
  assign T6 = T7 ? chosen : last_grant;
  assign T7 = io_out_ready & io_out_valid;
  assign T8 = io_in_1_valid & T9;
  assign T9 = last_grant < 2'h1;
  assign T107 = reset ? 2'h2 : T10;
  assign T10 = T15 ? T11 : lockIdx;
  assign T11 = T14 ? 2'h0 : T12;
  assign T12 = T13 ? 2'h1 : 2'h2;
  assign T13 = io_in_1_ready & io_in_1_valid;
  assign T14 = io_in_0_ready & io_in_0_valid;
  assign T15 = T17 & T16;
  assign T16 = locked ^ 1'h1;
  assign T17 = T23 & T18;
  assign T18 = T20 | T19;
  assign T19 = 3'h2 == io_out_bits_payload_r_type;
  assign T20 = T22 | T21;
  assign T21 = 3'h1 == io_out_bits_payload_r_type;
  assign T22 = 3'h0 == io_out_bits_payload_r_type;
  assign T23 = io_out_ready & io_out_valid;
  assign T108 = reset ? 1'h0 : T24;
  assign T24 = T26 ? 1'h0 : T25;
  assign T25 = T15 ? 1'h1 : locked;
  assign T26 = T23 & T27;
  assign T27 = T28 == 2'h0;
  assign T28 = R29 + 2'h1;
  assign T109 = reset ? 2'h0 : T30;
  assign T30 = T17 ? T28 : R29;
  assign io_out_bits_payload_data = T31;
  assign T31 = T35 ? io_in_2_bits_payload_data : T32;
  assign T32 = T33 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T33 = T34[1'h0:1'h0];
  assign T34 = chosen;
  assign T35 = T34[1'h1:1'h1];
  assign io_out_bits_payload_r_type = T36;
  assign T36 = T39 ? io_in_2_bits_payload_r_type : T37;
  assign T37 = T38 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T38 = T34[1'h0:1'h0];
  assign T39 = T34[1'h1:1'h1];
  assign io_out_bits_payload_voluntary = T40;
  assign T40 = T43 ? io_in_2_bits_payload_voluntary : T41;
  assign T41 = T42 ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign T42 = T34[1'h0:1'h0];
  assign T43 = T34[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T44;
  assign T44 = T47 ? io_in_2_bits_payload_client_xact_id : T45;
  assign T45 = T46 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T46 = T34[1'h0:1'h0];
  assign T47 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_block = T48;
  assign T48 = T51 ? io_in_2_bits_payload_addr_block : T49;
  assign T49 = T50 ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign T50 = T34[1'h0:1'h0];
  assign T51 = T34[1'h1:1'h1];
  assign io_out_bits_payload_addr_beat = T52;
  assign T52 = T55 ? io_in_2_bits_payload_addr_beat : T53;
  assign T53 = T54 ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign T54 = T34[1'h0:1'h0];
  assign T55 = T34[1'h1:1'h1];
  assign io_out_bits_header_dst = T56;
  assign T56 = T59 ? io_in_2_bits_header_dst : T57;
  assign T57 = T58 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T58 = T34[1'h0:1'h0];
  assign T59 = T34[1'h1:1'h1];
  assign io_out_bits_header_src = T60;
  assign T60 = T63 ? io_in_2_bits_header_src : T61;
  assign T61 = T62 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T62 = T34[1'h0:1'h0];
  assign T63 = T34[1'h1:1'h1];
  assign io_out_valid = T64;
  assign T64 = T67 ? io_in_2_valid : T65;
  assign T65 = T66 ? io_in_1_valid : io_in_0_valid;
  assign T66 = T34[1'h0:1'h0];
  assign T67 = T34[1'h1:1'h1];
  assign io_in_0_ready = T68;
  assign T68 = T69 & io_out_ready;
  assign T69 = locked ? T81 : T70;
  assign T70 = T80 | T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T75 | T73;
  assign T73 = io_in_2_valid & T74;
  assign T74 = last_grant < 2'h2;
  assign T75 = T78 | T76;
  assign T76 = io_in_1_valid & T77;
  assign T77 = last_grant < 2'h1;
  assign T78 = io_in_0_valid & T79;
  assign T79 = last_grant < 2'h0;
  assign T80 = last_grant < 2'h0;
  assign T81 = lockIdx == 2'h0;
  assign io_in_1_ready = T82;
  assign T82 = T83 & io_out_ready;
  assign T83 = locked ? T92 : T84;
  assign T84 = T89 | T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T87 | io_in_0_valid;
  assign T87 = T88 | T73;
  assign T88 = T78 | T76;
  assign T89 = T91 & T90;
  assign T90 = last_grant < 2'h1;
  assign T91 = T78 ^ 1'h1;
  assign T92 = lockIdx == 2'h1;
  assign io_in_2_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = locked ? T105 : T95;
  assign T95 = T101 | T96;
  assign T96 = T97 ^ 1'h1;
  assign T97 = T98 | io_in_1_valid;
  assign T98 = T99 | io_in_0_valid;
  assign T99 = T100 | T73;
  assign T100 = T78 | T76;
  assign T101 = T103 & T102;
  assign T102 = last_grant < 2'h2;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T78 | T76;
  assign T105 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T7) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T15) begin
      lockIdx <= T11;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T26) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R29 <= 2'h0;
    end else if(T17) begin
      R29 <= T28;
    end
  end
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_manager_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_manager_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_manager_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_manager_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire T3;
  wire T4;
  reg [1:0] last_grant;
  wire[1:0] T58;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T7 ? 2'h1 : T0;
  assign T0 = T3 ? 2'h2 : T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T3 = io_in_2_valid & T4;
  assign T4 = last_grant < 2'h2;
  assign T58 = reset ? 2'h0 : T5;
  assign T5 = T6 ? chosen : last_grant;
  assign T6 = io_out_ready & io_out_valid;
  assign T7 = io_in_1_valid & T8;
  assign T8 = last_grant < 2'h1;
  assign io_out_bits_payload_manager_xact_id = T9;
  assign T9 = T13 ? io_in_2_bits_payload_manager_xact_id : T10;
  assign T10 = T11 ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = chosen;
  assign T13 = T12[1'h1:1'h1];
  assign io_out_bits_header_dst = T14;
  assign T14 = T17 ? io_in_2_bits_header_dst : T15;
  assign T15 = T16 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T16 = T12[1'h0:1'h0];
  assign T17 = T12[1'h1:1'h1];
  assign io_out_bits_header_src = T18;
  assign T18 = T21 ? io_in_2_bits_header_src : T19;
  assign T19 = T20 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign io_out_valid = T22;
  assign T22 = T25 ? io_in_2_valid : T23;
  assign T23 = T24 ? io_in_1_valid : io_in_0_valid;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T12[1'h1:1'h1];
  assign io_in_0_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T37 | T28;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T32 | T30;
  assign T30 = io_in_2_valid & T31;
  assign T31 = last_grant < 2'h2;
  assign T32 = T35 | T33;
  assign T33 = io_in_1_valid & T34;
  assign T34 = last_grant < 2'h1;
  assign T35 = io_in_0_valid & T36;
  assign T36 = last_grant < 2'h0;
  assign T37 = last_grant < 2'h0;
  assign io_in_1_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T44 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T42 | io_in_0_valid;
  assign T42 = T43 | T30;
  assign T43 = T35 | T33;
  assign T44 = T46 & T45;
  assign T45 = last_grant < 2'h1;
  assign T46 = T35 ^ 1'h1;
  assign io_in_2_ready = T47;
  assign T47 = T48 & io_out_ready;
  assign T48 = T54 | T49;
  assign T49 = T50 ^ 1'h1;
  assign T50 = T51 | io_in_1_valid;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T30;
  assign T53 = T35 | T33;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h2;
  assign T56 = T57 ^ 1'h1;
  assign T57 = T35 | T33;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T6) begin
      last_grant <= chosen;
    end
  end
endmodule

module RocketChipTileLinkArbiter(input clk, input reset,
    output io_clients_2_acquire_ready,
    input  io_clients_2_acquire_valid,
    input [25:0] io_clients_2_acquire_bits_addr_block,
    input [1:0] io_clients_2_acquire_bits_client_xact_id,
    input [1:0] io_clients_2_acquire_bits_addr_beat,
    input  io_clients_2_acquire_bits_is_builtin_type,
    input [2:0] io_clients_2_acquire_bits_a_type,
    input [16:0] io_clients_2_acquire_bits_union,
    input [127:0] io_clients_2_acquire_bits_data,
    input  io_clients_2_grant_ready,
    output io_clients_2_grant_valid,
    output[1:0] io_clients_2_grant_bits_addr_beat,
    output[1:0] io_clients_2_grant_bits_client_xact_id,
    output[2:0] io_clients_2_grant_bits_manager_xact_id,
    output io_clients_2_grant_bits_is_builtin_type,
    output[3:0] io_clients_2_grant_bits_g_type,
    output[127:0] io_clients_2_grant_bits_data,
    input  io_clients_2_probe_ready,
    output io_clients_2_probe_valid,
    output[25:0] io_clients_2_probe_bits_addr_block,
    output[1:0] io_clients_2_probe_bits_p_type,
    output io_clients_2_release_ready,
    input  io_clients_2_release_valid,
    input [1:0] io_clients_2_release_bits_addr_beat,
    input [25:0] io_clients_2_release_bits_addr_block,
    input [1:0] io_clients_2_release_bits_client_xact_id,
    input  io_clients_2_release_bits_voluntary,
    input [2:0] io_clients_2_release_bits_r_type,
    input [127:0] io_clients_2_release_bits_data,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [25:0] io_clients_1_acquire_bits_addr_block,
    input [1:0] io_clients_1_acquire_bits_client_xact_id,
    input [1:0] io_clients_1_acquire_bits_addr_beat,
    input  io_clients_1_acquire_bits_is_builtin_type,
    input [2:0] io_clients_1_acquire_bits_a_type,
    input [16:0] io_clients_1_acquire_bits_union,
    input [127:0] io_clients_1_acquire_bits_data,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_addr_beat,
    output[1:0] io_clients_1_grant_bits_client_xact_id,
    output[2:0] io_clients_1_grant_bits_manager_xact_id,
    output io_clients_1_grant_bits_is_builtin_type,
    output[3:0] io_clients_1_grant_bits_g_type,
    output[127:0] io_clients_1_grant_bits_data,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[25:0] io_clients_1_probe_bits_addr_block,
    output[1:0] io_clients_1_probe_bits_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_addr_beat,
    input [25:0] io_clients_1_release_bits_addr_block,
    input [1:0] io_clients_1_release_bits_client_xact_id,
    input  io_clients_1_release_bits_voluntary,
    input [2:0] io_clients_1_release_bits_r_type,
    input [127:0] io_clients_1_release_bits_data,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [25:0] io_clients_0_acquire_bits_addr_block,
    input [1:0] io_clients_0_acquire_bits_client_xact_id,
    input [1:0] io_clients_0_acquire_bits_addr_beat,
    input  io_clients_0_acquire_bits_is_builtin_type,
    input [2:0] io_clients_0_acquire_bits_a_type,
    input [16:0] io_clients_0_acquire_bits_union,
    input [127:0] io_clients_0_acquire_bits_data,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_addr_beat,
    output[1:0] io_clients_0_grant_bits_client_xact_id,
    output[2:0] io_clients_0_grant_bits_manager_xact_id,
    output io_clients_0_grant_bits_is_builtin_type,
    output[3:0] io_clients_0_grant_bits_g_type,
    output[127:0] io_clients_0_grant_bits_data,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[25:0] io_clients_0_probe_bits_addr_block,
    output[1:0] io_clients_0_probe_bits_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_addr_beat,
    input [25:0] io_clients_0_release_bits_addr_block,
    input [1:0] io_clients_0_release_bits_client_xact_id,
    input  io_clients_0_release_bits_voluntary,
    input [2:0] io_clients_0_release_bits_r_type,
    input [127:0] io_clients_0_release_bits_data,
    input  io_managers_0_acquire_ready,
    output io_managers_0_acquire_valid,
    output[25:0] io_managers_0_acquire_bits_addr_block,
    output[1:0] io_managers_0_acquire_bits_client_xact_id,
    output[1:0] io_managers_0_acquire_bits_addr_beat,
    output io_managers_0_acquire_bits_is_builtin_type,
    output[2:0] io_managers_0_acquire_bits_a_type,
    output[16:0] io_managers_0_acquire_bits_union,
    output[127:0] io_managers_0_acquire_bits_data,
    output[1:0] io_managers_0_acquire_bits_client_id,
    output io_managers_0_grant_ready,
    input  io_managers_0_grant_valid,
    input [1:0] io_managers_0_grant_bits_addr_beat,
    input [1:0] io_managers_0_grant_bits_client_xact_id,
    input [2:0] io_managers_0_grant_bits_manager_xact_id,
    input  io_managers_0_grant_bits_is_builtin_type,
    input [3:0] io_managers_0_grant_bits_g_type,
    input [127:0] io_managers_0_grant_bits_data,
    input [1:0] io_managers_0_grant_bits_client_id,
    input  io_managers_0_finish_ready,
    output io_managers_0_finish_valid,
    output[2:0] io_managers_0_finish_bits_manager_xact_id,
    output io_managers_0_probe_ready,
    input  io_managers_0_probe_valid,
    input [25:0] io_managers_0_probe_bits_addr_block,
    input [1:0] io_managers_0_probe_bits_p_type,
    input [1:0] io_managers_0_probe_bits_client_id,
    input  io_managers_0_release_ready,
    output io_managers_0_release_valid,
    output[1:0] io_managers_0_release_bits_addr_beat,
    output[25:0] io_managers_0_release_bits_addr_block,
    output[1:0] io_managers_0_release_bits_client_xact_id,
    output io_managers_0_release_bits_voluntary,
    output[2:0] io_managers_0_release_bits_r_type,
    output[127:0] io_managers_0_release_bits_data,
    output[1:0] io_managers_0_release_bits_client_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  wire ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  wire[16:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_manager_grant_ready;
  wire ManagerTileLinkNetworkPort_io_manager_finish_valid;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_probe_ready;
  wire ManagerTileLinkNetworkPort_io_manager_release_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  wire[25:0] ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  wire ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  wire[2:0] ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  wire[127:0] ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  wire[1:0] ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  wire ManagerTileLinkNetworkPort_io_network_acquire_ready;
  wire ManagerTileLinkNetworkPort_io_network_grant_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id;
  wire[2:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id;
  wire ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type;
  wire[3:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type;
  wire[127:0] ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data;
  wire ManagerTileLinkNetworkPort_io_network_finish_ready;
  wire ManagerTileLinkNetworkPort_io_network_probe_valid;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_src;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst;
  wire[25:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block;
  wire[1:0] ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type;
  wire ManagerTileLinkNetworkPort_io_network_release_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[1:0] LockingRRArbiter_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_io_out_bits_header_dst;
  wire[25:0] LockingRRArbiter_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_payload_addr_beat;
  wire LockingRRArbiter_io_out_bits_payload_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_payload_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_payload_union;
  wire[127:0] LockingRRArbiter_io_out_bits_payload_data;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_addr_beat;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire LockingRRArbiter_1_io_out_bits_payload_voluntary;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire[127:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire RRArbiter_io_in_2_ready;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[1:0] RRArbiter_io_out_bits_header_src;
  wire[1:0] RRArbiter_io_out_bits_header_dst;
  wire[2:0] RRArbiter_io_out_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_acquire_ready;
  wire TileLinkEnqueuer_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_io_client_finish_ready;
  wire TileLinkEnqueuer_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_io_client_release_ready;
  wire TileLinkEnqueuer_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_io_manager_grant_ready;
  wire TileLinkEnqueuer_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_io_manager_probe_ready;
  wire TileLinkEnqueuer_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_acquire_ready;
  wire TileLinkEnqueuer_1_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_1_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_1_io_client_finish_ready;
  wire TileLinkEnqueuer_1_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_1_io_client_release_ready;
  wire TileLinkEnqueuer_1_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_1_io_manager_grant_ready;
  wire TileLinkEnqueuer_1_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_1_io_manager_probe_ready;
  wire TileLinkEnqueuer_1_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_1_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_acquire_ready;
  wire TileLinkEnqueuer_2_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_2_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_2_io_client_finish_ready;
  wire TileLinkEnqueuer_2_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_2_io_client_release_ready;
  wire TileLinkEnqueuer_2_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_2_io_manager_grant_ready;
  wire TileLinkEnqueuer_2_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_2_io_manager_probe_ready;
  wire TileLinkEnqueuer_2_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_2_io_manager_release_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_acquire_ready;
  wire TileLinkEnqueuer_3_io_client_grant_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat;
  wire[1:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id;
  wire[2:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type;
  wire[3:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type;
  wire[127:0] TileLinkEnqueuer_3_io_client_grant_bits_payload_data;
  wire TileLinkEnqueuer_3_io_client_finish_ready;
  wire TileLinkEnqueuer_3_io_client_probe_valid;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type;
  wire TileLinkEnqueuer_3_io_client_release_ready;
  wire TileLinkEnqueuer_3_io_manager_acquire_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst;
  wire[25:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id;
  wire[1:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat;
  wire TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type;
  wire[2:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type;
  wire[16:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union;
  wire[127:0] TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data;
  wire TileLinkEnqueuer_3_io_manager_grant_ready;
  wire TileLinkEnqueuer_3_io_manager_finish_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_finish_bits_header_dst;
  wire[2:0] TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id;
  wire TileLinkEnqueuer_3_io_manager_probe_ready;
  wire TileLinkEnqueuer_3_io_manager_release_valid;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_src;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_header_dst;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat;
  wire[25:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block;
  wire[1:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id;
  wire TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary;
  wire[2:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type;
  wire[127:0] TileLinkEnqueuer_3_io_manager_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_io_client_release_ready;
  wire ClientTileLinkNetworkPort_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  wire ClientTileLinkNetworkPort_2_io_client_grant_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  wire[127:0] ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  wire ClientTileLinkNetworkPort_2_io_client_probe_valid;
  wire[25:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  wire ClientTileLinkNetworkPort_2_io_client_release_ready;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire[16:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire ClientTileLinkNetworkPort_2_io_network_grant_ready;
  wire ClientTileLinkNetworkPort_2_io_network_finish_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_probe_ready;
  wire ClientTileLinkNetworkPort_2_io_network_release_valid;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire[25:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire[1:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire[2:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire[127:0] ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data;


  assign T0 = T5 ? TileLinkEnqueuer_2_io_manager_probe_ready : T1;
  assign T1 = T4 ? TileLinkEnqueuer_1_io_manager_probe_ready : T2;
  assign T2 = T3 ? TileLinkEnqueuer_io_manager_probe_ready : 1'h0;
  assign T3 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h0;
  assign T4 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h1;
  assign T5 = TileLinkEnqueuer_3_io_client_probe_bits_header_dst == 2'h2;
  assign T6 = T11 ? TileLinkEnqueuer_2_io_manager_grant_ready : T7;
  assign T7 = T10 ? TileLinkEnqueuer_1_io_manager_grant_ready : T8;
  assign T8 = T9 ? TileLinkEnqueuer_io_manager_grant_ready : 1'h0;
  assign T9 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h0;
  assign T10 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h1;
  assign T11 = TileLinkEnqueuer_3_io_client_grant_bits_header_dst == 2'h2;
  assign T12 = T5 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T13 = T11 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T14 = T4 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T15 = T10 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign T16 = T3 ? TileLinkEnqueuer_3_io_client_probe_valid : 1'h0;
  assign T17 = T9 ? TileLinkEnqueuer_3_io_client_grant_valid : 1'h0;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_id;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_io_manager_release_bits_data;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_io_manager_release_valid;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_io_manager_probe_ready;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_io_manager_finish_valid;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_io_manager_grant_ready;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_io_manager_acquire_valid;
  assign io_clients_0_release_ready = ClientTileLinkNetworkPort_io_client_release_ready;
  assign io_clients_0_probe_bits_p_type = ClientTileLinkNetworkPort_io_client_probe_bits_p_type;
  assign io_clients_0_probe_bits_addr_block = ClientTileLinkNetworkPort_io_client_probe_bits_addr_block;
  assign io_clients_0_probe_valid = ClientTileLinkNetworkPort_io_client_probe_valid;
  assign io_clients_0_grant_bits_data = ClientTileLinkNetworkPort_io_client_grant_bits_data;
  assign io_clients_0_grant_bits_g_type = ClientTileLinkNetworkPort_io_client_grant_bits_g_type;
  assign io_clients_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type;
  assign io_clients_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id;
  assign io_clients_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id;
  assign io_clients_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat;
  assign io_clients_0_grant_valid = ClientTileLinkNetworkPort_io_client_grant_valid;
  assign io_clients_0_acquire_ready = ClientTileLinkNetworkPort_io_client_acquire_ready;
  assign io_clients_1_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_1_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_1_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_1_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_1_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_1_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_1_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_1_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_1_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_1_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_1_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_1_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_2_release_ready = ClientTileLinkNetworkPort_2_io_client_release_ready;
  assign io_clients_2_probe_bits_p_type = ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type;
  assign io_clients_2_probe_bits_addr_block = ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block;
  assign io_clients_2_probe_valid = ClientTileLinkNetworkPort_2_io_client_probe_valid;
  assign io_clients_2_grant_bits_data = ClientTileLinkNetworkPort_2_io_client_grant_bits_data;
  assign io_clients_2_grant_bits_g_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type;
  assign io_clients_2_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type;
  assign io_clients_2_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id;
  assign io_clients_2_grant_bits_client_xact_id = ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id;
  assign io_clients_2_grant_bits_addr_beat = ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat;
  assign io_clients_2_grant_valid = ClientTileLinkNetworkPort_2_io_client_grant_valid;
  assign io_clients_2_acquire_ready = ClientTileLinkNetworkPort_2_io_client_acquire_ready;
  ClientTileLinkNetworkPort_0 ClientTileLinkNetworkPort(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_0_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_0_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_0_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_0_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_0_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_0_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_0_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_0_acquire_bits_data ),
       .io_client_grant_ready( io_clients_0_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_0_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_io_client_release_ready ),
       .io_client_release_valid( io_clients_0_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_0_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_0_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_0_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_0_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_0_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_0_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_0_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_io_manager_grant_ready ),
       .io_manager_grant_valid( T17 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_0_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_io_manager_probe_ready ),
       .io_manager_probe_valid( T16 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_1 ClientTileLinkNetworkPort_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_1_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_1_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_1_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_1_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_1_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_1_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_1_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_1_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_1_acquire_bits_data ),
       .io_client_grant_ready( io_clients_1_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_1_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_1_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_1_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_1_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_1_io_client_release_ready ),
       .io_client_release_valid( io_clients_1_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_1_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_1_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_1_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_1_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_1_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_1_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_1(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_1_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_1_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_1_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_1_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_1_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_1_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_1_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_1_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_1_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_1_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_1_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_1_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_1_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_1_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_1_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_1_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_1_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_1_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_1_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_1_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_1_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_1_io_manager_grant_ready ),
       .io_manager_grant_valid( T15 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_1_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_1_io_manager_probe_ready ),
       .io_manager_probe_valid( T14 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data )
  );
  ClientTileLinkNetworkPort_2 ClientTileLinkNetworkPort_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( ClientTileLinkNetworkPort_2_io_client_acquire_ready ),
       .io_client_acquire_valid( io_clients_2_acquire_valid ),
       .io_client_acquire_bits_addr_block( io_clients_2_acquire_bits_addr_block ),
       .io_client_acquire_bits_client_xact_id( io_clients_2_acquire_bits_client_xact_id ),
       .io_client_acquire_bits_addr_beat( io_clients_2_acquire_bits_addr_beat ),
       .io_client_acquire_bits_is_builtin_type( io_clients_2_acquire_bits_is_builtin_type ),
       .io_client_acquire_bits_a_type( io_clients_2_acquire_bits_a_type ),
       .io_client_acquire_bits_union( io_clients_2_acquire_bits_union ),
       .io_client_acquire_bits_data( io_clients_2_acquire_bits_data ),
       .io_client_grant_ready( io_clients_2_grant_ready ),
       .io_client_grant_valid( ClientTileLinkNetworkPort_2_io_client_grant_valid ),
       .io_client_grant_bits_addr_beat( ClientTileLinkNetworkPort_2_io_client_grant_bits_addr_beat ),
       .io_client_grant_bits_client_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_client_xact_id ),
       .io_client_grant_bits_manager_xact_id( ClientTileLinkNetworkPort_2_io_client_grant_bits_manager_xact_id ),
       .io_client_grant_bits_is_builtin_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_is_builtin_type ),
       .io_client_grant_bits_g_type( ClientTileLinkNetworkPort_2_io_client_grant_bits_g_type ),
       .io_client_grant_bits_data( ClientTileLinkNetworkPort_2_io_client_grant_bits_data ),
       .io_client_probe_ready( io_clients_2_probe_ready ),
       .io_client_probe_valid( ClientTileLinkNetworkPort_2_io_client_probe_valid ),
       .io_client_probe_bits_addr_block( ClientTileLinkNetworkPort_2_io_client_probe_bits_addr_block ),
       .io_client_probe_bits_p_type( ClientTileLinkNetworkPort_2_io_client_probe_bits_p_type ),
       .io_client_release_ready( ClientTileLinkNetworkPort_2_io_client_release_ready ),
       .io_client_release_valid( io_clients_2_release_valid ),
       .io_client_release_bits_addr_beat( io_clients_2_release_bits_addr_beat ),
       .io_client_release_bits_addr_block( io_clients_2_release_bits_addr_block ),
       .io_client_release_bits_client_xact_id( io_clients_2_release_bits_client_xact_id ),
       .io_client_release_bits_voluntary( io_clients_2_release_bits_voluntary ),
       .io_client_release_bits_r_type( io_clients_2_release_bits_r_type ),
       .io_client_release_bits_data( io_clients_2_release_bits_data ),
       .io_network_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_network_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_network_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_network_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_network_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_network_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_network_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_network_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_network_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_network_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_network_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_network_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_network_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_network_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_network_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data )
  );
  TileLinkEnqueuer_0 TileLinkEnqueuer_2(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_2_io_client_acquire_ready ),
       .io_client_acquire_valid( ClientTileLinkNetworkPort_2_io_network_acquire_valid ),
       .io_client_acquire_bits_header_src( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_src ),
       .io_client_acquire_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_acquire_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_union ),
       .io_client_acquire_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_acquire_bits_payload_data ),
       .io_client_grant_ready( ClientTileLinkNetworkPort_2_io_network_grant_ready ),
       .io_client_grant_valid( TileLinkEnqueuer_2_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_2_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_2_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_2_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_2_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_2_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_2_io_client_finish_ready ),
       .io_client_finish_valid( ClientTileLinkNetworkPort_2_io_network_finish_valid ),
       .io_client_finish_bits_header_src( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_src ),
       .io_client_finish_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_finish_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( ClientTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id ),
       .io_client_probe_ready( ClientTileLinkNetworkPort_2_io_network_probe_ready ),
       .io_client_probe_valid( TileLinkEnqueuer_2_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_2_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_2_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_2_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_2_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_2_io_client_release_ready ),
       .io_client_release_valid( ClientTileLinkNetworkPort_2_io_network_release_valid ),
       .io_client_release_bits_header_src( ClientTileLinkNetworkPort_2_io_network_release_bits_header_src ),
       .io_client_release_bits_header_dst( ClientTileLinkNetworkPort_2_io_network_release_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_r_type ),
       .io_client_release_bits_payload_data( ClientTileLinkNetworkPort_2_io_network_release_bits_payload_data ),
       .io_manager_acquire_ready( LockingRRArbiter_io_in_2_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_2_io_manager_grant_ready ),
       .io_manager_grant_valid( T13 ),
       .io_manager_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_manager_finish_ready( RRArbiter_io_in_2_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_2_io_manager_probe_ready ),
       .io_manager_probe_valid( T12 ),
       .io_manager_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_manager_release_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data )
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort(
       .io_manager_acquire_ready( io_managers_0_acquire_ready ),
       .io_manager_acquire_valid( ManagerTileLinkNetworkPort_io_manager_acquire_valid ),
       .io_manager_acquire_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_block ),
       .io_manager_acquire_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_xact_id ),
       .io_manager_acquire_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_acquire_bits_addr_beat ),
       .io_manager_acquire_bits_is_builtin_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_is_builtin_type ),
       .io_manager_acquire_bits_a_type( ManagerTileLinkNetworkPort_io_manager_acquire_bits_a_type ),
       .io_manager_acquire_bits_union( ManagerTileLinkNetworkPort_io_manager_acquire_bits_union ),
       .io_manager_acquire_bits_data( ManagerTileLinkNetworkPort_io_manager_acquire_bits_data ),
       .io_manager_acquire_bits_client_id( ManagerTileLinkNetworkPort_io_manager_acquire_bits_client_id ),
       .io_manager_grant_ready( ManagerTileLinkNetworkPort_io_manager_grant_ready ),
       .io_manager_grant_valid( io_managers_0_grant_valid ),
       .io_manager_grant_bits_addr_beat( io_managers_0_grant_bits_addr_beat ),
       .io_manager_grant_bits_client_xact_id( io_managers_0_grant_bits_client_xact_id ),
       .io_manager_grant_bits_manager_xact_id( io_managers_0_grant_bits_manager_xact_id ),
       .io_manager_grant_bits_is_builtin_type( io_managers_0_grant_bits_is_builtin_type ),
       .io_manager_grant_bits_g_type( io_managers_0_grant_bits_g_type ),
       .io_manager_grant_bits_data( io_managers_0_grant_bits_data ),
       .io_manager_grant_bits_client_id( io_managers_0_grant_bits_client_id ),
       .io_manager_finish_ready( io_managers_0_finish_ready ),
       .io_manager_finish_valid( ManagerTileLinkNetworkPort_io_manager_finish_valid ),
       .io_manager_finish_bits_manager_xact_id( ManagerTileLinkNetworkPort_io_manager_finish_bits_manager_xact_id ),
       .io_manager_probe_ready( ManagerTileLinkNetworkPort_io_manager_probe_ready ),
       .io_manager_probe_valid( io_managers_0_probe_valid ),
       .io_manager_probe_bits_addr_block( io_managers_0_probe_bits_addr_block ),
       .io_manager_probe_bits_p_type( io_managers_0_probe_bits_p_type ),
       .io_manager_probe_bits_client_id( io_managers_0_probe_bits_client_id ),
       .io_manager_release_ready( io_managers_0_release_ready ),
       .io_manager_release_valid( ManagerTileLinkNetworkPort_io_manager_release_valid ),
       .io_manager_release_bits_addr_beat( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_beat ),
       .io_manager_release_bits_addr_block( ManagerTileLinkNetworkPort_io_manager_release_bits_addr_block ),
       .io_manager_release_bits_client_xact_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_xact_id ),
       .io_manager_release_bits_voluntary( ManagerTileLinkNetworkPort_io_manager_release_bits_voluntary ),
       .io_manager_release_bits_r_type( ManagerTileLinkNetworkPort_io_manager_release_bits_r_type ),
       .io_manager_release_bits_data( ManagerTileLinkNetworkPort_io_manager_release_bits_data ),
       .io_manager_release_bits_client_id( ManagerTileLinkNetworkPort_io_manager_release_bits_client_id ),
       .io_network_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_network_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_network_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_network_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_network_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_network_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_network_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_network_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_network_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_network_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_network_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_network_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_network_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_network_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_network_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_network_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_network_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_network_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_network_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_network_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_network_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_network_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_network_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_network_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_network_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_network_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_network_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_network_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_network_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_network_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_network_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_network_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_network_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_network_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_network_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_network_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_network_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_network_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_network_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_network_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_network_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_network_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_3(.clk(clk), .reset(reset),
       .io_client_acquire_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_client_acquire_valid( LockingRRArbiter_io_out_valid ),
       .io_client_acquire_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_client_acquire_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_client_acquire_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_client_acquire_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_client_acquire_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_client_acquire_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_client_acquire_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_client_acquire_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_client_acquire_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data ),
       .io_client_grant_ready( T6 ),
       .io_client_grant_valid( TileLinkEnqueuer_3_io_client_grant_valid ),
       .io_client_grant_bits_header_src( TileLinkEnqueuer_3_io_client_grant_bits_header_src ),
       .io_client_grant_bits_header_dst( TileLinkEnqueuer_3_io_client_grant_bits_header_dst ),
       .io_client_grant_bits_payload_addr_beat( TileLinkEnqueuer_3_io_client_grant_bits_payload_addr_beat ),
       .io_client_grant_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_client_xact_id ),
       .io_client_grant_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_client_grant_bits_payload_manager_xact_id ),
       .io_client_grant_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_is_builtin_type ),
       .io_client_grant_bits_payload_g_type( TileLinkEnqueuer_3_io_client_grant_bits_payload_g_type ),
       .io_client_grant_bits_payload_data( TileLinkEnqueuer_3_io_client_grant_bits_payload_data ),
       .io_client_finish_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_client_finish_valid( RRArbiter_io_out_valid ),
       .io_client_finish_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_client_finish_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_client_finish_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id ),
       .io_client_probe_ready( T0 ),
       .io_client_probe_valid( TileLinkEnqueuer_3_io_client_probe_valid ),
       .io_client_probe_bits_header_src( TileLinkEnqueuer_3_io_client_probe_bits_header_src ),
       .io_client_probe_bits_header_dst( TileLinkEnqueuer_3_io_client_probe_bits_header_dst ),
       .io_client_probe_bits_payload_addr_block( TileLinkEnqueuer_3_io_client_probe_bits_payload_addr_block ),
       .io_client_probe_bits_payload_p_type( TileLinkEnqueuer_3_io_client_probe_bits_payload_p_type ),
       .io_client_release_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_client_release_valid( LockingRRArbiter_1_io_out_valid ),
       .io_client_release_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_client_release_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_client_release_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_client_release_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_client_release_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_client_release_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_client_release_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_client_release_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_manager_acquire_ready( ManagerTileLinkNetworkPort_io_network_acquire_ready ),
       .io_manager_acquire_valid( TileLinkEnqueuer_3_io_manager_acquire_valid ),
       .io_manager_acquire_bits_header_src( TileLinkEnqueuer_3_io_manager_acquire_bits_header_src ),
       .io_manager_acquire_bits_header_dst( TileLinkEnqueuer_3_io_manager_acquire_bits_header_dst ),
       .io_manager_acquire_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_block ),
       .io_manager_acquire_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_client_xact_id ),
       .io_manager_acquire_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_addr_beat ),
       .io_manager_acquire_bits_payload_is_builtin_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_manager_acquire_bits_payload_a_type( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_a_type ),
       .io_manager_acquire_bits_payload_union( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_union ),
       .io_manager_acquire_bits_payload_data( TileLinkEnqueuer_3_io_manager_acquire_bits_payload_data ),
       .io_manager_grant_ready( TileLinkEnqueuer_3_io_manager_grant_ready ),
       .io_manager_grant_valid( ManagerTileLinkNetworkPort_io_network_grant_valid ),
       .io_manager_grant_bits_header_src( ManagerTileLinkNetworkPort_io_network_grant_bits_header_src ),
       .io_manager_grant_bits_header_dst( ManagerTileLinkNetworkPort_io_network_grant_bits_header_dst ),
       .io_manager_grant_bits_payload_addr_beat( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_addr_beat ),
       .io_manager_grant_bits_payload_client_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_client_xact_id ),
       .io_manager_grant_bits_payload_manager_xact_id( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_manager_xact_id ),
       .io_manager_grant_bits_payload_is_builtin_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_is_builtin_type ),
       .io_manager_grant_bits_payload_g_type( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_g_type ),
       .io_manager_grant_bits_payload_data( ManagerTileLinkNetworkPort_io_network_grant_bits_payload_data ),
       .io_manager_finish_ready( ManagerTileLinkNetworkPort_io_network_finish_ready ),
       .io_manager_finish_valid( TileLinkEnqueuer_3_io_manager_finish_valid ),
       .io_manager_finish_bits_header_src( TileLinkEnqueuer_3_io_manager_finish_bits_header_src ),
       .io_manager_finish_bits_header_dst( TileLinkEnqueuer_3_io_manager_finish_bits_header_dst ),
       .io_manager_finish_bits_payload_manager_xact_id( TileLinkEnqueuer_3_io_manager_finish_bits_payload_manager_xact_id ),
       .io_manager_probe_ready( TileLinkEnqueuer_3_io_manager_probe_ready ),
       .io_manager_probe_valid( ManagerTileLinkNetworkPort_io_network_probe_valid ),
       .io_manager_probe_bits_header_src( ManagerTileLinkNetworkPort_io_network_probe_bits_header_src ),
       .io_manager_probe_bits_header_dst( ManagerTileLinkNetworkPort_io_network_probe_bits_header_dst ),
       .io_manager_probe_bits_payload_addr_block( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_addr_block ),
       .io_manager_probe_bits_payload_p_type( ManagerTileLinkNetworkPort_io_network_probe_bits_payload_p_type ),
       .io_manager_release_ready( ManagerTileLinkNetworkPort_io_network_release_ready ),
       .io_manager_release_valid( TileLinkEnqueuer_3_io_manager_release_valid ),
       .io_manager_release_bits_header_src( TileLinkEnqueuer_3_io_manager_release_bits_header_src ),
       .io_manager_release_bits_header_dst( TileLinkEnqueuer_3_io_manager_release_bits_header_dst ),
       .io_manager_release_bits_payload_addr_beat( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_beat ),
       .io_manager_release_bits_payload_addr_block( TileLinkEnqueuer_3_io_manager_release_bits_payload_addr_block ),
       .io_manager_release_bits_payload_client_xact_id( TileLinkEnqueuer_3_io_manager_release_bits_payload_client_xact_id ),
       .io_manager_release_bits_payload_voluntary( TileLinkEnqueuer_3_io_manager_release_bits_payload_voluntary ),
       .io_manager_release_bits_payload_r_type( TileLinkEnqueuer_3_io_manager_release_bits_payload_r_type ),
       .io_manager_release_bits_payload_data( TileLinkEnqueuer_3_io_manager_release_bits_payload_data )
  );
  LockingRRArbiter_0 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_acquire_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_2_bits_payload_is_builtin_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_2_bits_payload_a_type( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_union( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_union ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_acquire_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_acquire_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_1_bits_payload_is_builtin_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_1_bits_payload_a_type( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_union( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_union ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_acquire_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_acquire_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_acquire_bits_payload_addr_beat ),
       .io_in_0_bits_payload_is_builtin_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_is_builtin_type ),
       .io_in_0_bits_payload_a_type( TileLinkEnqueuer_io_manager_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_union( TileLinkEnqueuer_io_manager_acquire_bits_payload_union ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_acquire_bits_payload_data ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_is_builtin_type( LockingRRArbiter_io_out_bits_payload_is_builtin_type ),
       .io_out_bits_payload_a_type( LockingRRArbiter_io_out_bits_payload_a_type ),
       .io_out_bits_payload_union( LockingRRArbiter_io_out_bits_payload_union ),
       .io_out_bits_payload_data( LockingRRArbiter_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_release_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_release_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_release_bits_header_dst ),
       .io_in_2_bits_payload_addr_beat( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_beat ),
       .io_in_2_bits_payload_addr_block( TileLinkEnqueuer_2_io_manager_release_bits_payload_addr_block ),
       .io_in_2_bits_payload_client_xact_id( TileLinkEnqueuer_2_io_manager_release_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_voluntary( TileLinkEnqueuer_2_io_manager_release_bits_payload_voluntary ),
       .io_in_2_bits_payload_r_type( TileLinkEnqueuer_2_io_manager_release_bits_payload_r_type ),
       .io_in_2_bits_payload_data( TileLinkEnqueuer_2_io_manager_release_bits_payload_data ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_release_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_release_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_release_bits_header_dst ),
       .io_in_1_bits_payload_addr_beat( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_beat ),
       .io_in_1_bits_payload_addr_block( TileLinkEnqueuer_1_io_manager_release_bits_payload_addr_block ),
       .io_in_1_bits_payload_client_xact_id( TileLinkEnqueuer_1_io_manager_release_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_voluntary( TileLinkEnqueuer_1_io_manager_release_bits_payload_voluntary ),
       .io_in_1_bits_payload_r_type( TileLinkEnqueuer_1_io_manager_release_bits_payload_r_type ),
       .io_in_1_bits_payload_data( TileLinkEnqueuer_1_io_manager_release_bits_payload_data ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_release_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_release_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_release_bits_header_dst ),
       .io_in_0_bits_payload_addr_beat( TileLinkEnqueuer_io_manager_release_bits_payload_addr_beat ),
       .io_in_0_bits_payload_addr_block( TileLinkEnqueuer_io_manager_release_bits_payload_addr_block ),
       .io_in_0_bits_payload_client_xact_id( TileLinkEnqueuer_io_manager_release_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_voluntary( TileLinkEnqueuer_io_manager_release_bits_payload_voluntary ),
       .io_in_0_bits_payload_r_type( TileLinkEnqueuer_io_manager_release_bits_payload_r_type ),
       .io_in_0_bits_payload_data( TileLinkEnqueuer_io_manager_release_bits_payload_data ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_release_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr_beat( LockingRRArbiter_1_io_out_bits_payload_addr_beat ),
       .io_out_bits_payload_addr_block( LockingRRArbiter_1_io_out_bits_payload_addr_block ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_voluntary( LockingRRArbiter_1_io_out_bits_payload_voluntary ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data )
       //.io_chosen(  )
  );
  RRArbiter_3 RRArbiter(.clk(clk), .reset(reset),
       .io_in_2_ready( RRArbiter_io_in_2_ready ),
       .io_in_2_valid( TileLinkEnqueuer_2_io_manager_finish_valid ),
       .io_in_2_bits_header_src( TileLinkEnqueuer_2_io_manager_finish_bits_header_src ),
       .io_in_2_bits_header_dst( TileLinkEnqueuer_2_io_manager_finish_bits_header_dst ),
       .io_in_2_bits_payload_manager_xact_id( TileLinkEnqueuer_2_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( TileLinkEnqueuer_1_io_manager_finish_valid ),
       .io_in_1_bits_header_src( TileLinkEnqueuer_1_io_manager_finish_bits_header_src ),
       .io_in_1_bits_header_dst( TileLinkEnqueuer_1_io_manager_finish_bits_header_dst ),
       .io_in_1_bits_payload_manager_xact_id( TileLinkEnqueuer_1_io_manager_finish_bits_payload_manager_xact_id ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( TileLinkEnqueuer_io_manager_finish_valid ),
       .io_in_0_bits_header_src( TileLinkEnqueuer_io_manager_finish_bits_header_src ),
       .io_in_0_bits_header_dst( TileLinkEnqueuer_io_manager_finish_bits_header_dst ),
       .io_in_0_bits_payload_manager_xact_id( TileLinkEnqueuer_io_manager_finish_bits_payload_manager_xact_id ),
       .io_out_ready( TileLinkEnqueuer_3_io_client_finish_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_io_out_bits_header_dst ),
       .io_out_bits_payload_manager_xact_id( RRArbiter_io_out_bits_payload_manager_xact_id )
       //.io_chosen(  )
  );
endmodule

module BroadcastVoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[25:0] io_inner_probe_bits_addr_block
    //output[1:0] io_inner_probe_bits_p_type
    //output[1:0] io_inner_probe_bits_client_id
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T133;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire oacq_data_done;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] R18;
  wire[1:0] T134;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T36;
  wire[3:0] T37;
  wire T38;
  wire T39;
  wire[3:0] T40;
  wire[1:0] T41;
  wire T42;
  reg  collect_irel_data;
  wire T135;
  wire T43;
  wire T44;
  wire T45;
  wire irel_data_done;
  wire T46;
  wire T47;
  wire T48;
  reg [1:0] R49;
  wire[1:0] T136;
  wire[1:0] T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire[3:0] T65;
  wire[1:0] T66;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T67;
  wire[3:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[1:0] T74;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T75;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T76;
  wire[3:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire[16:0] T90;
  wire[16:0] T91;
  wire[15:0] T92;
  wire[2:0] T93;
  wire T94;
  wire[1:0] T95;
  wire[2:0] T137;
  wire[1:0] T96;
  wire[25:0] T97;
  reg [25:0] xact_addr_block;
  wire[25:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire T106;
  reg [3:0] irel_data_valid;
  wire[3:0] T138;
  wire[3:0] T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T139;
  wire T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[1:0] T123;
  reg [1:0] xact_client_id;
  wire[1:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire T127;
  wire[2:0] T128;
  wire[1:0] T129;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T130;
  wire[1:0] T131;
  wire T132;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    R18 = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    collect_irel_data = {1{$random}};
    R49 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_addr_block = {1{$random}};
    irel_data_valid = {1{$random}};
    xact_client_id = {1{$random}};
    xact_client_xact_id = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_inner_probe_bits_client_id = {1{$random}};
//  assign io_inner_probe_bits_p_type = {1{$random}};
//  assign io_inner_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign io_has_release_match = io_inner_release_bits_voluntary;
  assign io_has_acquire_match = 1'h0;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = T0;
  assign T0 = T1 ? io_inner_grant_ready : 1'h0;
  assign T1 = 2'h2 == state;
  assign T133 = reset ? 2'h0 : T2;
  assign T2 = T31 ? 2'h0 : T3;
  assign T3 = T29 ? T25 : T4;
  assign T4 = T14 ? 2'h2 : T5;
  assign T5 = T12 ? T6 : state;
  assign T6 = T7 ? 2'h1 : 2'h3;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_inner_release_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_inner_release_bits_r_type;
  assign T11 = 3'h0 == io_inner_release_bits_r_type;
  assign T12 = T13 & io_inner_release_valid;
  assign T13 = 2'h0 == state;
  assign T14 = T24 & oacq_data_done;
  assign oacq_data_done = T22 ? T16 : T15;
  assign T15 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T16 = T21 & T17;
  assign T17 = R18 == 2'h3;
  assign T134 = reset ? 2'h0 : T19;
  assign T19 = T21 ? T20 : R18;
  assign T20 = R18 + 2'h1;
  assign T21 = T15 & T22;
  assign T22 = io_outer_acquire_bits_is_builtin_type & T23;
  assign T23 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T24 = 2'h1 == state;
  assign T25 = T26 ? 2'h3 : 2'h0;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_inner_grant_bits_is_builtin_type & T28;
  assign T28 = io_inner_grant_bits_g_type == 4'h0;
  assign T29 = T1 & T30;
  assign T30 = io_inner_grant_ready & io_inner_grant_valid;
  assign T31 = T32 & io_inner_finish_valid;
  assign T32 = 2'h3 == state;
  assign io_outer_acquire_bits_data = T33;
  assign T33 = T34;
  assign T34 = T89 ? T75 : T35;
  assign T35 = T73 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T36 = T63 ? io_inner_release_bits_data : T37;
  assign T37 = T38 ? io_inner_release_bits_data : xact_data_buffer_0;
  assign T38 = T42 & T39;
  assign T39 = T40[1'h0:1'h0];
  assign T40 = 1'h1 << T41;
  assign T41 = io_inner_release_bits_addr_beat;
  assign T42 = collect_irel_data & io_inner_release_valid;
  assign T135 = reset ? 1'h0 : T43;
  assign T43 = T12 ? T58 : T44;
  assign T44 = T45 ? 1'h0 : collect_irel_data;
  assign T45 = collect_irel_data & irel_data_done;
  assign irel_data_done = T53 ? T47 : T46;
  assign T46 = io_inner_release_ready & io_inner_release_valid;
  assign T47 = T52 & T48;
  assign T48 = R49 == 2'h3;
  assign T136 = reset ? 2'h0 : T50;
  assign T50 = T52 ? T51 : R49;
  assign T51 = R49 + 2'h1;
  assign T52 = T46 & T53;
  assign T53 = T55 | T54;
  assign T54 = 3'h2 == io_inner_release_bits_r_type;
  assign T55 = T57 | T56;
  assign T56 = 3'h1 == io_inner_release_bits_r_type;
  assign T57 = 3'h0 == io_inner_release_bits_r_type;
  assign T58 = T60 | T59;
  assign T59 = 3'h2 == io_inner_release_bits_r_type;
  assign T60 = T62 | T61;
  assign T61 = 3'h1 == io_inner_release_bits_r_type;
  assign T62 = 3'h0 == io_inner_release_bits_r_type;
  assign T63 = T12 & T64;
  assign T64 = T65[1'h0:1'h0];
  assign T65 = 1'h1 << T66;
  assign T66 = 2'h0;
  assign T67 = T71 ? io_inner_release_bits_data : T68;
  assign T68 = T69 ? io_inner_release_bits_data : xact_data_buffer_1;
  assign T69 = T42 & T70;
  assign T70 = T40[1'h1:1'h1];
  assign T71 = T12 & T72;
  assign T72 = T65[1'h1:1'h1];
  assign T73 = T74[1'h0:1'h0];
  assign T74 = oacq_data_cnt;
  assign oacq_data_cnt = T22 ? R18 : 2'h0;
  assign T75 = T88 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T76 = T80 ? io_inner_release_bits_data : T77;
  assign T77 = T78 ? io_inner_release_bits_data : xact_data_buffer_2;
  assign T78 = T42 & T79;
  assign T79 = T40[2'h2:2'h2];
  assign T80 = T12 & T81;
  assign T81 = T65[2'h2:2'h2];
  assign T82 = T86 ? io_inner_release_bits_data : T83;
  assign T83 = T84 ? io_inner_release_bits_data : xact_data_buffer_3;
  assign T84 = T42 & T85;
  assign T85 = T40[2'h3:2'h3];
  assign T86 = T12 & T87;
  assign T87 = T65[2'h3:2'h3];
  assign T88 = T74[1'h0:1'h0];
  assign T89 = T74[1'h1:1'h1];
  assign io_outer_acquire_bits_union = T90;
  assign T90 = T91;
  assign T91 = {T92, 1'h1};
  assign T92 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T93;
  assign T93 = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T94;
  assign T94 = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T95;
  assign T95 = oacq_data_cnt;
  assign io_outer_acquire_bits_client_xact_id = T137;
  assign T137 = {1'h0, T96};
  assign T96 = 2'h0;
  assign io_outer_acquire_bits_addr_block = T97;
  assign T97 = xact_addr_block;
  assign T98 = T12 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign io_outer_acquire_valid = T99;
  assign T99 = T24 ? T100 : 1'h0;
  assign T100 = T121 | T101;
  assign T101 = T106 & T102;
  assign T102 = T103 - 1'h1;
  assign T103 = 1'h1 << T104;
  assign T104 = T105 + 2'h1;
  assign T105 = oacq_data_cnt - oacq_data_cnt;
  assign T106 = irel_data_valid >> oacq_data_cnt;
  assign T138 = reset ? 4'h0 : T107;
  assign T107 = T12 ? T115 : T108;
  assign T108 = T42 ? T109 : irel_data_valid;
  assign T109 = T113 | T110;
  assign T110 = T139 & T111;
  assign T111 = 1'h1 << io_inner_release_bits_addr_beat;
  assign T139 = T112 ? 4'hf : 4'h0;
  assign T112 = 1'h1;
  assign T113 = irel_data_valid & T114;
  assign T114 = ~ T111;
  assign T115 = T116 << io_inner_release_bits_addr_beat;
  assign T116 = T118 | T117;
  assign T117 = 3'h2 == io_inner_release_bits_r_type;
  assign T118 = T120 | T119;
  assign T119 = 3'h1 == io_inner_release_bits_r_type;
  assign T120 = 3'h0 == io_inner_release_bits_r_type;
  assign T121 = collect_irel_data ^ 1'h1;
  assign io_inner_release_ready = T122;
  assign T122 = T13 ? 1'h1 : collect_irel_data;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_finish_ready = T32;
  assign io_inner_grant_bits_client_id = T123;
  assign T123 = xact_client_id;
  assign T124 = T12 ? io_inner_release_bits_client_id : xact_client_id;
  assign io_inner_grant_bits_data = T125;
  assign T125 = 4'h0;
  assign io_inner_grant_bits_g_type = T126;
  assign T126 = 4'h0;
  assign io_inner_grant_bits_is_builtin_type = T127;
  assign T127 = 1'h1;
  assign io_inner_grant_bits_manager_xact_id = T128;
  assign T128 = 3'h0;
  assign io_inner_grant_bits_client_xact_id = T129;
  assign T129 = xact_client_xact_id;
  assign T130 = T12 ? io_inner_release_bits_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T131;
  assign T131 = 2'h0;
  assign io_inner_grant_valid = T132;
  assign T132 = T1 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T31) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= T25;
    end else if(T14) begin
      state <= 2'h2;
    end else if(T12) begin
      state <= T6;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T21) begin
      R18 <= T20;
    end
    if(T63) begin
      xact_data_buffer_0 <= io_inner_release_bits_data;
    end else if(T38) begin
      xact_data_buffer_0 <= io_inner_release_bits_data;
    end
    if(reset) begin
      collect_irel_data <= 1'h0;
    end else if(T12) begin
      collect_irel_data <= T58;
    end else if(T45) begin
      collect_irel_data <= 1'h0;
    end
    if(reset) begin
      R49 <= 2'h0;
    end else if(T52) begin
      R49 <= T51;
    end
    if(T71) begin
      xact_data_buffer_1 <= io_inner_release_bits_data;
    end else if(T69) begin
      xact_data_buffer_1 <= io_inner_release_bits_data;
    end
    if(T80) begin
      xact_data_buffer_2 <= io_inner_release_bits_data;
    end else if(T78) begin
      xact_data_buffer_2 <= io_inner_release_bits_data;
    end
    if(T86) begin
      xact_data_buffer_3 <= io_inner_release_bits_data;
    end else if(T84) begin
      xact_data_buffer_3 <= io_inner_release_bits_data;
    end
    if(T12) begin
      xact_addr_block <= io_inner_release_bits_addr_block;
    end
    if(reset) begin
      irel_data_valid <= 4'h0;
    end else if(T12) begin
      irel_data_valid <= T115;
    end else if(T42) begin
      irel_data_valid <= T109;
    end
    if(T12) begin
      xact_client_id <= io_inner_release_bits_client_id;
    end
    if(T12) begin
      xact_client_xact_id <= io_inner_release_bits_client_xact_id;
    end
  end
endmodule

module BroadcastAcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T482;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T483;
  wire[2:0] T25;
  wire[2:0] T484;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T485;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T486;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T487;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T488;
  wire[2:0] T489;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T490;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T491;
  wire T88;
  wire[2:0] T492;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T493;
  wire T92;
  wire T93;
  wire[2:0] T494;
  wire T94;
  wire[2:0] T495;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire oacq_data_done;
  wire T106;
  wire T107;
  wire T108;
  reg [1:0] R109;
  wire[1:0] T496;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  wire[2:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[2:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire ignt_data_done;
  wire T132;
  wire T133;
  wire T134;
  reg [1:0] R135;
  wire[1:0] T497;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  reg  collect_iacq_data;
  wire T498;
  wire T162;
  wire T163;
  wire T164;
  wire iacq_data_done;
  wire T165;
  wire T166;
  wire T167;
  reg [1:0] R168;
  wire[1:0] T499;
  wire[1:0] T169;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg[0:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg [1:0] xact_client_id;
  wire[1:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  reg [25:0] xact_addr_block;
  wire[25:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg  pending_ognt_ack;
  wire T500;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[3:0] T224;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T225;
  wire[3:0] T226;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T227;
  wire[3:0] T228;
  wire T229;
  wire T230;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire[3:0] T236;
  wire[1:0] T237;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T238;
  wire[3:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire[1:0] T245;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T246;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T247;
  wire[3:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T253;
  wire[3:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[3:0] oacq_write_beat_data;
  wire T261;
  wire[3:0] oacq_probe_data;
  wire T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] T265;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T501;
  wire[12:0] T266;
  wire[6:0] T267;
  wire[2:0] T268;
  reg [16:0] xact_union;
  wire[16:0] T269;
  wire[3:0] T270;
  wire[16:0] T271;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire[15:0] T285;
  wire[15:0] T286;
  wire[7:0] T287;
  wire[7:0] T502;
  wire T288;
  wire[1:0] T289;
  wire T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T503;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[3:0] T298;
  wire[1:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire[15:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[15:0] T308;
  wire[15:0] T309;
  wire[7:0] T310;
  wire[7:0] T504;
  wire T311;
  wire[1:0] T312;
  wire T313;
  wire[3:0] T314;
  wire[7:0] T315;
  wire[7:0] T505;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[1:0] T322;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T323;
  wire[15:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[1:0] T330;
  wire[15:0] T331;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T332;
  wire[15:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T338;
  wire[15:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[15:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire[15:0] T355;
  wire[15:0] T356;
  wire[7:0] T357;
  wire[7:0] T506;
  wire T358;
  wire[1:0] T359;
  wire T360;
  wire[3:0] T361;
  wire[7:0] T362;
  wire[7:0] T507;
  wire T363;
  wire T364;
  wire T365;
  wire[16:0] oacq_probe_union;
  wire[16:0] T366;
  wire[15:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] T370;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T371;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T372;
  wire T373;
  wire T374;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T375;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] oacq_read_block_client_xact_id;
  wire[2:0] oacq_read_beat_client_xact_id;
  wire[2:0] T384;
  wire[2:0] oacq_write_block_client_xact_id;
  wire[2:0] oacq_write_beat_client_xact_id;
  wire[2:0] oacq_probe_client_xact_id;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] T387;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T388;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  reg [3:0] iacq_data_valid;
  wire[3:0] T508;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[3:0] T509;
  wire T404;
  wire[3:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T510;
  wire[1:0] T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire T436;
  wire T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[25:0] T452;
  wire T453;
  wire T454;
  reg  pending_probes;
  wire T511;
  wire[3:0] T512;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[1:0] T428;
  wire T429;
  wire T430;
  wire[1:0] T515;
  wire T431;
  wire[1:0] T455;
  wire[3:0] T456;
  wire[3:0] T457;
  wire[3:0] T516;
  wire[2:0] T458;
  wire[2:0] T517;
  wire[1:0] T459;
  wire T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[2:0] T476;
  wire[1:0] T477;
  wire[1:0] T478;
  wire T479;
  wire T480;
  wire T481;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R109 = {1{$random}};
    R135 = {1{$random}};
    T153 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R168 = {1{$random}};
    T177 = 1'b0;
    xact_client_id = {1{$random}};
    T187 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T482 = reset ? 3'h0 : T11;
  assign T11 = T151 ? 3'h0 : T12;
  assign T12 = T149 ? T145 : T13;
  assign T13 = T131 ? T127 : T14;
  assign T14 = T124 ? 3'h5 : T15;
  assign T15 = T122 ? T121 : T16;
  assign T16 = T119 ? T117 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T483;
  assign T483 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T484;
  assign T484 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T485;
  assign T485 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T486 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T486 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T487 & T59;
  assign T59 = ~ T56;
  assign T487 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T105 & T79;
  assign T79 = release_count == 1'h1;
  assign T488 = T489[1'h0:1'h0];
  assign T489 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T495 : T81;
  assign T81 = T105 ? T494 : T82;
  assign T82 = T93 ? T83 : T490;
  assign T490 = {2'h0, release_count};
  assign T83 = T492 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T491 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3:2'h3];
  assign T491 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2:2'h2];
  assign T492 = {1'h0, T89};
  assign T89 = T493 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1:1'h1];
  assign T493 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0:1'h0];
  assign T93 = T61 & T52;
  assign T494 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T495 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T104 & io_inner_release_valid;
  assign T104 = 3'h1 == state;
  assign T105 = T115 & oacq_data_done;
  assign oacq_data_done = T113 ? T107 : T106;
  assign T106 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T107 = T112 & T108;
  assign T108 = R109 == 2'h3;
  assign T496 = reset ? 2'h0 : T110;
  assign T110 = T112 ? T111 : R109;
  assign T111 = R109 + 2'h1;
  assign T112 = T106 & T113;
  assign T113 = io_outer_acquire_bits_is_builtin_type & T114;
  assign T114 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T115 = T116 & io_outer_acquire_ready;
  assign T116 = T103 & T98;
  assign T117 = pending_outer_write ? 3'h3 : T118;
  assign T118 = pending_outer_read ? 3'h2 : 3'h4;
  assign T119 = T96 & T120;
  assign T120 = release_count == 1'h1;
  assign T121 = pending_outer_read ? 3'h2 : 3'h5;
  assign T122 = T123 & oacq_data_done;
  assign T123 = 3'h3 == state;
  assign T124 = T126 & T125;
  assign T125 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T126 = 3'h2 == state;
  assign T127 = T128 ? 3'h6 : 3'h0;
  assign T128 = T129 ^ 1'h1;
  assign T129 = io_inner_grant_bits_is_builtin_type & T130;
  assign T130 = io_inner_grant_bits_g_type == 4'h0;
  assign T131 = T144 & ignt_data_done;
  assign ignt_data_done = T139 ? T133 : T132;
  assign T132 = io_inner_grant_ready & io_inner_grant_valid;
  assign T133 = T138 & T134;
  assign T134 = R135 == 2'h3;
  assign T497 = reset ? 2'h0 : T136;
  assign T136 = T138 ? T137 : R135;
  assign T137 = R135 + 2'h1;
  assign T138 = T132 & T139;
  assign T139 = io_inner_grant_bits_is_builtin_type ? T143 : T140;
  assign T140 = T142 | T141;
  assign T141 = 4'h1 == io_inner_grant_bits_g_type;
  assign T142 = 4'h0 == io_inner_grant_bits_g_type;
  assign T143 = 4'h5 == io_inner_grant_bits_g_type;
  assign T144 = 3'h5 == state;
  assign T145 = T146 ? 3'h6 : 3'h0;
  assign T146 = T147 ^ 1'h1;
  assign T147 = io_inner_grant_bits_is_builtin_type & T148;
  assign T148 = io_inner_grant_bits_g_type == 4'h0;
  assign T149 = T150 & io_inner_grant_ready;
  assign T150 = 3'h4 == state;
  assign T151 = T152 & io_inner_finish_valid;
  assign T152 = 3'h6 == state;
  assign T154 = T155 | reset;
  assign T155 = T156 ^ 1'h1;
  assign T156 = T159 & T157;
  assign T157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T158 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T159 = T161 & T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T176 & collect_iacq_data;
  assign T498 = reset ? 1'h0 : T162;
  assign T162 = T61 ? T174 : T163;
  assign T163 = T164 ? 1'h0 : collect_iacq_data;
  assign T164 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T172 ? T166 : T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T171 & T167;
  assign T167 = R168 == 2'h3;
  assign T499 = reset ? 2'h0 : T169;
  assign T169 = T171 ? T170 : R168;
  assign T170 = R168 + 2'h1;
  assign T171 = T165 & T172;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = io_inner_acquire_bits_is_builtin_type & T175;
  assign T175 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T176 = state != 3'h0;
  assign T178 = T179 | reset;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T183 & T181;
  assign T181 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T182 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T183 = T185 & T184;
  assign T184 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T185 = T186 & collect_iacq_data;
  assign T186 = state != 3'h0;
  assign T188 = T189 | reset;
  assign T189 = T190 ^ 1'h1;
  assign T190 = T196 & T191;
  assign T191 = T193 | T192;
  assign T192 = 3'h6 == xact_a_type;
  assign T193 = T195 | T194;
  assign T194 = 3'h5 == xact_a_type;
  assign T195 = 3'h4 == xact_a_type;
  assign T196 = T197 & xact_is_builtin_type;
  assign T197 = state != 3'h0;
  assign io_has_release_match = T198;
  assign T198 = T200 & T199;
  assign T199 = state == 3'h1;
  assign T200 = T202 & T201;
  assign T201 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T202 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T203 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T204;
  assign T204 = T205 & collect_iacq_data;
  assign T205 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T206;
  assign T206 = T208 & T207;
  assign T207 = collect_iacq_data ^ 1'h1;
  assign T208 = T210 & T209;
  assign T209 = state != 3'h0;
  assign T210 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T211;
  assign T211 = T144 ? io_inner_grant_ready : pending_ognt_ack;
  assign T500 = reset ? 1'h0 : T212;
  assign T212 = T122 ? 1'h1 : T213;
  assign T213 = T105 ? 1'h1 : T214;
  assign T214 = T215 ? 1'h0 : pending_ognt_ack;
  assign T215 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T216;
  assign T216 = T262 ? oacq_probe_data : T217;
  assign T217 = T261 ? T224 : T218;
  assign T218 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T219;
  assign T219 = T221 | T220;
  assign T220 = 3'h4 == xact_a_type;
  assign T221 = T223 | T222;
  assign T222 = 3'h0 == xact_a_type;
  assign T223 = 3'h2 == xact_a_type;
  assign T224 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T225;
  assign T225 = T260 ? T246 : T226;
  assign T226 = T244 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T227 = T234 ? io_inner_acquire_bits_data : T228;
  assign T228 = T229 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T229 = T233 & T230;
  assign T230 = T231[1'h0:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = io_inner_acquire_bits_addr_beat;
  assign T233 = collect_iacq_data & io_inner_acquire_valid;
  assign T234 = T61 & T235;
  assign T235 = T236[1'h0:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = 2'h0;
  assign T238 = T242 ? io_inner_acquire_bits_data : T239;
  assign T239 = T240 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T240 = T233 & T241;
  assign T241 = T231[1'h1:1'h1];
  assign T242 = T61 & T243;
  assign T243 = T236[1'h1:1'h1];
  assign T244 = T245[1'h0:1'h0];
  assign T245 = oacq_data_cnt;
  assign oacq_data_cnt = T113 ? R109 : 2'h0;
  assign T246 = T259 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T247 = T251 ? io_inner_acquire_bits_data : T248;
  assign T248 = T249 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T249 = T233 & T250;
  assign T250 = T231[2'h2:2'h2];
  assign T251 = T61 & T252;
  assign T252 = T236[2'h2:2'h2];
  assign T253 = T257 ? io_inner_acquire_bits_data : T254;
  assign T254 = T255 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T255 = T233 & T256;
  assign T256 = T231[2'h3:2'h3];
  assign T257 = T61 & T258;
  assign T258 = T236[2'h3:2'h3];
  assign T259 = T245[1'h0:1'h0];
  assign T260 = T245[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T261 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T262 = state == 3'h1;
  assign io_outer_acquire_bits_union = T263;
  assign T263 = T262 ? oacq_probe_union : T264;
  assign T264 = T261 ? T271 : T265;
  assign T265 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T501;
  assign T501 = {4'h0, T266};
  assign T266 = {T267, 6'h0};
  assign T267 = {T270, T268};
  assign T268 = xact_union[4'h8:3'h6];
  assign T269 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T270 = xact_union[4'hc:4'h9];
  assign T271 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T272;
  assign T272 = {T273, 1'h1};
  assign T273 = T345 ? T331 : T274;
  assign T274 = T329 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T275 = T319 ? T300 : T276;
  assign T276 = T296 ? T277 : xact_wmask_buffer_0;
  assign T277 = T294 ? T285 : T278;
  assign T278 = T280 ? T279 : 16'h0;
  assign T279 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T280 = T283 | T281;
  assign T281 = io_inner_acquire_bits_is_builtin_type & T282;
  assign T282 = io_inner_acquire_bits_a_type == 3'h2;
  assign T283 = io_inner_acquire_bits_is_builtin_type & T284;
  assign T284 = io_inner_acquire_bits_a_type == 3'h3;
  assign T285 = T286;
  assign T286 = {T292, T287};
  assign T287 = 8'h0 - T502;
  assign T502 = {7'h0, T288};
  assign T288 = T289[1'h0:1'h0];
  assign T289 = 1'h1 << T290;
  assign T290 = T291[2'h3:2'h3];
  assign T291 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T292 = 8'h0 - T503;
  assign T503 = {7'h0, T293};
  assign T293 = T289[1'h1:1'h1];
  assign T294 = io_inner_acquire_bits_is_builtin_type & T295;
  assign T295 = io_inner_acquire_bits_a_type == 3'h4;
  assign T296 = T233 & T297;
  assign T297 = T298[1'h0:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = io_inner_acquire_bits_addr_beat;
  assign T300 = T317 ? T308 : T301;
  assign T301 = T303 ? T302 : 16'h0;
  assign T302 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T303 = T306 | T304;
  assign T304 = io_inner_acquire_bits_is_builtin_type & T305;
  assign T305 = io_inner_acquire_bits_a_type == 3'h2;
  assign T306 = io_inner_acquire_bits_is_builtin_type & T307;
  assign T307 = io_inner_acquire_bits_a_type == 3'h3;
  assign T308 = T309;
  assign T309 = {T315, T310};
  assign T310 = 8'h0 - T504;
  assign T504 = {7'h0, T311};
  assign T311 = T312[1'h0:1'h0];
  assign T312 = 1'h1 << T313;
  assign T313 = T314[2'h3:2'h3];
  assign T314 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T315 = 8'h0 - T505;
  assign T505 = {7'h0, T316};
  assign T316 = T312[1'h1:1'h1];
  assign T317 = io_inner_acquire_bits_is_builtin_type & T318;
  assign T318 = io_inner_acquire_bits_a_type == 3'h4;
  assign T319 = T61 & T320;
  assign T320 = T321[1'h0:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = 2'h0;
  assign T323 = T327 ? T300 : T324;
  assign T324 = T325 ? T277 : xact_wmask_buffer_1;
  assign T325 = T233 & T326;
  assign T326 = T298[1'h1:1'h1];
  assign T327 = T61 & T328;
  assign T328 = T321[1'h1:1'h1];
  assign T329 = T330[1'h0:1'h0];
  assign T330 = oacq_data_cnt;
  assign T331 = T344 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T332 = T336 ? T300 : T333;
  assign T333 = T334 ? T277 : xact_wmask_buffer_2;
  assign T334 = T233 & T335;
  assign T335 = T298[2'h2:2'h2];
  assign T336 = T61 & T337;
  assign T337 = T321[2'h2:2'h2];
  assign T338 = T342 ? T300 : T339;
  assign T339 = T340 ? T277 : xact_wmask_buffer_3;
  assign T340 = T233 & T341;
  assign T341 = T298[2'h3:2'h3];
  assign T342 = T61 & T343;
  assign T343 = T321[2'h3:2'h3];
  assign T344 = T330[1'h0:1'h0];
  assign T345 = T330[1'h1:1'h1];
  assign oacq_write_beat_union = T346;
  assign T346 = {T347, 1'h1};
  assign T347 = T364 ? T355 : T348;
  assign T348 = T350 ? T349 : 16'h0;
  assign T349 = xact_union[5'h10:1'h1];
  assign T350 = T353 | T351;
  assign T351 = xact_is_builtin_type & T352;
  assign T352 = xact_a_type == 3'h2;
  assign T353 = xact_is_builtin_type & T354;
  assign T354 = xact_a_type == 3'h3;
  assign T355 = T356;
  assign T356 = {T362, T357};
  assign T357 = 8'h0 - T506;
  assign T506 = {7'h0, T358};
  assign T358 = T359[1'h0:1'h0];
  assign T359 = 1'h1 << T360;
  assign T360 = T361[2'h3:2'h3];
  assign T361 = xact_union[4'hc:4'h9];
  assign T362 = 8'h0 - T507;
  assign T507 = {7'h0, T363};
  assign T363 = T359[1'h1:1'h1];
  assign T364 = xact_is_builtin_type & T365;
  assign T365 = xact_a_type == 3'h4;
  assign oacq_probe_union = T366;
  assign T366 = {T367, 1'h1};
  assign T367 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T368;
  assign T368 = T262 ? oacq_probe_a_type : T369;
  assign T369 = T261 ? T371 : T370;
  assign T370 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T371 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T372;
  assign T372 = T262 ? oacq_probe_is_builtin_type : T373;
  assign T373 = T261 ? T375 : T374;
  assign T374 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T375 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T376;
  assign T376 = T262 ? oacq_probe_addr_beat : T377;
  assign T377 = T261 ? T380 : T378;
  assign T378 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T379 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T380 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T381;
  assign T381 = T262 ? oacq_probe_client_xact_id : T382;
  assign T382 = T261 ? T384 : T383;
  assign T383 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 3'h1;
  assign oacq_read_beat_client_xact_id = 3'h1;
  assign T384 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 3'h1;
  assign oacq_write_beat_client_xact_id = 3'h1;
  assign oacq_probe_client_xact_id = 3'h1;
  assign io_outer_acquire_bits_addr_block = T385;
  assign T385 = T262 ? oacq_probe_addr_block : T386;
  assign T386 = T261 ? T388 : T387;
  assign T387 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T388 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T389;
  assign T389 = T126 ? T416 : T390;
  assign T390 = T123 ? T391 : T116;
  assign T391 = T415 & T392;
  assign T392 = T414 | T393;
  assign T393 = T398 & T394;
  assign T394 = T395 - 1'h1;
  assign T395 = 1'h1 << T396;
  assign T396 = T397 + 2'h1;
  assign T397 = oacq_data_cnt - oacq_data_cnt;
  assign T398 = iacq_data_valid >> oacq_data_cnt;
  assign T508 = reset ? 4'h0 : T399;
  assign T399 = T61 ? T407 : T400;
  assign T400 = T233 ? T401 : iacq_data_valid;
  assign T401 = T405 | T402;
  assign T402 = T509 & T403;
  assign T403 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T509 = T404 ? 4'hf : 4'h0;
  assign T404 = 1'h1;
  assign T405 = iacq_data_valid & T406;
  assign T406 = ~ T403;
  assign T407 = T408 << io_inner_acquire_bits_addr_beat;
  assign T408 = io_inner_acquire_bits_is_builtin_type & T409;
  assign T409 = T411 | T410;
  assign T410 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T411 = T413 | T412;
  assign T412 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T413 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T414 = collect_iacq_data ^ 1'h1;
  assign T415 = pending_ognt_ack ^ 1'h1;
  assign T416 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T417;
  assign T417 = T104 ? T418 : 1'h0;
  assign T418 = T419 | io_outer_acquire_ready;
  assign T419 = T420 ^ 1'h1;
  assign T420 = T422 | T421;
  assign T421 = 3'h2 == io_inner_release_bits_r_type;
  assign T422 = T424 | T423;
  assign T423 = 3'h1 == io_inner_release_bits_r_type;
  assign T424 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T425;
  assign T425 = T510;
  assign T510 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T432;
  assign T432 = T433;
  assign T433 = xact_is_builtin_type ? T438 : T434;
  assign T434 = T437 ? 2'h1 : T435;
  assign T435 = T436 ? 2'h0 : 2'h2;
  assign T436 = xact_a_type == 3'h1;
  assign T437 = xact_a_type == 3'h0;
  assign T438 = T451 ? 2'h2 : T439;
  assign T439 = T450 ? 2'h0 : T440;
  assign T440 = T449 ? 2'h2 : T441;
  assign T441 = T448 ? 2'h0 : T442;
  assign T442 = T447 ? 2'h2 : T443;
  assign T443 = T446 ? 2'h0 : T444;
  assign T444 = T445 ? 2'h0 : 2'h2;
  assign T445 = xact_a_type == 3'h4;
  assign T446 = xact_a_type == 3'h6;
  assign T447 = xact_a_type == 3'h5;
  assign T448 = xact_a_type == 3'h2;
  assign T449 = xact_a_type == 3'h0;
  assign T450 = xact_a_type == 3'h3;
  assign T451 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T452;
  assign T452 = xact_addr_block;
  assign io_inner_probe_valid = T453;
  assign T453 = T104 ? T454 : 1'h0;
  assign T454 = pending_probes != 1'h0;
  assign T511 = T512[1'h0:1'h0];
  assign T512 = reset ? 4'h0 : T426;
  assign T426 = T431 ? T514 : T427;
  assign T427 = T93 ? mask_incoherent : T513;
  assign T513 = {3'h0, pending_probes};
  assign T514 = {2'h0, T428};
  assign T428 = T515 & T429;
  assign T429 = ~ T430;
  assign T430 = 1'h1 << 1'h0;
  assign T515 = {1'h0, pending_probes};
  assign T431 = T104 & io_inner_probe_ready;
  assign io_inner_finish_ready = T152;
  assign io_inner_grant_bits_client_id = T455;
  assign T455 = xact_client_id;
  assign io_inner_grant_bits_data = T456;
  assign T456 = 4'h0;
  assign io_inner_grant_bits_g_type = T457;
  assign T457 = T516;
  assign T516 = {1'h0, T458};
  assign T458 = xact_is_builtin_type ? T461 : T517;
  assign T517 = {1'h0, T459};
  assign T459 = T460 ? 2'h0 : 2'h1;
  assign T460 = xact_a_type == 3'h0;
  assign T461 = T474 ? 3'h4 : T462;
  assign T462 = T473 ? 3'h5 : T463;
  assign T463 = T472 ? 3'h3 : T464;
  assign T464 = T471 ? 3'h3 : T465;
  assign T465 = T470 ? 3'h4 : T466;
  assign T466 = T469 ? 3'h1 : T467;
  assign T467 = T468 ? 3'h1 : 3'h3;
  assign T468 = xact_a_type == 3'h6;
  assign T469 = xact_a_type == 3'h5;
  assign T470 = xact_a_type == 3'h4;
  assign T471 = xact_a_type == 3'h3;
  assign T472 = xact_a_type == 3'h2;
  assign T473 = xact_a_type == 3'h1;
  assign T474 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T475;
  assign T475 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T476;
  assign T476 = 3'h1;
  assign io_inner_grant_bits_client_xact_id = T477;
  assign T477 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T478;
  assign T478 = 2'h0;
  assign io_inner_grant_valid = T479;
  assign T479 = T150 ? 1'h1 : T480;
  assign T480 = T144 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T481;
  assign T481 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T187 <= 1'b1;
  if(!T188 && T187 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T177 <= 1'b1;
  if(!T178 && T177 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T153 <= 1'b1;
  if(!T154 && T153 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T151) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= T145;
    end else if(T131) begin
      state <= T127;
    end else if(T124) begin
      state <= 3'h5;
    end else if(T122) begin
      state <= T121;
    end else if(T119) begin
      state <= T117;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T488;
    if(reset) begin
      R109 <= 2'h0;
    end else if(T112) begin
      R109 <= T111;
    end
    if(reset) begin
      R135 <= 2'h0;
    end else if(T138) begin
      R135 <= T137;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T174;
    end else if(T164) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R168 <= 2'h0;
    end else if(T171) begin
      R168 <= T170;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T122) begin
      pending_ognt_ack <= 1'h1;
    end else if(T105) begin
      pending_ognt_ack <= 1'h1;
    end else if(T215) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T234) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T229) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T242) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T240) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T251) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T249) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T257) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T255) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T319) begin
      xact_wmask_buffer_0 <= T300;
    end else if(T296) begin
      xact_wmask_buffer_0 <= T277;
    end
    if(T327) begin
      xact_wmask_buffer_1 <= T300;
    end else if(T325) begin
      xact_wmask_buffer_1 <= T277;
    end
    if(T336) begin
      xact_wmask_buffer_2 <= T300;
    end else if(T334) begin
      xact_wmask_buffer_2 <= T277;
    end
    if(T342) begin
      xact_wmask_buffer_3 <= T300;
    end else if(T340) begin
      xact_wmask_buffer_3 <= T277;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T407;
    end else if(T233) begin
      iacq_data_valid <= T401;
    end
    pending_probes <= T511;
  end
endmodule

module BroadcastAcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T482;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T483;
  wire[2:0] T25;
  wire[2:0] T484;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T485;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T486;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T487;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T488;
  wire[2:0] T489;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T490;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T491;
  wire T88;
  wire[2:0] T492;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T493;
  wire T92;
  wire T93;
  wire[2:0] T494;
  wire T94;
  wire[2:0] T495;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire oacq_data_done;
  wire T106;
  wire T107;
  wire T108;
  reg [1:0] R109;
  wire[1:0] T496;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  wire[2:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[2:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire ignt_data_done;
  wire T132;
  wire T133;
  wire T134;
  reg [1:0] R135;
  wire[1:0] T497;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  reg  collect_iacq_data;
  wire T498;
  wire T162;
  wire T163;
  wire T164;
  wire iacq_data_done;
  wire T165;
  wire T166;
  wire T167;
  reg [1:0] R168;
  wire[1:0] T499;
  wire[1:0] T169;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg[0:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg [1:0] xact_client_id;
  wire[1:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  reg [25:0] xact_addr_block;
  wire[25:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg  pending_ognt_ack;
  wire T500;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[3:0] T224;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T225;
  wire[3:0] T226;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T227;
  wire[3:0] T228;
  wire T229;
  wire T230;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire[3:0] T236;
  wire[1:0] T237;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T238;
  wire[3:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire[1:0] T245;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T246;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T247;
  wire[3:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T253;
  wire[3:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[3:0] oacq_write_beat_data;
  wire T261;
  wire[3:0] oacq_probe_data;
  wire T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] T265;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T501;
  wire[12:0] T266;
  wire[6:0] T267;
  wire[2:0] T268;
  reg [16:0] xact_union;
  wire[16:0] T269;
  wire[3:0] T270;
  wire[16:0] T271;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire[15:0] T285;
  wire[15:0] T286;
  wire[7:0] T287;
  wire[7:0] T502;
  wire T288;
  wire[1:0] T289;
  wire T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T503;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[3:0] T298;
  wire[1:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire[15:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[15:0] T308;
  wire[15:0] T309;
  wire[7:0] T310;
  wire[7:0] T504;
  wire T311;
  wire[1:0] T312;
  wire T313;
  wire[3:0] T314;
  wire[7:0] T315;
  wire[7:0] T505;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[1:0] T322;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T323;
  wire[15:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[1:0] T330;
  wire[15:0] T331;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T332;
  wire[15:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T338;
  wire[15:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[15:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire[15:0] T355;
  wire[15:0] T356;
  wire[7:0] T357;
  wire[7:0] T506;
  wire T358;
  wire[1:0] T359;
  wire T360;
  wire[3:0] T361;
  wire[7:0] T362;
  wire[7:0] T507;
  wire T363;
  wire T364;
  wire T365;
  wire[16:0] oacq_probe_union;
  wire[16:0] T366;
  wire[15:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] T370;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T371;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T372;
  wire T373;
  wire T374;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T375;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] oacq_read_block_client_xact_id;
  wire[2:0] oacq_read_beat_client_xact_id;
  wire[2:0] T384;
  wire[2:0] oacq_write_block_client_xact_id;
  wire[2:0] oacq_write_beat_client_xact_id;
  wire[2:0] oacq_probe_client_xact_id;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] T387;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T388;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  reg [3:0] iacq_data_valid;
  wire[3:0] T508;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[3:0] T509;
  wire T404;
  wire[3:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T510;
  wire[1:0] T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire T436;
  wire T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[25:0] T452;
  wire T453;
  wire T454;
  reg  pending_probes;
  wire T511;
  wire[3:0] T512;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[1:0] T428;
  wire T429;
  wire T430;
  wire[1:0] T515;
  wire T431;
  wire[1:0] T455;
  wire[3:0] T456;
  wire[3:0] T457;
  wire[3:0] T516;
  wire[2:0] T458;
  wire[2:0] T517;
  wire[1:0] T459;
  wire T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[2:0] T476;
  wire[1:0] T477;
  wire[1:0] T478;
  wire T479;
  wire T480;
  wire T481;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R109 = {1{$random}};
    R135 = {1{$random}};
    T153 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R168 = {1{$random}};
    T177 = 1'b0;
    xact_client_id = {1{$random}};
    T187 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T482 = reset ? 3'h0 : T11;
  assign T11 = T151 ? 3'h0 : T12;
  assign T12 = T149 ? T145 : T13;
  assign T13 = T131 ? T127 : T14;
  assign T14 = T124 ? 3'h5 : T15;
  assign T15 = T122 ? T121 : T16;
  assign T16 = T119 ? T117 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T483;
  assign T483 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T484;
  assign T484 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T485;
  assign T485 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T486 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T486 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T487 & T59;
  assign T59 = ~ T56;
  assign T487 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T105 & T79;
  assign T79 = release_count == 1'h1;
  assign T488 = T489[1'h0:1'h0];
  assign T489 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T495 : T81;
  assign T81 = T105 ? T494 : T82;
  assign T82 = T93 ? T83 : T490;
  assign T490 = {2'h0, release_count};
  assign T83 = T492 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T491 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3:2'h3];
  assign T491 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2:2'h2];
  assign T492 = {1'h0, T89};
  assign T89 = T493 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1:1'h1];
  assign T493 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0:1'h0];
  assign T93 = T61 & T52;
  assign T494 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T495 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T104 & io_inner_release_valid;
  assign T104 = 3'h1 == state;
  assign T105 = T115 & oacq_data_done;
  assign oacq_data_done = T113 ? T107 : T106;
  assign T106 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T107 = T112 & T108;
  assign T108 = R109 == 2'h3;
  assign T496 = reset ? 2'h0 : T110;
  assign T110 = T112 ? T111 : R109;
  assign T111 = R109 + 2'h1;
  assign T112 = T106 & T113;
  assign T113 = io_outer_acquire_bits_is_builtin_type & T114;
  assign T114 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T115 = T116 & io_outer_acquire_ready;
  assign T116 = T103 & T98;
  assign T117 = pending_outer_write ? 3'h3 : T118;
  assign T118 = pending_outer_read ? 3'h2 : 3'h4;
  assign T119 = T96 & T120;
  assign T120 = release_count == 1'h1;
  assign T121 = pending_outer_read ? 3'h2 : 3'h5;
  assign T122 = T123 & oacq_data_done;
  assign T123 = 3'h3 == state;
  assign T124 = T126 & T125;
  assign T125 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T126 = 3'h2 == state;
  assign T127 = T128 ? 3'h6 : 3'h0;
  assign T128 = T129 ^ 1'h1;
  assign T129 = io_inner_grant_bits_is_builtin_type & T130;
  assign T130 = io_inner_grant_bits_g_type == 4'h0;
  assign T131 = T144 & ignt_data_done;
  assign ignt_data_done = T139 ? T133 : T132;
  assign T132 = io_inner_grant_ready & io_inner_grant_valid;
  assign T133 = T138 & T134;
  assign T134 = R135 == 2'h3;
  assign T497 = reset ? 2'h0 : T136;
  assign T136 = T138 ? T137 : R135;
  assign T137 = R135 + 2'h1;
  assign T138 = T132 & T139;
  assign T139 = io_inner_grant_bits_is_builtin_type ? T143 : T140;
  assign T140 = T142 | T141;
  assign T141 = 4'h1 == io_inner_grant_bits_g_type;
  assign T142 = 4'h0 == io_inner_grant_bits_g_type;
  assign T143 = 4'h5 == io_inner_grant_bits_g_type;
  assign T144 = 3'h5 == state;
  assign T145 = T146 ? 3'h6 : 3'h0;
  assign T146 = T147 ^ 1'h1;
  assign T147 = io_inner_grant_bits_is_builtin_type & T148;
  assign T148 = io_inner_grant_bits_g_type == 4'h0;
  assign T149 = T150 & io_inner_grant_ready;
  assign T150 = 3'h4 == state;
  assign T151 = T152 & io_inner_finish_valid;
  assign T152 = 3'h6 == state;
  assign T154 = T155 | reset;
  assign T155 = T156 ^ 1'h1;
  assign T156 = T159 & T157;
  assign T157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T158 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T159 = T161 & T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T176 & collect_iacq_data;
  assign T498 = reset ? 1'h0 : T162;
  assign T162 = T61 ? T174 : T163;
  assign T163 = T164 ? 1'h0 : collect_iacq_data;
  assign T164 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T172 ? T166 : T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T171 & T167;
  assign T167 = R168 == 2'h3;
  assign T499 = reset ? 2'h0 : T169;
  assign T169 = T171 ? T170 : R168;
  assign T170 = R168 + 2'h1;
  assign T171 = T165 & T172;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = io_inner_acquire_bits_is_builtin_type & T175;
  assign T175 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T176 = state != 3'h0;
  assign T178 = T179 | reset;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T183 & T181;
  assign T181 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T182 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T183 = T185 & T184;
  assign T184 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T185 = T186 & collect_iacq_data;
  assign T186 = state != 3'h0;
  assign T188 = T189 | reset;
  assign T189 = T190 ^ 1'h1;
  assign T190 = T196 & T191;
  assign T191 = T193 | T192;
  assign T192 = 3'h6 == xact_a_type;
  assign T193 = T195 | T194;
  assign T194 = 3'h5 == xact_a_type;
  assign T195 = 3'h4 == xact_a_type;
  assign T196 = T197 & xact_is_builtin_type;
  assign T197 = state != 3'h0;
  assign io_has_release_match = T198;
  assign T198 = T200 & T199;
  assign T199 = state == 3'h1;
  assign T200 = T202 & T201;
  assign T201 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T202 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T203 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T204;
  assign T204 = T205 & collect_iacq_data;
  assign T205 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T206;
  assign T206 = T208 & T207;
  assign T207 = collect_iacq_data ^ 1'h1;
  assign T208 = T210 & T209;
  assign T209 = state != 3'h0;
  assign T210 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T211;
  assign T211 = T144 ? io_inner_grant_ready : pending_ognt_ack;
  assign T500 = reset ? 1'h0 : T212;
  assign T212 = T122 ? 1'h1 : T213;
  assign T213 = T105 ? 1'h1 : T214;
  assign T214 = T215 ? 1'h0 : pending_ognt_ack;
  assign T215 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T216;
  assign T216 = T262 ? oacq_probe_data : T217;
  assign T217 = T261 ? T224 : T218;
  assign T218 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T219;
  assign T219 = T221 | T220;
  assign T220 = 3'h4 == xact_a_type;
  assign T221 = T223 | T222;
  assign T222 = 3'h0 == xact_a_type;
  assign T223 = 3'h2 == xact_a_type;
  assign T224 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T225;
  assign T225 = T260 ? T246 : T226;
  assign T226 = T244 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T227 = T234 ? io_inner_acquire_bits_data : T228;
  assign T228 = T229 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T229 = T233 & T230;
  assign T230 = T231[1'h0:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = io_inner_acquire_bits_addr_beat;
  assign T233 = collect_iacq_data & io_inner_acquire_valid;
  assign T234 = T61 & T235;
  assign T235 = T236[1'h0:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = 2'h0;
  assign T238 = T242 ? io_inner_acquire_bits_data : T239;
  assign T239 = T240 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T240 = T233 & T241;
  assign T241 = T231[1'h1:1'h1];
  assign T242 = T61 & T243;
  assign T243 = T236[1'h1:1'h1];
  assign T244 = T245[1'h0:1'h0];
  assign T245 = oacq_data_cnt;
  assign oacq_data_cnt = T113 ? R109 : 2'h0;
  assign T246 = T259 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T247 = T251 ? io_inner_acquire_bits_data : T248;
  assign T248 = T249 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T249 = T233 & T250;
  assign T250 = T231[2'h2:2'h2];
  assign T251 = T61 & T252;
  assign T252 = T236[2'h2:2'h2];
  assign T253 = T257 ? io_inner_acquire_bits_data : T254;
  assign T254 = T255 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T255 = T233 & T256;
  assign T256 = T231[2'h3:2'h3];
  assign T257 = T61 & T258;
  assign T258 = T236[2'h3:2'h3];
  assign T259 = T245[1'h0:1'h0];
  assign T260 = T245[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T261 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T262 = state == 3'h1;
  assign io_outer_acquire_bits_union = T263;
  assign T263 = T262 ? oacq_probe_union : T264;
  assign T264 = T261 ? T271 : T265;
  assign T265 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T501;
  assign T501 = {4'h0, T266};
  assign T266 = {T267, 6'h0};
  assign T267 = {T270, T268};
  assign T268 = xact_union[4'h8:3'h6];
  assign T269 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T270 = xact_union[4'hc:4'h9];
  assign T271 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T272;
  assign T272 = {T273, 1'h1};
  assign T273 = T345 ? T331 : T274;
  assign T274 = T329 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T275 = T319 ? T300 : T276;
  assign T276 = T296 ? T277 : xact_wmask_buffer_0;
  assign T277 = T294 ? T285 : T278;
  assign T278 = T280 ? T279 : 16'h0;
  assign T279 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T280 = T283 | T281;
  assign T281 = io_inner_acquire_bits_is_builtin_type & T282;
  assign T282 = io_inner_acquire_bits_a_type == 3'h2;
  assign T283 = io_inner_acquire_bits_is_builtin_type & T284;
  assign T284 = io_inner_acquire_bits_a_type == 3'h3;
  assign T285 = T286;
  assign T286 = {T292, T287};
  assign T287 = 8'h0 - T502;
  assign T502 = {7'h0, T288};
  assign T288 = T289[1'h0:1'h0];
  assign T289 = 1'h1 << T290;
  assign T290 = T291[2'h3:2'h3];
  assign T291 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T292 = 8'h0 - T503;
  assign T503 = {7'h0, T293};
  assign T293 = T289[1'h1:1'h1];
  assign T294 = io_inner_acquire_bits_is_builtin_type & T295;
  assign T295 = io_inner_acquire_bits_a_type == 3'h4;
  assign T296 = T233 & T297;
  assign T297 = T298[1'h0:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = io_inner_acquire_bits_addr_beat;
  assign T300 = T317 ? T308 : T301;
  assign T301 = T303 ? T302 : 16'h0;
  assign T302 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T303 = T306 | T304;
  assign T304 = io_inner_acquire_bits_is_builtin_type & T305;
  assign T305 = io_inner_acquire_bits_a_type == 3'h2;
  assign T306 = io_inner_acquire_bits_is_builtin_type & T307;
  assign T307 = io_inner_acquire_bits_a_type == 3'h3;
  assign T308 = T309;
  assign T309 = {T315, T310};
  assign T310 = 8'h0 - T504;
  assign T504 = {7'h0, T311};
  assign T311 = T312[1'h0:1'h0];
  assign T312 = 1'h1 << T313;
  assign T313 = T314[2'h3:2'h3];
  assign T314 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T315 = 8'h0 - T505;
  assign T505 = {7'h0, T316};
  assign T316 = T312[1'h1:1'h1];
  assign T317 = io_inner_acquire_bits_is_builtin_type & T318;
  assign T318 = io_inner_acquire_bits_a_type == 3'h4;
  assign T319 = T61 & T320;
  assign T320 = T321[1'h0:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = 2'h0;
  assign T323 = T327 ? T300 : T324;
  assign T324 = T325 ? T277 : xact_wmask_buffer_1;
  assign T325 = T233 & T326;
  assign T326 = T298[1'h1:1'h1];
  assign T327 = T61 & T328;
  assign T328 = T321[1'h1:1'h1];
  assign T329 = T330[1'h0:1'h0];
  assign T330 = oacq_data_cnt;
  assign T331 = T344 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T332 = T336 ? T300 : T333;
  assign T333 = T334 ? T277 : xact_wmask_buffer_2;
  assign T334 = T233 & T335;
  assign T335 = T298[2'h2:2'h2];
  assign T336 = T61 & T337;
  assign T337 = T321[2'h2:2'h2];
  assign T338 = T342 ? T300 : T339;
  assign T339 = T340 ? T277 : xact_wmask_buffer_3;
  assign T340 = T233 & T341;
  assign T341 = T298[2'h3:2'h3];
  assign T342 = T61 & T343;
  assign T343 = T321[2'h3:2'h3];
  assign T344 = T330[1'h0:1'h0];
  assign T345 = T330[1'h1:1'h1];
  assign oacq_write_beat_union = T346;
  assign T346 = {T347, 1'h1};
  assign T347 = T364 ? T355 : T348;
  assign T348 = T350 ? T349 : 16'h0;
  assign T349 = xact_union[5'h10:1'h1];
  assign T350 = T353 | T351;
  assign T351 = xact_is_builtin_type & T352;
  assign T352 = xact_a_type == 3'h2;
  assign T353 = xact_is_builtin_type & T354;
  assign T354 = xact_a_type == 3'h3;
  assign T355 = T356;
  assign T356 = {T362, T357};
  assign T357 = 8'h0 - T506;
  assign T506 = {7'h0, T358};
  assign T358 = T359[1'h0:1'h0];
  assign T359 = 1'h1 << T360;
  assign T360 = T361[2'h3:2'h3];
  assign T361 = xact_union[4'hc:4'h9];
  assign T362 = 8'h0 - T507;
  assign T507 = {7'h0, T363};
  assign T363 = T359[1'h1:1'h1];
  assign T364 = xact_is_builtin_type & T365;
  assign T365 = xact_a_type == 3'h4;
  assign oacq_probe_union = T366;
  assign T366 = {T367, 1'h1};
  assign T367 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T368;
  assign T368 = T262 ? oacq_probe_a_type : T369;
  assign T369 = T261 ? T371 : T370;
  assign T370 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T371 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T372;
  assign T372 = T262 ? oacq_probe_is_builtin_type : T373;
  assign T373 = T261 ? T375 : T374;
  assign T374 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T375 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T376;
  assign T376 = T262 ? oacq_probe_addr_beat : T377;
  assign T377 = T261 ? T380 : T378;
  assign T378 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T379 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T380 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T381;
  assign T381 = T262 ? oacq_probe_client_xact_id : T382;
  assign T382 = T261 ? T384 : T383;
  assign T383 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 3'h2;
  assign oacq_read_beat_client_xact_id = 3'h2;
  assign T384 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 3'h2;
  assign oacq_write_beat_client_xact_id = 3'h2;
  assign oacq_probe_client_xact_id = 3'h2;
  assign io_outer_acquire_bits_addr_block = T385;
  assign T385 = T262 ? oacq_probe_addr_block : T386;
  assign T386 = T261 ? T388 : T387;
  assign T387 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T388 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T389;
  assign T389 = T126 ? T416 : T390;
  assign T390 = T123 ? T391 : T116;
  assign T391 = T415 & T392;
  assign T392 = T414 | T393;
  assign T393 = T398 & T394;
  assign T394 = T395 - 1'h1;
  assign T395 = 1'h1 << T396;
  assign T396 = T397 + 2'h1;
  assign T397 = oacq_data_cnt - oacq_data_cnt;
  assign T398 = iacq_data_valid >> oacq_data_cnt;
  assign T508 = reset ? 4'h0 : T399;
  assign T399 = T61 ? T407 : T400;
  assign T400 = T233 ? T401 : iacq_data_valid;
  assign T401 = T405 | T402;
  assign T402 = T509 & T403;
  assign T403 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T509 = T404 ? 4'hf : 4'h0;
  assign T404 = 1'h1;
  assign T405 = iacq_data_valid & T406;
  assign T406 = ~ T403;
  assign T407 = T408 << io_inner_acquire_bits_addr_beat;
  assign T408 = io_inner_acquire_bits_is_builtin_type & T409;
  assign T409 = T411 | T410;
  assign T410 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T411 = T413 | T412;
  assign T412 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T413 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T414 = collect_iacq_data ^ 1'h1;
  assign T415 = pending_ognt_ack ^ 1'h1;
  assign T416 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T417;
  assign T417 = T104 ? T418 : 1'h0;
  assign T418 = T419 | io_outer_acquire_ready;
  assign T419 = T420 ^ 1'h1;
  assign T420 = T422 | T421;
  assign T421 = 3'h2 == io_inner_release_bits_r_type;
  assign T422 = T424 | T423;
  assign T423 = 3'h1 == io_inner_release_bits_r_type;
  assign T424 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T425;
  assign T425 = T510;
  assign T510 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T432;
  assign T432 = T433;
  assign T433 = xact_is_builtin_type ? T438 : T434;
  assign T434 = T437 ? 2'h1 : T435;
  assign T435 = T436 ? 2'h0 : 2'h2;
  assign T436 = xact_a_type == 3'h1;
  assign T437 = xact_a_type == 3'h0;
  assign T438 = T451 ? 2'h2 : T439;
  assign T439 = T450 ? 2'h0 : T440;
  assign T440 = T449 ? 2'h2 : T441;
  assign T441 = T448 ? 2'h0 : T442;
  assign T442 = T447 ? 2'h2 : T443;
  assign T443 = T446 ? 2'h0 : T444;
  assign T444 = T445 ? 2'h0 : 2'h2;
  assign T445 = xact_a_type == 3'h4;
  assign T446 = xact_a_type == 3'h6;
  assign T447 = xact_a_type == 3'h5;
  assign T448 = xact_a_type == 3'h2;
  assign T449 = xact_a_type == 3'h0;
  assign T450 = xact_a_type == 3'h3;
  assign T451 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T452;
  assign T452 = xact_addr_block;
  assign io_inner_probe_valid = T453;
  assign T453 = T104 ? T454 : 1'h0;
  assign T454 = pending_probes != 1'h0;
  assign T511 = T512[1'h0:1'h0];
  assign T512 = reset ? 4'h0 : T426;
  assign T426 = T431 ? T514 : T427;
  assign T427 = T93 ? mask_incoherent : T513;
  assign T513 = {3'h0, pending_probes};
  assign T514 = {2'h0, T428};
  assign T428 = T515 & T429;
  assign T429 = ~ T430;
  assign T430 = 1'h1 << 1'h0;
  assign T515 = {1'h0, pending_probes};
  assign T431 = T104 & io_inner_probe_ready;
  assign io_inner_finish_ready = T152;
  assign io_inner_grant_bits_client_id = T455;
  assign T455 = xact_client_id;
  assign io_inner_grant_bits_data = T456;
  assign T456 = 4'h0;
  assign io_inner_grant_bits_g_type = T457;
  assign T457 = T516;
  assign T516 = {1'h0, T458};
  assign T458 = xact_is_builtin_type ? T461 : T517;
  assign T517 = {1'h0, T459};
  assign T459 = T460 ? 2'h0 : 2'h1;
  assign T460 = xact_a_type == 3'h0;
  assign T461 = T474 ? 3'h4 : T462;
  assign T462 = T473 ? 3'h5 : T463;
  assign T463 = T472 ? 3'h3 : T464;
  assign T464 = T471 ? 3'h3 : T465;
  assign T465 = T470 ? 3'h4 : T466;
  assign T466 = T469 ? 3'h1 : T467;
  assign T467 = T468 ? 3'h1 : 3'h3;
  assign T468 = xact_a_type == 3'h6;
  assign T469 = xact_a_type == 3'h5;
  assign T470 = xact_a_type == 3'h4;
  assign T471 = xact_a_type == 3'h3;
  assign T472 = xact_a_type == 3'h2;
  assign T473 = xact_a_type == 3'h1;
  assign T474 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T475;
  assign T475 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T476;
  assign T476 = 3'h2;
  assign io_inner_grant_bits_client_xact_id = T477;
  assign T477 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T478;
  assign T478 = 2'h0;
  assign io_inner_grant_valid = T479;
  assign T479 = T150 ? 1'h1 : T480;
  assign T480 = T144 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T481;
  assign T481 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T187 <= 1'b1;
  if(!T188 && T187 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T177 <= 1'b1;
  if(!T178 && T177 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T153 <= 1'b1;
  if(!T154 && T153 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T151) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= T145;
    end else if(T131) begin
      state <= T127;
    end else if(T124) begin
      state <= 3'h5;
    end else if(T122) begin
      state <= T121;
    end else if(T119) begin
      state <= T117;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T488;
    if(reset) begin
      R109 <= 2'h0;
    end else if(T112) begin
      R109 <= T111;
    end
    if(reset) begin
      R135 <= 2'h0;
    end else if(T138) begin
      R135 <= T137;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T174;
    end else if(T164) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R168 <= 2'h0;
    end else if(T171) begin
      R168 <= T170;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T122) begin
      pending_ognt_ack <= 1'h1;
    end else if(T105) begin
      pending_ognt_ack <= 1'h1;
    end else if(T215) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T234) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T229) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T242) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T240) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T251) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T249) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T257) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T255) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T319) begin
      xact_wmask_buffer_0 <= T300;
    end else if(T296) begin
      xact_wmask_buffer_0 <= T277;
    end
    if(T327) begin
      xact_wmask_buffer_1 <= T300;
    end else if(T325) begin
      xact_wmask_buffer_1 <= T277;
    end
    if(T336) begin
      xact_wmask_buffer_2 <= T300;
    end else if(T334) begin
      xact_wmask_buffer_2 <= T277;
    end
    if(T342) begin
      xact_wmask_buffer_3 <= T300;
    end else if(T340) begin
      xact_wmask_buffer_3 <= T277;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T407;
    end else if(T233) begin
      iacq_data_valid <= T401;
    end
    pending_probes <= T511;
  end
endmodule

module BroadcastAcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T482;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T483;
  wire[2:0] T25;
  wire[2:0] T484;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T485;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T486;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T487;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T488;
  wire[2:0] T489;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T490;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T491;
  wire T88;
  wire[2:0] T492;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T493;
  wire T92;
  wire T93;
  wire[2:0] T494;
  wire T94;
  wire[2:0] T495;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire oacq_data_done;
  wire T106;
  wire T107;
  wire T108;
  reg [1:0] R109;
  wire[1:0] T496;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  wire[2:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[2:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire ignt_data_done;
  wire T132;
  wire T133;
  wire T134;
  reg [1:0] R135;
  wire[1:0] T497;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  reg  collect_iacq_data;
  wire T498;
  wire T162;
  wire T163;
  wire T164;
  wire iacq_data_done;
  wire T165;
  wire T166;
  wire T167;
  reg [1:0] R168;
  wire[1:0] T499;
  wire[1:0] T169;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg[0:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg [1:0] xact_client_id;
  wire[1:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  reg [25:0] xact_addr_block;
  wire[25:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg  pending_ognt_ack;
  wire T500;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[3:0] T224;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T225;
  wire[3:0] T226;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T227;
  wire[3:0] T228;
  wire T229;
  wire T230;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire[3:0] T236;
  wire[1:0] T237;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T238;
  wire[3:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire[1:0] T245;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T246;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T247;
  wire[3:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T253;
  wire[3:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[3:0] oacq_write_beat_data;
  wire T261;
  wire[3:0] oacq_probe_data;
  wire T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] T265;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T501;
  wire[12:0] T266;
  wire[6:0] T267;
  wire[2:0] T268;
  reg [16:0] xact_union;
  wire[16:0] T269;
  wire[3:0] T270;
  wire[16:0] T271;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire[15:0] T285;
  wire[15:0] T286;
  wire[7:0] T287;
  wire[7:0] T502;
  wire T288;
  wire[1:0] T289;
  wire T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T503;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[3:0] T298;
  wire[1:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire[15:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[15:0] T308;
  wire[15:0] T309;
  wire[7:0] T310;
  wire[7:0] T504;
  wire T311;
  wire[1:0] T312;
  wire T313;
  wire[3:0] T314;
  wire[7:0] T315;
  wire[7:0] T505;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[1:0] T322;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T323;
  wire[15:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[1:0] T330;
  wire[15:0] T331;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T332;
  wire[15:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T338;
  wire[15:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[15:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire[15:0] T355;
  wire[15:0] T356;
  wire[7:0] T357;
  wire[7:0] T506;
  wire T358;
  wire[1:0] T359;
  wire T360;
  wire[3:0] T361;
  wire[7:0] T362;
  wire[7:0] T507;
  wire T363;
  wire T364;
  wire T365;
  wire[16:0] oacq_probe_union;
  wire[16:0] T366;
  wire[15:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] T370;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T371;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T372;
  wire T373;
  wire T374;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T375;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] oacq_read_block_client_xact_id;
  wire[2:0] oacq_read_beat_client_xact_id;
  wire[2:0] T384;
  wire[2:0] oacq_write_block_client_xact_id;
  wire[2:0] oacq_write_beat_client_xact_id;
  wire[2:0] oacq_probe_client_xact_id;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] T387;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T388;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  reg [3:0] iacq_data_valid;
  wire[3:0] T508;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[3:0] T509;
  wire T404;
  wire[3:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T510;
  wire[1:0] T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire T436;
  wire T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[25:0] T452;
  wire T453;
  wire T454;
  reg  pending_probes;
  wire T511;
  wire[3:0] T512;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[1:0] T428;
  wire T429;
  wire T430;
  wire[1:0] T515;
  wire T431;
  wire[1:0] T455;
  wire[3:0] T456;
  wire[3:0] T457;
  wire[3:0] T516;
  wire[2:0] T458;
  wire[2:0] T517;
  wire[1:0] T459;
  wire T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[2:0] T476;
  wire[1:0] T477;
  wire[1:0] T478;
  wire T479;
  wire T480;
  wire T481;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R109 = {1{$random}};
    R135 = {1{$random}};
    T153 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R168 = {1{$random}};
    T177 = 1'b0;
    xact_client_id = {1{$random}};
    T187 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T482 = reset ? 3'h0 : T11;
  assign T11 = T151 ? 3'h0 : T12;
  assign T12 = T149 ? T145 : T13;
  assign T13 = T131 ? T127 : T14;
  assign T14 = T124 ? 3'h5 : T15;
  assign T15 = T122 ? T121 : T16;
  assign T16 = T119 ? T117 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T483;
  assign T483 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T484;
  assign T484 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T485;
  assign T485 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T486 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T486 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T487 & T59;
  assign T59 = ~ T56;
  assign T487 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T105 & T79;
  assign T79 = release_count == 1'h1;
  assign T488 = T489[1'h0:1'h0];
  assign T489 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T495 : T81;
  assign T81 = T105 ? T494 : T82;
  assign T82 = T93 ? T83 : T490;
  assign T490 = {2'h0, release_count};
  assign T83 = T492 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T491 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3:2'h3];
  assign T491 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2:2'h2];
  assign T492 = {1'h0, T89};
  assign T89 = T493 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1:1'h1];
  assign T493 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0:1'h0];
  assign T93 = T61 & T52;
  assign T494 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T495 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T104 & io_inner_release_valid;
  assign T104 = 3'h1 == state;
  assign T105 = T115 & oacq_data_done;
  assign oacq_data_done = T113 ? T107 : T106;
  assign T106 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T107 = T112 & T108;
  assign T108 = R109 == 2'h3;
  assign T496 = reset ? 2'h0 : T110;
  assign T110 = T112 ? T111 : R109;
  assign T111 = R109 + 2'h1;
  assign T112 = T106 & T113;
  assign T113 = io_outer_acquire_bits_is_builtin_type & T114;
  assign T114 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T115 = T116 & io_outer_acquire_ready;
  assign T116 = T103 & T98;
  assign T117 = pending_outer_write ? 3'h3 : T118;
  assign T118 = pending_outer_read ? 3'h2 : 3'h4;
  assign T119 = T96 & T120;
  assign T120 = release_count == 1'h1;
  assign T121 = pending_outer_read ? 3'h2 : 3'h5;
  assign T122 = T123 & oacq_data_done;
  assign T123 = 3'h3 == state;
  assign T124 = T126 & T125;
  assign T125 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T126 = 3'h2 == state;
  assign T127 = T128 ? 3'h6 : 3'h0;
  assign T128 = T129 ^ 1'h1;
  assign T129 = io_inner_grant_bits_is_builtin_type & T130;
  assign T130 = io_inner_grant_bits_g_type == 4'h0;
  assign T131 = T144 & ignt_data_done;
  assign ignt_data_done = T139 ? T133 : T132;
  assign T132 = io_inner_grant_ready & io_inner_grant_valid;
  assign T133 = T138 & T134;
  assign T134 = R135 == 2'h3;
  assign T497 = reset ? 2'h0 : T136;
  assign T136 = T138 ? T137 : R135;
  assign T137 = R135 + 2'h1;
  assign T138 = T132 & T139;
  assign T139 = io_inner_grant_bits_is_builtin_type ? T143 : T140;
  assign T140 = T142 | T141;
  assign T141 = 4'h1 == io_inner_grant_bits_g_type;
  assign T142 = 4'h0 == io_inner_grant_bits_g_type;
  assign T143 = 4'h5 == io_inner_grant_bits_g_type;
  assign T144 = 3'h5 == state;
  assign T145 = T146 ? 3'h6 : 3'h0;
  assign T146 = T147 ^ 1'h1;
  assign T147 = io_inner_grant_bits_is_builtin_type & T148;
  assign T148 = io_inner_grant_bits_g_type == 4'h0;
  assign T149 = T150 & io_inner_grant_ready;
  assign T150 = 3'h4 == state;
  assign T151 = T152 & io_inner_finish_valid;
  assign T152 = 3'h6 == state;
  assign T154 = T155 | reset;
  assign T155 = T156 ^ 1'h1;
  assign T156 = T159 & T157;
  assign T157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T158 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T159 = T161 & T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T176 & collect_iacq_data;
  assign T498 = reset ? 1'h0 : T162;
  assign T162 = T61 ? T174 : T163;
  assign T163 = T164 ? 1'h0 : collect_iacq_data;
  assign T164 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T172 ? T166 : T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T171 & T167;
  assign T167 = R168 == 2'h3;
  assign T499 = reset ? 2'h0 : T169;
  assign T169 = T171 ? T170 : R168;
  assign T170 = R168 + 2'h1;
  assign T171 = T165 & T172;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = io_inner_acquire_bits_is_builtin_type & T175;
  assign T175 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T176 = state != 3'h0;
  assign T178 = T179 | reset;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T183 & T181;
  assign T181 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T182 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T183 = T185 & T184;
  assign T184 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T185 = T186 & collect_iacq_data;
  assign T186 = state != 3'h0;
  assign T188 = T189 | reset;
  assign T189 = T190 ^ 1'h1;
  assign T190 = T196 & T191;
  assign T191 = T193 | T192;
  assign T192 = 3'h6 == xact_a_type;
  assign T193 = T195 | T194;
  assign T194 = 3'h5 == xact_a_type;
  assign T195 = 3'h4 == xact_a_type;
  assign T196 = T197 & xact_is_builtin_type;
  assign T197 = state != 3'h0;
  assign io_has_release_match = T198;
  assign T198 = T200 & T199;
  assign T199 = state == 3'h1;
  assign T200 = T202 & T201;
  assign T201 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T202 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T203 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T204;
  assign T204 = T205 & collect_iacq_data;
  assign T205 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T206;
  assign T206 = T208 & T207;
  assign T207 = collect_iacq_data ^ 1'h1;
  assign T208 = T210 & T209;
  assign T209 = state != 3'h0;
  assign T210 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T211;
  assign T211 = T144 ? io_inner_grant_ready : pending_ognt_ack;
  assign T500 = reset ? 1'h0 : T212;
  assign T212 = T122 ? 1'h1 : T213;
  assign T213 = T105 ? 1'h1 : T214;
  assign T214 = T215 ? 1'h0 : pending_ognt_ack;
  assign T215 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T216;
  assign T216 = T262 ? oacq_probe_data : T217;
  assign T217 = T261 ? T224 : T218;
  assign T218 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T219;
  assign T219 = T221 | T220;
  assign T220 = 3'h4 == xact_a_type;
  assign T221 = T223 | T222;
  assign T222 = 3'h0 == xact_a_type;
  assign T223 = 3'h2 == xact_a_type;
  assign T224 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T225;
  assign T225 = T260 ? T246 : T226;
  assign T226 = T244 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T227 = T234 ? io_inner_acquire_bits_data : T228;
  assign T228 = T229 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T229 = T233 & T230;
  assign T230 = T231[1'h0:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = io_inner_acquire_bits_addr_beat;
  assign T233 = collect_iacq_data & io_inner_acquire_valid;
  assign T234 = T61 & T235;
  assign T235 = T236[1'h0:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = 2'h0;
  assign T238 = T242 ? io_inner_acquire_bits_data : T239;
  assign T239 = T240 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T240 = T233 & T241;
  assign T241 = T231[1'h1:1'h1];
  assign T242 = T61 & T243;
  assign T243 = T236[1'h1:1'h1];
  assign T244 = T245[1'h0:1'h0];
  assign T245 = oacq_data_cnt;
  assign oacq_data_cnt = T113 ? R109 : 2'h0;
  assign T246 = T259 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T247 = T251 ? io_inner_acquire_bits_data : T248;
  assign T248 = T249 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T249 = T233 & T250;
  assign T250 = T231[2'h2:2'h2];
  assign T251 = T61 & T252;
  assign T252 = T236[2'h2:2'h2];
  assign T253 = T257 ? io_inner_acquire_bits_data : T254;
  assign T254 = T255 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T255 = T233 & T256;
  assign T256 = T231[2'h3:2'h3];
  assign T257 = T61 & T258;
  assign T258 = T236[2'h3:2'h3];
  assign T259 = T245[1'h0:1'h0];
  assign T260 = T245[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T261 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T262 = state == 3'h1;
  assign io_outer_acquire_bits_union = T263;
  assign T263 = T262 ? oacq_probe_union : T264;
  assign T264 = T261 ? T271 : T265;
  assign T265 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T501;
  assign T501 = {4'h0, T266};
  assign T266 = {T267, 6'h0};
  assign T267 = {T270, T268};
  assign T268 = xact_union[4'h8:3'h6];
  assign T269 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T270 = xact_union[4'hc:4'h9];
  assign T271 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T272;
  assign T272 = {T273, 1'h1};
  assign T273 = T345 ? T331 : T274;
  assign T274 = T329 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T275 = T319 ? T300 : T276;
  assign T276 = T296 ? T277 : xact_wmask_buffer_0;
  assign T277 = T294 ? T285 : T278;
  assign T278 = T280 ? T279 : 16'h0;
  assign T279 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T280 = T283 | T281;
  assign T281 = io_inner_acquire_bits_is_builtin_type & T282;
  assign T282 = io_inner_acquire_bits_a_type == 3'h2;
  assign T283 = io_inner_acquire_bits_is_builtin_type & T284;
  assign T284 = io_inner_acquire_bits_a_type == 3'h3;
  assign T285 = T286;
  assign T286 = {T292, T287};
  assign T287 = 8'h0 - T502;
  assign T502 = {7'h0, T288};
  assign T288 = T289[1'h0:1'h0];
  assign T289 = 1'h1 << T290;
  assign T290 = T291[2'h3:2'h3];
  assign T291 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T292 = 8'h0 - T503;
  assign T503 = {7'h0, T293};
  assign T293 = T289[1'h1:1'h1];
  assign T294 = io_inner_acquire_bits_is_builtin_type & T295;
  assign T295 = io_inner_acquire_bits_a_type == 3'h4;
  assign T296 = T233 & T297;
  assign T297 = T298[1'h0:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = io_inner_acquire_bits_addr_beat;
  assign T300 = T317 ? T308 : T301;
  assign T301 = T303 ? T302 : 16'h0;
  assign T302 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T303 = T306 | T304;
  assign T304 = io_inner_acquire_bits_is_builtin_type & T305;
  assign T305 = io_inner_acquire_bits_a_type == 3'h2;
  assign T306 = io_inner_acquire_bits_is_builtin_type & T307;
  assign T307 = io_inner_acquire_bits_a_type == 3'h3;
  assign T308 = T309;
  assign T309 = {T315, T310};
  assign T310 = 8'h0 - T504;
  assign T504 = {7'h0, T311};
  assign T311 = T312[1'h0:1'h0];
  assign T312 = 1'h1 << T313;
  assign T313 = T314[2'h3:2'h3];
  assign T314 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T315 = 8'h0 - T505;
  assign T505 = {7'h0, T316};
  assign T316 = T312[1'h1:1'h1];
  assign T317 = io_inner_acquire_bits_is_builtin_type & T318;
  assign T318 = io_inner_acquire_bits_a_type == 3'h4;
  assign T319 = T61 & T320;
  assign T320 = T321[1'h0:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = 2'h0;
  assign T323 = T327 ? T300 : T324;
  assign T324 = T325 ? T277 : xact_wmask_buffer_1;
  assign T325 = T233 & T326;
  assign T326 = T298[1'h1:1'h1];
  assign T327 = T61 & T328;
  assign T328 = T321[1'h1:1'h1];
  assign T329 = T330[1'h0:1'h0];
  assign T330 = oacq_data_cnt;
  assign T331 = T344 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T332 = T336 ? T300 : T333;
  assign T333 = T334 ? T277 : xact_wmask_buffer_2;
  assign T334 = T233 & T335;
  assign T335 = T298[2'h2:2'h2];
  assign T336 = T61 & T337;
  assign T337 = T321[2'h2:2'h2];
  assign T338 = T342 ? T300 : T339;
  assign T339 = T340 ? T277 : xact_wmask_buffer_3;
  assign T340 = T233 & T341;
  assign T341 = T298[2'h3:2'h3];
  assign T342 = T61 & T343;
  assign T343 = T321[2'h3:2'h3];
  assign T344 = T330[1'h0:1'h0];
  assign T345 = T330[1'h1:1'h1];
  assign oacq_write_beat_union = T346;
  assign T346 = {T347, 1'h1};
  assign T347 = T364 ? T355 : T348;
  assign T348 = T350 ? T349 : 16'h0;
  assign T349 = xact_union[5'h10:1'h1];
  assign T350 = T353 | T351;
  assign T351 = xact_is_builtin_type & T352;
  assign T352 = xact_a_type == 3'h2;
  assign T353 = xact_is_builtin_type & T354;
  assign T354 = xact_a_type == 3'h3;
  assign T355 = T356;
  assign T356 = {T362, T357};
  assign T357 = 8'h0 - T506;
  assign T506 = {7'h0, T358};
  assign T358 = T359[1'h0:1'h0];
  assign T359 = 1'h1 << T360;
  assign T360 = T361[2'h3:2'h3];
  assign T361 = xact_union[4'hc:4'h9];
  assign T362 = 8'h0 - T507;
  assign T507 = {7'h0, T363};
  assign T363 = T359[1'h1:1'h1];
  assign T364 = xact_is_builtin_type & T365;
  assign T365 = xact_a_type == 3'h4;
  assign oacq_probe_union = T366;
  assign T366 = {T367, 1'h1};
  assign T367 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T368;
  assign T368 = T262 ? oacq_probe_a_type : T369;
  assign T369 = T261 ? T371 : T370;
  assign T370 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T371 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T372;
  assign T372 = T262 ? oacq_probe_is_builtin_type : T373;
  assign T373 = T261 ? T375 : T374;
  assign T374 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T375 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T376;
  assign T376 = T262 ? oacq_probe_addr_beat : T377;
  assign T377 = T261 ? T380 : T378;
  assign T378 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T379 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T380 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T381;
  assign T381 = T262 ? oacq_probe_client_xact_id : T382;
  assign T382 = T261 ? T384 : T383;
  assign T383 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 3'h3;
  assign oacq_read_beat_client_xact_id = 3'h3;
  assign T384 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 3'h3;
  assign oacq_write_beat_client_xact_id = 3'h3;
  assign oacq_probe_client_xact_id = 3'h3;
  assign io_outer_acquire_bits_addr_block = T385;
  assign T385 = T262 ? oacq_probe_addr_block : T386;
  assign T386 = T261 ? T388 : T387;
  assign T387 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T388 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T389;
  assign T389 = T126 ? T416 : T390;
  assign T390 = T123 ? T391 : T116;
  assign T391 = T415 & T392;
  assign T392 = T414 | T393;
  assign T393 = T398 & T394;
  assign T394 = T395 - 1'h1;
  assign T395 = 1'h1 << T396;
  assign T396 = T397 + 2'h1;
  assign T397 = oacq_data_cnt - oacq_data_cnt;
  assign T398 = iacq_data_valid >> oacq_data_cnt;
  assign T508 = reset ? 4'h0 : T399;
  assign T399 = T61 ? T407 : T400;
  assign T400 = T233 ? T401 : iacq_data_valid;
  assign T401 = T405 | T402;
  assign T402 = T509 & T403;
  assign T403 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T509 = T404 ? 4'hf : 4'h0;
  assign T404 = 1'h1;
  assign T405 = iacq_data_valid & T406;
  assign T406 = ~ T403;
  assign T407 = T408 << io_inner_acquire_bits_addr_beat;
  assign T408 = io_inner_acquire_bits_is_builtin_type & T409;
  assign T409 = T411 | T410;
  assign T410 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T411 = T413 | T412;
  assign T412 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T413 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T414 = collect_iacq_data ^ 1'h1;
  assign T415 = pending_ognt_ack ^ 1'h1;
  assign T416 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T417;
  assign T417 = T104 ? T418 : 1'h0;
  assign T418 = T419 | io_outer_acquire_ready;
  assign T419 = T420 ^ 1'h1;
  assign T420 = T422 | T421;
  assign T421 = 3'h2 == io_inner_release_bits_r_type;
  assign T422 = T424 | T423;
  assign T423 = 3'h1 == io_inner_release_bits_r_type;
  assign T424 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T425;
  assign T425 = T510;
  assign T510 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T432;
  assign T432 = T433;
  assign T433 = xact_is_builtin_type ? T438 : T434;
  assign T434 = T437 ? 2'h1 : T435;
  assign T435 = T436 ? 2'h0 : 2'h2;
  assign T436 = xact_a_type == 3'h1;
  assign T437 = xact_a_type == 3'h0;
  assign T438 = T451 ? 2'h2 : T439;
  assign T439 = T450 ? 2'h0 : T440;
  assign T440 = T449 ? 2'h2 : T441;
  assign T441 = T448 ? 2'h0 : T442;
  assign T442 = T447 ? 2'h2 : T443;
  assign T443 = T446 ? 2'h0 : T444;
  assign T444 = T445 ? 2'h0 : 2'h2;
  assign T445 = xact_a_type == 3'h4;
  assign T446 = xact_a_type == 3'h6;
  assign T447 = xact_a_type == 3'h5;
  assign T448 = xact_a_type == 3'h2;
  assign T449 = xact_a_type == 3'h0;
  assign T450 = xact_a_type == 3'h3;
  assign T451 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T452;
  assign T452 = xact_addr_block;
  assign io_inner_probe_valid = T453;
  assign T453 = T104 ? T454 : 1'h0;
  assign T454 = pending_probes != 1'h0;
  assign T511 = T512[1'h0:1'h0];
  assign T512 = reset ? 4'h0 : T426;
  assign T426 = T431 ? T514 : T427;
  assign T427 = T93 ? mask_incoherent : T513;
  assign T513 = {3'h0, pending_probes};
  assign T514 = {2'h0, T428};
  assign T428 = T515 & T429;
  assign T429 = ~ T430;
  assign T430 = 1'h1 << 1'h0;
  assign T515 = {1'h0, pending_probes};
  assign T431 = T104 & io_inner_probe_ready;
  assign io_inner_finish_ready = T152;
  assign io_inner_grant_bits_client_id = T455;
  assign T455 = xact_client_id;
  assign io_inner_grant_bits_data = T456;
  assign T456 = 4'h0;
  assign io_inner_grant_bits_g_type = T457;
  assign T457 = T516;
  assign T516 = {1'h0, T458};
  assign T458 = xact_is_builtin_type ? T461 : T517;
  assign T517 = {1'h0, T459};
  assign T459 = T460 ? 2'h0 : 2'h1;
  assign T460 = xact_a_type == 3'h0;
  assign T461 = T474 ? 3'h4 : T462;
  assign T462 = T473 ? 3'h5 : T463;
  assign T463 = T472 ? 3'h3 : T464;
  assign T464 = T471 ? 3'h3 : T465;
  assign T465 = T470 ? 3'h4 : T466;
  assign T466 = T469 ? 3'h1 : T467;
  assign T467 = T468 ? 3'h1 : 3'h3;
  assign T468 = xact_a_type == 3'h6;
  assign T469 = xact_a_type == 3'h5;
  assign T470 = xact_a_type == 3'h4;
  assign T471 = xact_a_type == 3'h3;
  assign T472 = xact_a_type == 3'h2;
  assign T473 = xact_a_type == 3'h1;
  assign T474 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T475;
  assign T475 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T476;
  assign T476 = 3'h3;
  assign io_inner_grant_bits_client_xact_id = T477;
  assign T477 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T478;
  assign T478 = 2'h0;
  assign io_inner_grant_valid = T479;
  assign T479 = T150 ? 1'h1 : T480;
  assign T480 = T144 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T481;
  assign T481 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T187 <= 1'b1;
  if(!T188 && T187 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T177 <= 1'b1;
  if(!T178 && T177 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T153 <= 1'b1;
  if(!T154 && T153 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T151) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= T145;
    end else if(T131) begin
      state <= T127;
    end else if(T124) begin
      state <= 3'h5;
    end else if(T122) begin
      state <= T121;
    end else if(T119) begin
      state <= T117;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T488;
    if(reset) begin
      R109 <= 2'h0;
    end else if(T112) begin
      R109 <= T111;
    end
    if(reset) begin
      R135 <= 2'h0;
    end else if(T138) begin
      R135 <= T137;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T174;
    end else if(T164) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R168 <= 2'h0;
    end else if(T171) begin
      R168 <= T170;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T122) begin
      pending_ognt_ack <= 1'h1;
    end else if(T105) begin
      pending_ognt_ack <= 1'h1;
    end else if(T215) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T234) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T229) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T242) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T240) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T251) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T249) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T257) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T255) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T319) begin
      xact_wmask_buffer_0 <= T300;
    end else if(T296) begin
      xact_wmask_buffer_0 <= T277;
    end
    if(T327) begin
      xact_wmask_buffer_1 <= T300;
    end else if(T325) begin
      xact_wmask_buffer_1 <= T277;
    end
    if(T336) begin
      xact_wmask_buffer_2 <= T300;
    end else if(T334) begin
      xact_wmask_buffer_2 <= T277;
    end
    if(T342) begin
      xact_wmask_buffer_3 <= T300;
    end else if(T340) begin
      xact_wmask_buffer_3 <= T277;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T407;
    end else if(T233) begin
      iacq_data_valid <= T401;
    end
    pending_probes <= T511;
  end
endmodule

module BroadcastAcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [3:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[3:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [3:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[3:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [3:0] io_outer_grant_bits_data,
    output io_has_acquire_conflict,
    output io_has_acquire_match,
    output io_has_release_match
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  reg [2:0] state;
  wire[2:0] T482;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire pending_outer_read_;
  wire T22;
  wire T23;
  wire[3:0] T24;
  wire[3:0] T483;
  wire[2:0] T25;
  wire[2:0] T484;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire[2:0] T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire pending_outer_write_;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] mask_incoherent;
  wire[3:0] T485;
  wire T53;
  wire T54;
  wire[3:0] mask_self;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T486;
  wire T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] T487;
  wire T60;
  wire T61;
  wire T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire pending_outer_read;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire pending_outer_write;
  wire T71;
  wire T72;
  reg [2:0] xact_a_type;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  reg  xact_is_builtin_type;
  wire T77;
  wire T78;
  wire T79;
  reg  release_count;
  wire T488;
  wire[2:0] T489;
  wire[2:0] T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T490;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T491;
  wire T88;
  wire[2:0] T492;
  wire[1:0] T89;
  wire[1:0] T90;
  wire T91;
  wire[1:0] T493;
  wire T92;
  wire T93;
  wire[2:0] T494;
  wire T94;
  wire[2:0] T495;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire oacq_data_done;
  wire T106;
  wire T107;
  wire T108;
  reg [1:0] R109;
  wire[1:0] T496;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  wire[2:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire[2:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire ignt_data_done;
  wire T132;
  wire T133;
  wire T134;
  reg [1:0] R135;
  wire[1:0] T497;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  reg[0:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T158;
  wire T159;
  wire T160;
  wire T161;
  reg  collect_iacq_data;
  wire T498;
  wire T162;
  wire T163;
  wire T164;
  wire iacq_data_done;
  wire T165;
  wire T166;
  wire T167;
  reg [1:0] R168;
  wire[1:0] T499;
  wire[1:0] T169;
  wire[1:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  reg[0:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  reg [1:0] xact_client_id;
  wire[1:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  reg[0:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  reg [25:0] xact_addr_block;
  wire[25:0] T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  reg  pending_ognt_ack;
  wire T500;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] oacq_read_block_data;
  wire[3:0] oacq_read_beat_data;
  wire subblock_type;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire[3:0] T224;
  wire[3:0] oacq_write_block_data;
  wire[3:0] T225;
  wire[3:0] T226;
  reg [3:0] xact_data_buffer_0;
  wire[3:0] T227;
  wire[3:0] T228;
  wire T229;
  wire T230;
  wire[3:0] T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire T235;
  wire[3:0] T236;
  wire[1:0] T237;
  reg [3:0] xact_data_buffer_1;
  wire[3:0] T238;
  wire[3:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire[1:0] T245;
  wire[1:0] oacq_data_cnt;
  wire[3:0] T246;
  reg [3:0] xact_data_buffer_2;
  wire[3:0] T247;
  wire[3:0] T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg [3:0] xact_data_buffer_3;
  wire[3:0] T253;
  wire[3:0] T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[3:0] oacq_write_beat_data;
  wire T261;
  wire[3:0] oacq_probe_data;
  wire T262;
  wire[16:0] T263;
  wire[16:0] T264;
  wire[16:0] T265;
  wire[16:0] oacq_read_block_union;
  wire[16:0] oacq_read_beat_union;
  wire[16:0] T501;
  wire[12:0] T266;
  wire[6:0] T267;
  wire[2:0] T268;
  reg [16:0] xact_union;
  wire[16:0] T269;
  wire[3:0] T270;
  wire[16:0] T271;
  wire[16:0] oacq_write_block_union;
  wire[16:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  reg [15:0] xact_wmask_buffer_0;
  wire[15:0] T275;
  wire[15:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire[15:0] T285;
  wire[15:0] T286;
  wire[7:0] T287;
  wire[7:0] T502;
  wire T288;
  wire[1:0] T289;
  wire T290;
  wire[3:0] T291;
  wire[7:0] T292;
  wire[7:0] T503;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire[3:0] T298;
  wire[1:0] T299;
  wire[15:0] T300;
  wire[15:0] T301;
  wire[15:0] T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[15:0] T308;
  wire[15:0] T309;
  wire[7:0] T310;
  wire[7:0] T504;
  wire T311;
  wire[1:0] T312;
  wire T313;
  wire[3:0] T314;
  wire[7:0] T315;
  wire[7:0] T505;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[1:0] T322;
  reg [15:0] xact_wmask_buffer_1;
  wire[15:0] T323;
  wire[15:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[1:0] T330;
  wire[15:0] T331;
  reg [15:0] xact_wmask_buffer_2;
  wire[15:0] T332;
  wire[15:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  reg [15:0] xact_wmask_buffer_3;
  wire[15:0] T338;
  wire[15:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire[16:0] oacq_write_beat_union;
  wire[16:0] T346;
  wire[15:0] T347;
  wire[15:0] T348;
  wire[15:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire[15:0] T355;
  wire[15:0] T356;
  wire[7:0] T357;
  wire[7:0] T506;
  wire T358;
  wire[1:0] T359;
  wire T360;
  wire[3:0] T361;
  wire[7:0] T362;
  wire[7:0] T507;
  wire T363;
  wire T364;
  wire T365;
  wire[16:0] oacq_probe_union;
  wire[16:0] T366;
  wire[15:0] T367;
  wire[2:0] T368;
  wire[2:0] T369;
  wire[2:0] T370;
  wire[2:0] oacq_read_block_a_type;
  wire[2:0] oacq_read_beat_a_type;
  wire[2:0] T371;
  wire[2:0] oacq_write_block_a_type;
  wire[2:0] oacq_write_beat_a_type;
  wire[2:0] oacq_probe_a_type;
  wire T372;
  wire T373;
  wire T374;
  wire oacq_read_block_is_builtin_type;
  wire oacq_read_beat_is_builtin_type;
  wire T375;
  wire oacq_write_block_is_builtin_type;
  wire oacq_write_beat_is_builtin_type;
  wire oacq_probe_is_builtin_type;
  wire[1:0] T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] oacq_read_block_addr_beat;
  wire[1:0] oacq_read_beat_addr_beat;
  reg [1:0] xact_addr_beat;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] oacq_write_block_addr_beat;
  wire[1:0] oacq_write_beat_addr_beat;
  wire[1:0] oacq_probe_addr_beat;
  wire[2:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire[2:0] oacq_read_block_client_xact_id;
  wire[2:0] oacq_read_beat_client_xact_id;
  wire[2:0] T384;
  wire[2:0] oacq_write_block_client_xact_id;
  wire[2:0] oacq_write_beat_client_xact_id;
  wire[2:0] oacq_probe_client_xact_id;
  wire[25:0] T385;
  wire[25:0] T386;
  wire[25:0] T387;
  wire[25:0] oacq_read_block_addr_block;
  wire[25:0] oacq_read_beat_addr_block;
  wire[25:0] T388;
  wire[25:0] oacq_write_block_addr_block;
  wire[25:0] oacq_write_beat_addr_block;
  wire[25:0] oacq_probe_addr_block;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  reg [3:0] iacq_data_valid;
  wire[3:0] T508;
  wire[3:0] T399;
  wire[3:0] T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[3:0] T509;
  wire T404;
  wire[3:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T510;
  wire[1:0] T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire T436;
  wire T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[25:0] T452;
  wire T453;
  wire T454;
  reg  pending_probes;
  wire T511;
  wire[3:0] T512;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[1:0] T428;
  wire T429;
  wire T430;
  wire[1:0] T515;
  wire T431;
  wire[1:0] T455;
  wire[3:0] T456;
  wire[3:0] T457;
  wire[3:0] T516;
  wire[2:0] T458;
  wire[2:0] T517;
  wire[1:0] T459;
  wire T460;
  wire[2:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire[2:0] T466;
  wire[2:0] T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[2:0] T476;
  wire[1:0] T477;
  wire[1:0] T478;
  wire T479;
  wire T480;
  wire T481;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    xact_is_builtin_type = {1{$random}};
    release_count = {1{$random}};
    R109 = {1{$random}};
    R135 = {1{$random}};
    T153 = 1'b0;
    xact_client_xact_id = {1{$random}};
    collect_iacq_data = {1{$random}};
    R168 = {1{$random}};
    T177 = 1'b0;
    xact_client_id = {1{$random}};
    T187 = 1'b0;
    xact_addr_block = {1{$random}};
    pending_ognt_ack = {1{$random}};
    xact_data_buffer_0 = {1{$random}};
    xact_data_buffer_1 = {1{$random}};
    xact_data_buffer_2 = {1{$random}};
    xact_data_buffer_3 = {1{$random}};
    xact_union = {1{$random}};
    xact_wmask_buffer_0 = {1{$random}};
    xact_wmask_buffer_1 = {1{$random}};
    xact_wmask_buffer_2 = {1{$random}};
    xact_wmask_buffer_3 = {1{$random}};
    xact_addr_beat = {1{$random}};
    iacq_data_valid = {1{$random}};
    pending_probes = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 & T4;
  assign T4 = io_inner_acquire_bits_addr_beat != 2'h0;
  assign T5 = T8 & T6;
  assign T6 = io_inner_acquire_bits_is_builtin_type & T7;
  assign T7 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T8 = T10 & T9;
  assign T9 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T10 = state == 3'h0;
  assign T482 = reset ? 3'h0 : T11;
  assign T11 = T151 ? 3'h0 : T12;
  assign T12 = T149 ? T145 : T13;
  assign T13 = T131 ? T127 : T14;
  assign T14 = T124 ? 3'h5 : T15;
  assign T15 = T122 ? T121 : T16;
  assign T16 = T119 ? T117 : T17;
  assign T17 = T78 ? T63 : T18;
  assign T18 = T61 ? T19 : state;
  assign T19 = T52 ? 3'h1 : T20;
  assign T20 = pending_outer_write_ ? 3'h3 : T21;
  assign T21 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign pending_outer_read_ = T46 ? T43 : T22;
  assign T22 = T42 | T23;
  assign T23 = 4'h1 == T24;
  assign T24 = T483;
  assign T483 = {1'h0, T25};
  assign T25 = io_inner_acquire_bits_is_builtin_type ? T28 : T484;
  assign T484 = {1'h0, T26};
  assign T26 = T27 ? 2'h0 : 2'h1;
  assign T27 = io_inner_acquire_bits_a_type == 3'h0;
  assign T28 = T41 ? 3'h4 : T29;
  assign T29 = T40 ? 3'h5 : T30;
  assign T30 = T39 ? 3'h3 : T31;
  assign T31 = T38 ? 3'h3 : T32;
  assign T32 = T37 ? 3'h4 : T33;
  assign T33 = T36 ? 3'h1 : T34;
  assign T34 = T35 ? 3'h1 : 3'h3;
  assign T35 = io_inner_acquire_bits_a_type == 3'h6;
  assign T36 = io_inner_acquire_bits_a_type == 3'h5;
  assign T37 = io_inner_acquire_bits_a_type == 3'h4;
  assign T38 = io_inner_acquire_bits_a_type == 3'h3;
  assign T39 = io_inner_acquire_bits_a_type == 3'h2;
  assign T40 = io_inner_acquire_bits_a_type == 3'h1;
  assign T41 = io_inner_acquire_bits_a_type == 3'h0;
  assign T42 = 4'h0 == T24;
  assign T43 = T45 | T44;
  assign T44 = 4'h4 == T24;
  assign T45 = 4'h5 == T24;
  assign T46 = io_inner_acquire_bits_is_builtin_type;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T47;
  assign T47 = T49 | T48;
  assign T48 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T51 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T52 = mask_incoherent != 4'h0;
  assign mask_incoherent = mask_self & T485;
  assign T485 = {3'h0, T53};
  assign T53 = ~ T54;
  assign T54 = io_incoherent_0;
  assign mask_self = T58 | T55;
  assign T55 = T486 & T56;
  assign T56 = 1'h1 << io_inner_acquire_bits_client_id;
  assign T486 = T57 ? 4'hf : 4'h0;
  assign T57 = 1'h0;
  assign T58 = T487 & T59;
  assign T59 = ~ T56;
  assign T487 = {3'h0, T60};
  assign T60 = 1'h1;
  assign T61 = T62 & io_inner_acquire_valid;
  assign T62 = 3'h0 == state;
  assign T63 = pending_outer_write ? 3'h3 : T64;
  assign T64 = pending_outer_read ? 3'h2 : 3'h4;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T68 : T65;
  assign T65 = T67 | T66;
  assign T66 = 4'h1 == io_inner_grant_bits_g_type;
  assign T67 = 4'h0 == io_inner_grant_bits_g_type;
  assign T68 = T70 | T69;
  assign T69 = 4'h4 == io_inner_grant_bits_g_type;
  assign T70 = 4'h5 == io_inner_grant_bits_g_type;
  assign pending_outer_write = xact_is_builtin_type & T71;
  assign T71 = T74 | T72;
  assign T72 = 3'h4 == xact_a_type;
  assign T73 = T61 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign T74 = T76 | T75;
  assign T75 = 3'h3 == xact_a_type;
  assign T76 = 3'h2 == xact_a_type;
  assign T77 = T61 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign T78 = T105 & T79;
  assign T79 = release_count == 1'h1;
  assign T488 = T489[1'h0:1'h0];
  assign T489 = reset ? 3'h0 : T80;
  assign T80 = T96 ? T495 : T81;
  assign T81 = T105 ? T494 : T82;
  assign T82 = T93 ? T83 : T490;
  assign T490 = {2'h0, release_count};
  assign T83 = T492 + T84;
  assign T84 = {1'h0, T85};
  assign T85 = T491 + T86;
  assign T86 = {1'h0, T87};
  assign T87 = mask_incoherent[2'h3:2'h3];
  assign T491 = {1'h0, T88};
  assign T88 = mask_incoherent[2'h2:2'h2];
  assign T492 = {1'h0, T89};
  assign T89 = T493 + T90;
  assign T90 = {1'h0, T91};
  assign T91 = mask_incoherent[1'h1:1'h1];
  assign T493 = {1'h0, T92};
  assign T92 = mask_incoherent[1'h0:1'h0];
  assign T93 = T61 & T52;
  assign T494 = {2'h0, T94};
  assign T94 = release_count - 1'h1;
  assign T495 = {2'h0, T95};
  assign T95 = release_count - 1'h1;
  assign T96 = T103 & T97;
  assign T97 = T98 ^ 1'h1;
  assign T98 = T100 | T99;
  assign T99 = 3'h2 == io_inner_release_bits_r_type;
  assign T100 = T102 | T101;
  assign T101 = 3'h1 == io_inner_release_bits_r_type;
  assign T102 = 3'h0 == io_inner_release_bits_r_type;
  assign T103 = T104 & io_inner_release_valid;
  assign T104 = 3'h1 == state;
  assign T105 = T115 & oacq_data_done;
  assign oacq_data_done = T113 ? T107 : T106;
  assign T106 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T107 = T112 & T108;
  assign T108 = R109 == 2'h3;
  assign T496 = reset ? 2'h0 : T110;
  assign T110 = T112 ? T111 : R109;
  assign T111 = R109 + 2'h1;
  assign T112 = T106 & T113;
  assign T113 = io_outer_acquire_bits_is_builtin_type & T114;
  assign T114 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T115 = T116 & io_outer_acquire_ready;
  assign T116 = T103 & T98;
  assign T117 = pending_outer_write ? 3'h3 : T118;
  assign T118 = pending_outer_read ? 3'h2 : 3'h4;
  assign T119 = T96 & T120;
  assign T120 = release_count == 1'h1;
  assign T121 = pending_outer_read ? 3'h2 : 3'h5;
  assign T122 = T123 & oacq_data_done;
  assign T123 = 3'h3 == state;
  assign T124 = T126 & T125;
  assign T125 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T126 = 3'h2 == state;
  assign T127 = T128 ? 3'h6 : 3'h0;
  assign T128 = T129 ^ 1'h1;
  assign T129 = io_inner_grant_bits_is_builtin_type & T130;
  assign T130 = io_inner_grant_bits_g_type == 4'h0;
  assign T131 = T144 & ignt_data_done;
  assign ignt_data_done = T139 ? T133 : T132;
  assign T132 = io_inner_grant_ready & io_inner_grant_valid;
  assign T133 = T138 & T134;
  assign T134 = R135 == 2'h3;
  assign T497 = reset ? 2'h0 : T136;
  assign T136 = T138 ? T137 : R135;
  assign T137 = R135 + 2'h1;
  assign T138 = T132 & T139;
  assign T139 = io_inner_grant_bits_is_builtin_type ? T143 : T140;
  assign T140 = T142 | T141;
  assign T141 = 4'h1 == io_inner_grant_bits_g_type;
  assign T142 = 4'h0 == io_inner_grant_bits_g_type;
  assign T143 = 4'h5 == io_inner_grant_bits_g_type;
  assign T144 = 3'h5 == state;
  assign T145 = T146 ? 3'h6 : 3'h0;
  assign T146 = T147 ^ 1'h1;
  assign T147 = io_inner_grant_bits_is_builtin_type & T148;
  assign T148 = io_inner_grant_bits_g_type == 4'h0;
  assign T149 = T150 & io_inner_grant_ready;
  assign T150 = 3'h4 == state;
  assign T151 = T152 & io_inner_finish_valid;
  assign T152 = 3'h6 == state;
  assign T154 = T155 | reset;
  assign T155 = T156 ^ 1'h1;
  assign T156 = T159 & T157;
  assign T157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T158 = T61 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign T159 = T161 & T160;
  assign T160 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T161 = T176 & collect_iacq_data;
  assign T498 = reset ? 1'h0 : T162;
  assign T162 = T61 ? T174 : T163;
  assign T163 = T164 ? 1'h0 : collect_iacq_data;
  assign T164 = collect_iacq_data & iacq_data_done;
  assign iacq_data_done = T172 ? T166 : T165;
  assign T165 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T166 = T171 & T167;
  assign T167 = R168 == 2'h3;
  assign T499 = reset ? 2'h0 : T169;
  assign T169 = T171 ? T170 : R168;
  assign T170 = R168 + 2'h1;
  assign T171 = T165 & T172;
  assign T172 = io_inner_acquire_bits_is_builtin_type & T173;
  assign T173 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T174 = io_inner_acquire_bits_is_builtin_type & T175;
  assign T175 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T176 = state != 3'h0;
  assign T178 = T179 | reset;
  assign T179 = T180 ^ 1'h1;
  assign T180 = T183 & T181;
  assign T181 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T182 = T61 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign T183 = T185 & T184;
  assign T184 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T185 = T186 & collect_iacq_data;
  assign T186 = state != 3'h0;
  assign T188 = T189 | reset;
  assign T189 = T190 ^ 1'h1;
  assign T190 = T196 & T191;
  assign T191 = T193 | T192;
  assign T192 = 3'h6 == xact_a_type;
  assign T193 = T195 | T194;
  assign T194 = 3'h5 == xact_a_type;
  assign T195 = 3'h4 == xact_a_type;
  assign T196 = T197 & xact_is_builtin_type;
  assign T197 = state != 3'h0;
  assign io_has_release_match = T198;
  assign T198 = T200 & T199;
  assign T199 = state == 3'h1;
  assign T200 = T202 & T201;
  assign T201 = io_inner_release_bits_voluntary ^ 1'h1;
  assign T202 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T203 = T61 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign io_has_acquire_match = T204;
  assign T204 = T205 & collect_iacq_data;
  assign T205 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_has_acquire_conflict = T206;
  assign T206 = T208 & T207;
  assign T207 = collect_iacq_data ^ 1'h1;
  assign T208 = T210 & T209;
  assign T209 = state != 3'h0;
  assign T210 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign io_outer_grant_ready = T211;
  assign T211 = T144 ? io_inner_grant_ready : pending_ognt_ack;
  assign T500 = reset ? 1'h0 : T212;
  assign T212 = T122 ? 1'h1 : T213;
  assign T213 = T105 ? 1'h1 : T214;
  assign T214 = T215 ? 1'h0 : pending_ognt_ack;
  assign T215 = pending_ognt_ack & io_outer_grant_valid;
  assign io_outer_acquire_bits_data = T216;
  assign T216 = T262 ? oacq_probe_data : T217;
  assign T217 = T261 ? T224 : T218;
  assign T218 = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign oacq_read_block_data = 4'h0;
  assign oacq_read_beat_data = 4'h0;
  assign subblock_type = xact_is_builtin_type & T219;
  assign T219 = T221 | T220;
  assign T220 = 3'h4 == xact_a_type;
  assign T221 = T223 | T222;
  assign T222 = 3'h0 == xact_a_type;
  assign T223 = 3'h2 == xact_a_type;
  assign T224 = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign oacq_write_block_data = T225;
  assign T225 = T260 ? T246 : T226;
  assign T226 = T244 ? xact_data_buffer_1 : xact_data_buffer_0;
  assign T227 = T234 ? io_inner_acquire_bits_data : T228;
  assign T228 = T229 ? io_inner_acquire_bits_data : xact_data_buffer_0;
  assign T229 = T233 & T230;
  assign T230 = T231[1'h0:1'h0];
  assign T231 = 1'h1 << T232;
  assign T232 = io_inner_acquire_bits_addr_beat;
  assign T233 = collect_iacq_data & io_inner_acquire_valid;
  assign T234 = T61 & T235;
  assign T235 = T236[1'h0:1'h0];
  assign T236 = 1'h1 << T237;
  assign T237 = 2'h0;
  assign T238 = T242 ? io_inner_acquire_bits_data : T239;
  assign T239 = T240 ? io_inner_acquire_bits_data : xact_data_buffer_1;
  assign T240 = T233 & T241;
  assign T241 = T231[1'h1:1'h1];
  assign T242 = T61 & T243;
  assign T243 = T236[1'h1:1'h1];
  assign T244 = T245[1'h0:1'h0];
  assign T245 = oacq_data_cnt;
  assign oacq_data_cnt = T113 ? R109 : 2'h0;
  assign T246 = T259 ? xact_data_buffer_3 : xact_data_buffer_2;
  assign T247 = T251 ? io_inner_acquire_bits_data : T248;
  assign T248 = T249 ? io_inner_acquire_bits_data : xact_data_buffer_2;
  assign T249 = T233 & T250;
  assign T250 = T231[2'h2:2'h2];
  assign T251 = T61 & T252;
  assign T252 = T236[2'h2:2'h2];
  assign T253 = T257 ? io_inner_acquire_bits_data : T254;
  assign T254 = T255 ? io_inner_acquire_bits_data : xact_data_buffer_3;
  assign T255 = T233 & T256;
  assign T256 = T231[2'h3:2'h3];
  assign T257 = T61 & T258;
  assign T258 = T236[2'h3:2'h3];
  assign T259 = T245[1'h0:1'h0];
  assign T260 = T245[1'h1:1'h1];
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign T261 = state == 3'h3;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T262 = state == 3'h1;
  assign io_outer_acquire_bits_union = T263;
  assign T263 = T262 ? oacq_probe_union : T264;
  assign T264 = T261 ? T271 : T265;
  assign T265 = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign oacq_read_block_union = 17'h1c1;
  assign oacq_read_beat_union = T501;
  assign T501 = {4'h0, T266};
  assign T266 = {T267, 6'h0};
  assign T267 = {T270, T268};
  assign T268 = xact_union[4'h8:3'h6];
  assign T269 = T61 ? io_inner_acquire_bits_union : xact_union;
  assign T270 = xact_union[4'hc:4'h9];
  assign T271 = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign oacq_write_block_union = T272;
  assign T272 = {T273, 1'h1};
  assign T273 = T345 ? T331 : T274;
  assign T274 = T329 ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign T275 = T319 ? T300 : T276;
  assign T276 = T296 ? T277 : xact_wmask_buffer_0;
  assign T277 = T294 ? T285 : T278;
  assign T278 = T280 ? T279 : 16'h0;
  assign T279 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T280 = T283 | T281;
  assign T281 = io_inner_acquire_bits_is_builtin_type & T282;
  assign T282 = io_inner_acquire_bits_a_type == 3'h2;
  assign T283 = io_inner_acquire_bits_is_builtin_type & T284;
  assign T284 = io_inner_acquire_bits_a_type == 3'h3;
  assign T285 = T286;
  assign T286 = {T292, T287};
  assign T287 = 8'h0 - T502;
  assign T502 = {7'h0, T288};
  assign T288 = T289[1'h0:1'h0];
  assign T289 = 1'h1 << T290;
  assign T290 = T291[2'h3:2'h3];
  assign T291 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T292 = 8'h0 - T503;
  assign T503 = {7'h0, T293};
  assign T293 = T289[1'h1:1'h1];
  assign T294 = io_inner_acquire_bits_is_builtin_type & T295;
  assign T295 = io_inner_acquire_bits_a_type == 3'h4;
  assign T296 = T233 & T297;
  assign T297 = T298[1'h0:1'h0];
  assign T298 = 1'h1 << T299;
  assign T299 = io_inner_acquire_bits_addr_beat;
  assign T300 = T317 ? T308 : T301;
  assign T301 = T303 ? T302 : 16'h0;
  assign T302 = io_inner_acquire_bits_union[5'h10:1'h1];
  assign T303 = T306 | T304;
  assign T304 = io_inner_acquire_bits_is_builtin_type & T305;
  assign T305 = io_inner_acquire_bits_a_type == 3'h2;
  assign T306 = io_inner_acquire_bits_is_builtin_type & T307;
  assign T307 = io_inner_acquire_bits_a_type == 3'h3;
  assign T308 = T309;
  assign T309 = {T315, T310};
  assign T310 = 8'h0 - T504;
  assign T504 = {7'h0, T311};
  assign T311 = T312[1'h0:1'h0];
  assign T312 = 1'h1 << T313;
  assign T313 = T314[2'h3:2'h3];
  assign T314 = io_inner_acquire_bits_union[4'hc:4'h9];
  assign T315 = 8'h0 - T505;
  assign T505 = {7'h0, T316};
  assign T316 = T312[1'h1:1'h1];
  assign T317 = io_inner_acquire_bits_is_builtin_type & T318;
  assign T318 = io_inner_acquire_bits_a_type == 3'h4;
  assign T319 = T61 & T320;
  assign T320 = T321[1'h0:1'h0];
  assign T321 = 1'h1 << T322;
  assign T322 = 2'h0;
  assign T323 = T327 ? T300 : T324;
  assign T324 = T325 ? T277 : xact_wmask_buffer_1;
  assign T325 = T233 & T326;
  assign T326 = T298[1'h1:1'h1];
  assign T327 = T61 & T328;
  assign T328 = T321[1'h1:1'h1];
  assign T329 = T330[1'h0:1'h0];
  assign T330 = oacq_data_cnt;
  assign T331 = T344 ? xact_wmask_buffer_3 : xact_wmask_buffer_2;
  assign T332 = T336 ? T300 : T333;
  assign T333 = T334 ? T277 : xact_wmask_buffer_2;
  assign T334 = T233 & T335;
  assign T335 = T298[2'h2:2'h2];
  assign T336 = T61 & T337;
  assign T337 = T321[2'h2:2'h2];
  assign T338 = T342 ? T300 : T339;
  assign T339 = T340 ? T277 : xact_wmask_buffer_3;
  assign T340 = T233 & T341;
  assign T341 = T298[2'h3:2'h3];
  assign T342 = T61 & T343;
  assign T343 = T321[2'h3:2'h3];
  assign T344 = T330[1'h0:1'h0];
  assign T345 = T330[1'h1:1'h1];
  assign oacq_write_beat_union = T346;
  assign T346 = {T347, 1'h1};
  assign T347 = T364 ? T355 : T348;
  assign T348 = T350 ? T349 : 16'h0;
  assign T349 = xact_union[5'h10:1'h1];
  assign T350 = T353 | T351;
  assign T351 = xact_is_builtin_type & T352;
  assign T352 = xact_a_type == 3'h2;
  assign T353 = xact_is_builtin_type & T354;
  assign T354 = xact_a_type == 3'h3;
  assign T355 = T356;
  assign T356 = {T362, T357};
  assign T357 = 8'h0 - T506;
  assign T506 = {7'h0, T358};
  assign T358 = T359[1'h0:1'h0];
  assign T359 = 1'h1 << T360;
  assign T360 = T361[2'h3:2'h3];
  assign T361 = xact_union[4'hc:4'h9];
  assign T362 = 8'h0 - T507;
  assign T507 = {7'h0, T363};
  assign T363 = T359[1'h1:1'h1];
  assign T364 = xact_is_builtin_type & T365;
  assign T365 = xact_a_type == 3'h4;
  assign oacq_probe_union = T366;
  assign T366 = {T367, 1'h1};
  assign T367 = 16'hffff;
  assign io_outer_acquire_bits_a_type = T368;
  assign T368 = T262 ? oacq_probe_a_type : T369;
  assign T369 = T261 ? T371 : T370;
  assign T370 = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign T371 = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_probe_a_type = 3'h3;
  assign io_outer_acquire_bits_is_builtin_type = T372;
  assign T372 = T262 ? oacq_probe_is_builtin_type : T373;
  assign T373 = T261 ? T375 : T374;
  assign T374 = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign T375 = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign io_outer_acquire_bits_addr_beat = T376;
  assign T376 = T262 ? oacq_probe_addr_beat : T377;
  assign T377 = T261 ? T380 : T378;
  assign T378 = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign oacq_read_block_addr_beat = 2'h0;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign T379 = T61 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign T380 = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = T381;
  assign T381 = T262 ? oacq_probe_client_xact_id : T382;
  assign T382 = T261 ? T384 : T383;
  assign T383 = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign oacq_read_block_client_xact_id = 3'h4;
  assign oacq_read_beat_client_xact_id = 3'h4;
  assign T384 = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign oacq_write_block_client_xact_id = 3'h4;
  assign oacq_write_beat_client_xact_id = 3'h4;
  assign oacq_probe_client_xact_id = 3'h4;
  assign io_outer_acquire_bits_addr_block = T385;
  assign T385 = T262 ? oacq_probe_addr_block : T386;
  assign T386 = T261 ? T388 : T387;
  assign T387 = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign T388 = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_acquire_valid = T389;
  assign T389 = T126 ? T416 : T390;
  assign T390 = T123 ? T391 : T116;
  assign T391 = T415 & T392;
  assign T392 = T414 | T393;
  assign T393 = T398 & T394;
  assign T394 = T395 - 1'h1;
  assign T395 = 1'h1 << T396;
  assign T396 = T397 + 2'h1;
  assign T397 = oacq_data_cnt - oacq_data_cnt;
  assign T398 = iacq_data_valid >> oacq_data_cnt;
  assign T508 = reset ? 4'h0 : T399;
  assign T399 = T61 ? T407 : T400;
  assign T400 = T233 ? T401 : iacq_data_valid;
  assign T401 = T405 | T402;
  assign T402 = T509 & T403;
  assign T403 = 1'h1 << io_inner_acquire_bits_addr_beat;
  assign T509 = T404 ? 4'hf : 4'h0;
  assign T404 = 1'h1;
  assign T405 = iacq_data_valid & T406;
  assign T406 = ~ T403;
  assign T407 = T408 << io_inner_acquire_bits_addr_beat;
  assign T408 = io_inner_acquire_bits_is_builtin_type & T409;
  assign T409 = T411 | T410;
  assign T410 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T411 = T413 | T412;
  assign T412 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T413 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T414 = collect_iacq_data ^ 1'h1;
  assign T415 = pending_ognt_ack ^ 1'h1;
  assign T416 = pending_ognt_ack ^ 1'h1;
  assign io_inner_release_ready = T417;
  assign T417 = T104 ? T418 : 1'h0;
  assign T418 = T419 | io_outer_acquire_ready;
  assign T419 = T420 ^ 1'h1;
  assign T420 = T422 | T421;
  assign T421 = 3'h2 == io_inner_release_bits_r_type;
  assign T422 = T424 | T423;
  assign T423 = 3'h1 == io_inner_release_bits_r_type;
  assign T424 = 3'h0 == io_inner_release_bits_r_type;
  assign io_inner_probe_bits_client_id = T425;
  assign T425 = T510;
  assign T510 = {1'h0, 1'h0};
  assign io_inner_probe_bits_p_type = T432;
  assign T432 = T433;
  assign T433 = xact_is_builtin_type ? T438 : T434;
  assign T434 = T437 ? 2'h1 : T435;
  assign T435 = T436 ? 2'h0 : 2'h2;
  assign T436 = xact_a_type == 3'h1;
  assign T437 = xact_a_type == 3'h0;
  assign T438 = T451 ? 2'h2 : T439;
  assign T439 = T450 ? 2'h0 : T440;
  assign T440 = T449 ? 2'h2 : T441;
  assign T441 = T448 ? 2'h0 : T442;
  assign T442 = T447 ? 2'h2 : T443;
  assign T443 = T446 ? 2'h0 : T444;
  assign T444 = T445 ? 2'h0 : 2'h2;
  assign T445 = xact_a_type == 3'h4;
  assign T446 = xact_a_type == 3'h6;
  assign T447 = xact_a_type == 3'h5;
  assign T448 = xact_a_type == 3'h2;
  assign T449 = xact_a_type == 3'h0;
  assign T450 = xact_a_type == 3'h3;
  assign T451 = xact_a_type == 3'h1;
  assign io_inner_probe_bits_addr_block = T452;
  assign T452 = xact_addr_block;
  assign io_inner_probe_valid = T453;
  assign T453 = T104 ? T454 : 1'h0;
  assign T454 = pending_probes != 1'h0;
  assign T511 = T512[1'h0:1'h0];
  assign T512 = reset ? 4'h0 : T426;
  assign T426 = T431 ? T514 : T427;
  assign T427 = T93 ? mask_incoherent : T513;
  assign T513 = {3'h0, pending_probes};
  assign T514 = {2'h0, T428};
  assign T428 = T515 & T429;
  assign T429 = ~ T430;
  assign T430 = 1'h1 << 1'h0;
  assign T515 = {1'h0, pending_probes};
  assign T431 = T104 & io_inner_probe_ready;
  assign io_inner_finish_ready = T152;
  assign io_inner_grant_bits_client_id = T455;
  assign T455 = xact_client_id;
  assign io_inner_grant_bits_data = T456;
  assign T456 = 4'h0;
  assign io_inner_grant_bits_g_type = T457;
  assign T457 = T516;
  assign T516 = {1'h0, T458};
  assign T458 = xact_is_builtin_type ? T461 : T517;
  assign T517 = {1'h0, T459};
  assign T459 = T460 ? 2'h0 : 2'h1;
  assign T460 = xact_a_type == 3'h0;
  assign T461 = T474 ? 3'h4 : T462;
  assign T462 = T473 ? 3'h5 : T463;
  assign T463 = T472 ? 3'h3 : T464;
  assign T464 = T471 ? 3'h3 : T465;
  assign T465 = T470 ? 3'h4 : T466;
  assign T466 = T469 ? 3'h1 : T467;
  assign T467 = T468 ? 3'h1 : 3'h3;
  assign T468 = xact_a_type == 3'h6;
  assign T469 = xact_a_type == 3'h5;
  assign T470 = xact_a_type == 3'h4;
  assign T471 = xact_a_type == 3'h3;
  assign T472 = xact_a_type == 3'h2;
  assign T473 = xact_a_type == 3'h1;
  assign T474 = xact_a_type == 3'h0;
  assign io_inner_grant_bits_is_builtin_type = T475;
  assign T475 = xact_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = T476;
  assign T476 = 3'h4;
  assign io_inner_grant_bits_client_xact_id = T477;
  assign T477 = xact_client_xact_id;
  assign io_inner_grant_bits_addr_beat = T478;
  assign T478 = 2'h0;
  assign io_inner_grant_valid = T479;
  assign T479 = T150 ? 1'h1 : T480;
  assign T480 = T144 ? io_outer_grant_valid : 1'h0;
  assign io_inner_acquire_ready = T481;
  assign T481 = T62 ? 1'h1 : collect_iacq_data;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T187 <= 1'b1;
  if(!T188 && T187 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Broadcast Hub does not support PutAtomics or prefetches");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T177 <= 1'b1;
  if(!T178 && T177 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different network source than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T153 <= 1'b1;
  if(!T154 && T153 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker accepted data beat from different client transaction than initial request.");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "AcquireTracker initialized with a tail data beat.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T151) begin
      state <= 3'h0;
    end else if(T149) begin
      state <= T145;
    end else if(T131) begin
      state <= T127;
    end else if(T124) begin
      state <= 3'h5;
    end else if(T122) begin
      state <= T121;
    end else if(T119) begin
      state <= T117;
    end else if(T78) begin
      state <= T63;
    end else if(T61) begin
      state <= T19;
    end
    if(T61) begin
      xact_a_type <= io_inner_acquire_bits_a_type;
    end
    if(T61) begin
      xact_is_builtin_type <= io_inner_acquire_bits_is_builtin_type;
    end
    release_count <= T488;
    if(reset) begin
      R109 <= 2'h0;
    end else if(T112) begin
      R109 <= T111;
    end
    if(reset) begin
      R135 <= 2'h0;
    end else if(T138) begin
      R135 <= T137;
    end
    if(T61) begin
      xact_client_xact_id <= io_inner_acquire_bits_client_xact_id;
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else if(T61) begin
      collect_iacq_data <= T174;
    end else if(T164) begin
      collect_iacq_data <= 1'h0;
    end
    if(reset) begin
      R168 <= 2'h0;
    end else if(T171) begin
      R168 <= T170;
    end
    if(T61) begin
      xact_client_id <= io_inner_acquire_bits_client_id;
    end
    if(T61) begin
      xact_addr_block <= io_inner_acquire_bits_addr_block;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else if(T122) begin
      pending_ognt_ack <= 1'h1;
    end else if(T105) begin
      pending_ognt_ack <= 1'h1;
    end else if(T215) begin
      pending_ognt_ack <= 1'h0;
    end
    if(T234) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end else if(T229) begin
      xact_data_buffer_0 <= io_inner_acquire_bits_data;
    end
    if(T242) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end else if(T240) begin
      xact_data_buffer_1 <= io_inner_acquire_bits_data;
    end
    if(T251) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end else if(T249) begin
      xact_data_buffer_2 <= io_inner_acquire_bits_data;
    end
    if(T257) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end else if(T255) begin
      xact_data_buffer_3 <= io_inner_acquire_bits_data;
    end
    if(T61) begin
      xact_union <= io_inner_acquire_bits_union;
    end
    if(T319) begin
      xact_wmask_buffer_0 <= T300;
    end else if(T296) begin
      xact_wmask_buffer_0 <= T277;
    end
    if(T327) begin
      xact_wmask_buffer_1 <= T300;
    end else if(T325) begin
      xact_wmask_buffer_1 <= T277;
    end
    if(T336) begin
      xact_wmask_buffer_2 <= T300;
    end else if(T334) begin
      xact_wmask_buffer_2 <= T277;
    end
    if(T342) begin
      xact_wmask_buffer_3 <= T300;
    end else if(T340) begin
      xact_wmask_buffer_3 <= T277;
    end
    if(T61) begin
      xact_addr_beat <= io_inner_acquire_bits_addr_beat;
    end
    if(reset) begin
      iacq_data_valid <= 4'h0;
    end else if(T61) begin
      iacq_data_valid <= T407;
    end else if(T233) begin
      iacq_data_valid <= T401;
    end
    pending_probes <= T511;
  end
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_addr_beat,
    input [1:0] io_in_4_bits_client_xact_id,
    input [2:0] io_in_4_bits_manager_xact_id,
    input  io_in_4_bits_is_builtin_type,
    input [3:0] io_in_4_bits_g_type,
    input [127:0] io_in_4_bits_data,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_addr_beat,
    input [1:0] io_in_3_bits_client_xact_id,
    input [2:0] io_in_3_bits_manager_xact_id,
    input  io_in_3_bits_is_builtin_type,
    input [3:0] io_in_3_bits_g_type,
    input [127:0] io_in_3_bits_data,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_addr_beat,
    input [1:0] io_in_2_bits_client_xact_id,
    input [2:0] io_in_2_bits_manager_xact_id,
    input  io_in_2_bits_is_builtin_type,
    input [3:0] io_in_2_bits_g_type,
    input [127:0] io_in_2_bits_data,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [127:0] io_in_1_bits_data,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [127:0] io_in_0_bits_data,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T192;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T193;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg  locked;
  wire T194;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  reg [1:0] R41;
  wire[1:0] T195;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[2:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire[127:0] T52;
  wire[127:0] T53;
  wire[127:0] T54;
  wire T55;
  wire[127:0] T56;
  wire T57;
  wire T58;
  wire T59;
  wire[3:0] T60;
  wire[3:0] T61;
  wire[3:0] T62;
  wire T63;
  wire[3:0] T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] T86;
  wire T87;
  wire[1:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire[1:0] T92;
  wire[1:0] T93;
  wire[1:0] T94;
  wire T95;
  wire[1:0] T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R41 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T192 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T193 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T35 & T30;
  assign T30 = io_out_bits_is_builtin_type ? T34 : T31;
  assign T31 = T33 | T32;
  assign T32 = 4'h1 == io_out_bits_g_type;
  assign T33 = 4'h0 == io_out_bits_g_type;
  assign T34 = 4'h5 == io_out_bits_g_type;
  assign T35 = io_out_ready & io_out_valid;
  assign T194 = reset ? 1'h0 : T36;
  assign T36 = T38 ? 1'h0 : T37;
  assign T37 = T27 ? 1'h1 : locked;
  assign T38 = T35 & T39;
  assign T39 = T40 == 2'h0;
  assign T40 = R41 + 2'h1;
  assign T195 = reset ? 2'h0 : T42;
  assign T42 = T29 ? T40 : R41;
  assign io_out_bits_client_id = T43;
  assign T43 = T51 ? io_in_4_bits_client_id : T44;
  assign T44 = T50 ? T48 : T45;
  assign T45 = T46 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T46 = T47[1'h0:1'h0];
  assign T47 = chosen;
  assign T48 = T49 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T49 = T47[1'h0:1'h0];
  assign T50 = T47[1'h1:1'h1];
  assign T51 = T47[2'h2:2'h2];
  assign io_out_bits_data = T52;
  assign T52 = T59 ? io_in_4_bits_data : T53;
  assign T53 = T58 ? T56 : T54;
  assign T54 = T55 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T55 = T47[1'h0:1'h0];
  assign T56 = T57 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T57 = T47[1'h0:1'h0];
  assign T58 = T47[1'h1:1'h1];
  assign T59 = T47[2'h2:2'h2];
  assign io_out_bits_g_type = T60;
  assign T60 = T67 ? io_in_4_bits_g_type : T61;
  assign T61 = T66 ? T64 : T62;
  assign T62 = T63 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign T63 = T47[1'h0:1'h0];
  assign T64 = T65 ? io_in_3_bits_g_type : io_in_2_bits_g_type;
  assign T65 = T47[1'h0:1'h0];
  assign T66 = T47[1'h1:1'h1];
  assign T67 = T47[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T68;
  assign T68 = T75 ? io_in_4_bits_is_builtin_type : T69;
  assign T69 = T74 ? T72 : T70;
  assign T70 = T71 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T71 = T47[1'h0:1'h0];
  assign T72 = T73 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T73 = T47[1'h0:1'h0];
  assign T74 = T47[1'h1:1'h1];
  assign T75 = T47[2'h2:2'h2];
  assign io_out_bits_manager_xact_id = T76;
  assign T76 = T83 ? io_in_4_bits_manager_xact_id : T77;
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign T79 = T47[1'h0:1'h0];
  assign T80 = T81 ? io_in_3_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign T81 = T47[1'h0:1'h0];
  assign T82 = T47[1'h1:1'h1];
  assign T83 = T47[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T84;
  assign T84 = T91 ? io_in_4_bits_client_xact_id : T85;
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T87 = T47[1'h0:1'h0];
  assign T88 = T89 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T89 = T47[1'h0:1'h0];
  assign T90 = T47[1'h1:1'h1];
  assign T91 = T47[2'h2:2'h2];
  assign io_out_bits_addr_beat = T92;
  assign T92 = T99 ? io_in_4_bits_addr_beat : T93;
  assign T93 = T98 ? T96 : T94;
  assign T94 = T95 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T95 = T47[1'h0:1'h0];
  assign T96 = T97 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T97 = T47[1'h0:1'h0];
  assign T98 = T47[1'h1:1'h1];
  assign T99 = T47[2'h2:2'h2];
  assign io_out_valid = T100;
  assign T100 = T107 ? io_in_4_valid : T101;
  assign T101 = T106 ? T104 : T102;
  assign T102 = T103 ? io_in_1_valid : io_in_0_valid;
  assign T103 = T47[1'h0:1'h0];
  assign T104 = T105 ? io_in_3_valid : io_in_2_valid;
  assign T105 = T47[1'h0:1'h0];
  assign T106 = T47[1'h1:1'h1];
  assign T107 = T47[2'h2:2'h2];
  assign io_in_0_ready = T108;
  assign T108 = T109 & io_out_ready;
  assign T109 = locked ? T127 : T110;
  assign T110 = T126 | T111;
  assign T111 = T112 ^ 1'h1;
  assign T112 = T115 | T113;
  assign T113 = io_in_4_valid & T114;
  assign T114 = last_grant < 3'h4;
  assign T115 = T118 | T116;
  assign T116 = io_in_3_valid & T117;
  assign T117 = last_grant < 3'h3;
  assign T118 = T121 | T119;
  assign T119 = io_in_2_valid & T120;
  assign T120 = last_grant < 3'h2;
  assign T121 = T124 | T122;
  assign T122 = io_in_1_valid & T123;
  assign T123 = last_grant < 3'h1;
  assign T124 = io_in_0_valid & T125;
  assign T125 = last_grant < 3'h0;
  assign T126 = last_grant < 3'h0;
  assign T127 = lockIdx == 3'h0;
  assign io_in_1_ready = T128;
  assign T128 = T129 & io_out_ready;
  assign T129 = locked ? T140 : T130;
  assign T130 = T137 | T131;
  assign T131 = T132 ^ 1'h1;
  assign T132 = T133 | io_in_0_valid;
  assign T133 = T134 | T113;
  assign T134 = T135 | T116;
  assign T135 = T136 | T119;
  assign T136 = T124 | T122;
  assign T137 = T139 & T138;
  assign T138 = last_grant < 3'h1;
  assign T139 = T124 ^ 1'h1;
  assign T140 = lockIdx == 3'h1;
  assign io_in_2_ready = T141;
  assign T141 = T142 & io_out_ready;
  assign T142 = locked ? T155 : T143;
  assign T143 = T151 | T144;
  assign T144 = T145 ^ 1'h1;
  assign T145 = T146 | io_in_1_valid;
  assign T146 = T147 | io_in_0_valid;
  assign T147 = T148 | T113;
  assign T148 = T149 | T116;
  assign T149 = T150 | T119;
  assign T150 = T124 | T122;
  assign T151 = T153 & T152;
  assign T152 = last_grant < 3'h2;
  assign T153 = T154 ^ 1'h1;
  assign T154 = T124 | T122;
  assign T155 = lockIdx == 3'h2;
  assign io_in_3_ready = T156;
  assign T156 = T157 & io_out_ready;
  assign T157 = locked ? T172 : T158;
  assign T158 = T167 | T159;
  assign T159 = T160 ^ 1'h1;
  assign T160 = T161 | io_in_2_valid;
  assign T161 = T162 | io_in_1_valid;
  assign T162 = T163 | io_in_0_valid;
  assign T163 = T164 | T113;
  assign T164 = T165 | T116;
  assign T165 = T166 | T119;
  assign T166 = T124 | T122;
  assign T167 = T169 & T168;
  assign T168 = last_grant < 3'h3;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T171 | T119;
  assign T171 = T124 | T122;
  assign T172 = lockIdx == 3'h3;
  assign io_in_4_ready = T173;
  assign T173 = T174 & io_out_ready;
  assign T174 = locked ? T191 : T175;
  assign T175 = T185 | T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T178 | io_in_3_valid;
  assign T178 = T179 | io_in_2_valid;
  assign T179 = T180 | io_in_1_valid;
  assign T180 = T181 | io_in_0_valid;
  assign T181 = T182 | T113;
  assign T182 = T183 | T116;
  assign T183 = T184 | T119;
  assign T184 = T124 | T122;
  assign T185 = T187 & T186;
  assign T186 = last_grant < 3'h4;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T189 | T116;
  assign T189 = T190 | T119;
  assign T190 = T124 | T122;
  assign T191 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T38) begin
      locked <= 1'h0;
    end else if(T27) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R41 <= 2'h0;
    end else if(T29) begin
      R41 <= T40;
    end
  end
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [1:0] io_in_4_bits_p_type,
    input [1:0] io_in_4_bits_client_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [1:0] io_in_3_bits_p_type,
    input [1:0] io_in_3_bits_client_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_p_type,
    input [1:0] io_in_2_bits_client_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_p_type,
    input [1:0] io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_p_type,
    input [1:0] io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_p_type,
    output[1:0] io_out_bits_client_id,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T141;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T142;
  reg  locked;
  wire T143;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  reg [1:0] R22;
  wire[1:0] T144;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire[2:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[25:0] T41;
  wire[25:0] T42;
  wire[25:0] T43;
  wire T44;
  wire[25:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R22 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T141 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T142 = reset ? 3'h4 : lockIdx;
  assign T143 = reset ? 1'h0 : T18;
  assign T18 = T19 ? 1'h0 : locked;
  assign T19 = T23 & T20;
  assign T20 = T21 == 2'h0;
  assign T21 = R22 + 2'h1;
  assign T144 = reset ? 2'h0 : R22;
  assign T23 = io_out_ready & io_out_valid;
  assign io_out_bits_client_id = T24;
  assign T24 = T32 ? io_in_4_bits_client_id : T25;
  assign T25 = T31 ? T29 : T26;
  assign T26 = T27 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T27 = T28[1'h0:1'h0];
  assign T28 = chosen;
  assign T29 = T30 ? io_in_3_bits_client_id : io_in_2_bits_client_id;
  assign T30 = T28[1'h0:1'h0];
  assign T31 = T28[1'h1:1'h1];
  assign T32 = T28[2'h2:2'h2];
  assign io_out_bits_p_type = T33;
  assign T33 = T40 ? io_in_4_bits_p_type : T34;
  assign T34 = T39 ? T37 : T35;
  assign T35 = T36 ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign T36 = T28[1'h0:1'h0];
  assign T37 = T38 ? io_in_3_bits_p_type : io_in_2_bits_p_type;
  assign T38 = T28[1'h0:1'h0];
  assign T39 = T28[1'h1:1'h1];
  assign T40 = T28[2'h2:2'h2];
  assign io_out_bits_addr_block = T41;
  assign T41 = T48 ? io_in_4_bits_addr_block : T42;
  assign T42 = T47 ? T45 : T43;
  assign T43 = T44 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T44 = T28[1'h0:1'h0];
  assign T45 = T46 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T46 = T28[1'h0:1'h0];
  assign T47 = T28[1'h1:1'h1];
  assign T48 = T28[2'h2:2'h2];
  assign io_out_valid = T49;
  assign T49 = T56 ? io_in_4_valid : T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52 ? io_in_1_valid : io_in_0_valid;
  assign T52 = T28[1'h0:1'h0];
  assign T53 = T54 ? io_in_3_valid : io_in_2_valid;
  assign T54 = T28[1'h0:1'h0];
  assign T55 = T28[1'h1:1'h1];
  assign T56 = T28[2'h2:2'h2];
  assign io_in_0_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = locked ? T76 : T59;
  assign T59 = T75 | T60;
  assign T60 = T61 ^ 1'h1;
  assign T61 = T64 | T62;
  assign T62 = io_in_4_valid & T63;
  assign T63 = last_grant < 3'h4;
  assign T64 = T67 | T65;
  assign T65 = io_in_3_valid & T66;
  assign T66 = last_grant < 3'h3;
  assign T67 = T70 | T68;
  assign T68 = io_in_2_valid & T69;
  assign T69 = last_grant < 3'h2;
  assign T70 = T73 | T71;
  assign T71 = io_in_1_valid & T72;
  assign T72 = last_grant < 3'h1;
  assign T73 = io_in_0_valid & T74;
  assign T74 = last_grant < 3'h0;
  assign T75 = last_grant < 3'h0;
  assign T76 = lockIdx == 3'h0;
  assign io_in_1_ready = T77;
  assign T77 = T78 & io_out_ready;
  assign T78 = locked ? T89 : T79;
  assign T79 = T86 | T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T82 | io_in_0_valid;
  assign T82 = T83 | T62;
  assign T83 = T84 | T65;
  assign T84 = T85 | T68;
  assign T85 = T73 | T71;
  assign T86 = T88 & T87;
  assign T87 = last_grant < 3'h1;
  assign T88 = T73 ^ 1'h1;
  assign T89 = lockIdx == 3'h1;
  assign io_in_2_ready = T90;
  assign T90 = T91 & io_out_ready;
  assign T91 = locked ? T104 : T92;
  assign T92 = T100 | T93;
  assign T93 = T94 ^ 1'h1;
  assign T94 = T95 | io_in_1_valid;
  assign T95 = T96 | io_in_0_valid;
  assign T96 = T97 | T62;
  assign T97 = T98 | T65;
  assign T98 = T99 | T68;
  assign T99 = T73 | T71;
  assign T100 = T102 & T101;
  assign T101 = last_grant < 3'h2;
  assign T102 = T103 ^ 1'h1;
  assign T103 = T73 | T71;
  assign T104 = lockIdx == 3'h2;
  assign io_in_3_ready = T105;
  assign T105 = T106 & io_out_ready;
  assign T106 = locked ? T121 : T107;
  assign T107 = T116 | T108;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T110 | io_in_2_valid;
  assign T110 = T111 | io_in_1_valid;
  assign T111 = T112 | io_in_0_valid;
  assign T112 = T113 | T62;
  assign T113 = T114 | T65;
  assign T114 = T115 | T68;
  assign T115 = T73 | T71;
  assign T116 = T118 & T117;
  assign T117 = last_grant < 3'h3;
  assign T118 = T119 ^ 1'h1;
  assign T119 = T120 | T68;
  assign T120 = T73 | T71;
  assign T121 = lockIdx == 3'h3;
  assign io_in_4_ready = T122;
  assign T122 = T123 & io_out_ready;
  assign T123 = locked ? T140 : T124;
  assign T124 = T134 | T125;
  assign T125 = T126 ^ 1'h1;
  assign T126 = T127 | io_in_3_valid;
  assign T127 = T128 | io_in_2_valid;
  assign T128 = T129 | io_in_1_valid;
  assign T129 = T130 | io_in_0_valid;
  assign T130 = T131 | T62;
  assign T131 = T132 | T65;
  assign T132 = T133 | T68;
  assign T133 = T73 | T71;
  assign T134 = T136 & T135;
  assign T135 = last_grant < 3'h4;
  assign T136 = T137 ^ 1'h1;
  assign T137 = T138 | T65;
  assign T138 = T139 | T68;
  assign T139 = T73 | T71;
  assign T140 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T19) begin
      locked <= 1'h0;
    end
    if(reset) begin
      R22 <= 2'h0;
    end
  end
endmodule

module LockingRRArbiter_5(input clk, input reset,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [25:0] io_in_4_bits_addr_block,
    input [2:0] io_in_4_bits_client_xact_id,
    input [1:0] io_in_4_bits_addr_beat,
    input  io_in_4_bits_is_builtin_type,
    input [2:0] io_in_4_bits_a_type,
    input [16:0] io_in_4_bits_union,
    input [3:0] io_in_4_bits_data,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [25:0] io_in_3_bits_addr_block,
    input [2:0] io_in_3_bits_client_xact_id,
    input [1:0] io_in_3_bits_addr_beat,
    input  io_in_3_bits_is_builtin_type,
    input [2:0] io_in_3_bits_a_type,
    input [16:0] io_in_3_bits_union,
    input [3:0] io_in_3_bits_data,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [2:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [3:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [2:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [3:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [2:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [3:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[2:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[3:0] io_out_bits_data,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] T0;
  wire[2:0] choose;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  reg [2:0] last_grant;
  wire[2:0] T189;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [2:0] lockIdx;
  wire[2:0] T190;
  wire[2:0] T18;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  locked;
  wire T191;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  reg [1:0] R38;
  wire[1:0] T192;
  wire[1:0] T39;
  wire[3:0] T40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire T43;
  wire[2:0] T44;
  wire[3:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire[16:0] T49;
  wire[16:0] T50;
  wire[16:0] T51;
  wire T52;
  wire[16:0] T53;
  wire T54;
  wire T55;
  wire T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire[2:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[2:0] T81;
  wire[2:0] T82;
  wire[2:0] T83;
  wire T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[25:0] T89;
  wire[25:0] T90;
  wire[25:0] T91;
  wire T92;
  wire[25:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R38 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T16 ? 3'h1 : T1;
  assign T1 = T14 ? 3'h2 : T2;
  assign T2 = T12 ? 3'h3 : T3;
  assign T3 = T8 ? 3'h4 : T4;
  assign T4 = io_in_0_valid ? 3'h0 : T5;
  assign T5 = io_in_1_valid ? 3'h1 : T6;
  assign T6 = io_in_2_valid ? 3'h2 : T7;
  assign T7 = io_in_3_valid ? 3'h3 : 3'h4;
  assign T8 = io_in_4_valid & T9;
  assign T9 = last_grant < 3'h4;
  assign T189 = reset ? 3'h0 : T10;
  assign T10 = T11 ? chosen : last_grant;
  assign T11 = io_out_ready & io_out_valid;
  assign T12 = io_in_3_valid & T13;
  assign T13 = last_grant < 3'h3;
  assign T14 = io_in_2_valid & T15;
  assign T15 = last_grant < 3'h2;
  assign T16 = io_in_1_valid & T17;
  assign T17 = last_grant < 3'h1;
  assign T190 = reset ? 3'h4 : T18;
  assign T18 = T27 ? T19 : lockIdx;
  assign T19 = T26 ? 3'h0 : T20;
  assign T20 = T25 ? 3'h1 : T21;
  assign T21 = T24 ? 3'h2 : T22;
  assign T22 = T23 ? 3'h3 : 3'h4;
  assign T23 = io_in_3_ready & io_in_3_valid;
  assign T24 = io_in_2_ready & io_in_2_valid;
  assign T25 = io_in_1_ready & io_in_1_valid;
  assign T26 = io_in_0_ready & io_in_0_valid;
  assign T27 = T29 & T28;
  assign T28 = locked ^ 1'h1;
  assign T29 = T32 & T30;
  assign T30 = io_out_bits_is_builtin_type & T31;
  assign T31 = 3'h3 == io_out_bits_a_type;
  assign T32 = io_out_ready & io_out_valid;
  assign T191 = reset ? 1'h0 : T33;
  assign T33 = T35 ? 1'h0 : T34;
  assign T34 = T27 ? 1'h1 : locked;
  assign T35 = T32 & T36;
  assign T36 = T37 == 2'h0;
  assign T37 = R38 + 2'h1;
  assign T192 = reset ? 2'h0 : T39;
  assign T39 = T29 ? T37 : R38;
  assign io_out_bits_data = T40;
  assign T40 = T48 ? io_in_4_bits_data : T41;
  assign T41 = T47 ? T45 : T42;
  assign T42 = T43 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = chosen;
  assign T45 = T46 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T46 = T44[1'h0:1'h0];
  assign T47 = T44[1'h1:1'h1];
  assign T48 = T44[2'h2:2'h2];
  assign io_out_bits_union = T49;
  assign T49 = T56 ? io_in_4_bits_union : T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T52 = T44[1'h0:1'h0];
  assign T53 = T54 ? io_in_3_bits_union : io_in_2_bits_union;
  assign T54 = T44[1'h0:1'h0];
  assign T55 = T44[1'h1:1'h1];
  assign T56 = T44[2'h2:2'h2];
  assign io_out_bits_a_type = T57;
  assign T57 = T64 ? io_in_4_bits_a_type : T58;
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T60 = T44[1'h0:1'h0];
  assign T61 = T62 ? io_in_3_bits_a_type : io_in_2_bits_a_type;
  assign T62 = T44[1'h0:1'h0];
  assign T63 = T44[1'h1:1'h1];
  assign T64 = T44[2'h2:2'h2];
  assign io_out_bits_is_builtin_type = T65;
  assign T65 = T72 ? io_in_4_bits_is_builtin_type : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T68 = T44[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_is_builtin_type : io_in_2_bits_is_builtin_type;
  assign T70 = T44[1'h0:1'h0];
  assign T71 = T44[1'h1:1'h1];
  assign T72 = T44[2'h2:2'h2];
  assign io_out_bits_addr_beat = T73;
  assign T73 = T80 ? io_in_4_bits_addr_beat : T74;
  assign T74 = T79 ? T77 : T75;
  assign T75 = T76 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T76 = T44[1'h0:1'h0];
  assign T77 = T78 ? io_in_3_bits_addr_beat : io_in_2_bits_addr_beat;
  assign T78 = T44[1'h0:1'h0];
  assign T79 = T44[1'h1:1'h1];
  assign T80 = T44[2'h2:2'h2];
  assign io_out_bits_client_xact_id = T81;
  assign T81 = T88 ? io_in_4_bits_client_xact_id : T82;
  assign T82 = T87 ? T85 : T83;
  assign T83 = T84 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T84 = T44[1'h0:1'h0];
  assign T85 = T86 ? io_in_3_bits_client_xact_id : io_in_2_bits_client_xact_id;
  assign T86 = T44[1'h0:1'h0];
  assign T87 = T44[1'h1:1'h1];
  assign T88 = T44[2'h2:2'h2];
  assign io_out_bits_addr_block = T89;
  assign T89 = T96 ? io_in_4_bits_addr_block : T90;
  assign T90 = T95 ? T93 : T91;
  assign T91 = T92 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T92 = T44[1'h0:1'h0];
  assign T93 = T94 ? io_in_3_bits_addr_block : io_in_2_bits_addr_block;
  assign T94 = T44[1'h0:1'h0];
  assign T95 = T44[1'h1:1'h1];
  assign T96 = T44[2'h2:2'h2];
  assign io_out_valid = T97;
  assign T97 = T104 ? io_in_4_valid : T98;
  assign T98 = T103 ? T101 : T99;
  assign T99 = T100 ? io_in_1_valid : io_in_0_valid;
  assign T100 = T44[1'h0:1'h0];
  assign T101 = T102 ? io_in_3_valid : io_in_2_valid;
  assign T102 = T44[1'h0:1'h0];
  assign T103 = T44[1'h1:1'h1];
  assign T104 = T44[2'h2:2'h2];
  assign io_in_0_ready = T105;
  assign T105 = T106 & io_out_ready;
  assign T106 = locked ? T124 : T107;
  assign T107 = T123 | T108;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T112 | T110;
  assign T110 = io_in_4_valid & T111;
  assign T111 = last_grant < 3'h4;
  assign T112 = T115 | T113;
  assign T113 = io_in_3_valid & T114;
  assign T114 = last_grant < 3'h3;
  assign T115 = T118 | T116;
  assign T116 = io_in_2_valid & T117;
  assign T117 = last_grant < 3'h2;
  assign T118 = T121 | T119;
  assign T119 = io_in_1_valid & T120;
  assign T120 = last_grant < 3'h1;
  assign T121 = io_in_0_valid & T122;
  assign T122 = last_grant < 3'h0;
  assign T123 = last_grant < 3'h0;
  assign T124 = lockIdx == 3'h0;
  assign io_in_1_ready = T125;
  assign T125 = T126 & io_out_ready;
  assign T126 = locked ? T137 : T127;
  assign T127 = T134 | T128;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | io_in_0_valid;
  assign T130 = T131 | T110;
  assign T131 = T132 | T113;
  assign T132 = T133 | T116;
  assign T133 = T121 | T119;
  assign T134 = T136 & T135;
  assign T135 = last_grant < 3'h1;
  assign T136 = T121 ^ 1'h1;
  assign T137 = lockIdx == 3'h1;
  assign io_in_2_ready = T138;
  assign T138 = T139 & io_out_ready;
  assign T139 = locked ? T152 : T140;
  assign T140 = T148 | T141;
  assign T141 = T142 ^ 1'h1;
  assign T142 = T143 | io_in_1_valid;
  assign T143 = T144 | io_in_0_valid;
  assign T144 = T145 | T110;
  assign T145 = T146 | T113;
  assign T146 = T147 | T116;
  assign T147 = T121 | T119;
  assign T148 = T150 & T149;
  assign T149 = last_grant < 3'h2;
  assign T150 = T151 ^ 1'h1;
  assign T151 = T121 | T119;
  assign T152 = lockIdx == 3'h2;
  assign io_in_3_ready = T153;
  assign T153 = T154 & io_out_ready;
  assign T154 = locked ? T169 : T155;
  assign T155 = T164 | T156;
  assign T156 = T157 ^ 1'h1;
  assign T157 = T158 | io_in_2_valid;
  assign T158 = T159 | io_in_1_valid;
  assign T159 = T160 | io_in_0_valid;
  assign T160 = T161 | T110;
  assign T161 = T162 | T113;
  assign T162 = T163 | T116;
  assign T163 = T121 | T119;
  assign T164 = T166 & T165;
  assign T165 = last_grant < 3'h3;
  assign T166 = T167 ^ 1'h1;
  assign T167 = T168 | T116;
  assign T168 = T121 | T119;
  assign T169 = lockIdx == 3'h3;
  assign io_in_4_ready = T170;
  assign T170 = T171 & io_out_ready;
  assign T171 = locked ? T188 : T172;
  assign T172 = T182 | T173;
  assign T173 = T174 ^ 1'h1;
  assign T174 = T175 | io_in_3_valid;
  assign T175 = T176 | io_in_2_valid;
  assign T176 = T177 | io_in_1_valid;
  assign T177 = T178 | io_in_0_valid;
  assign T178 = T179 | T110;
  assign T179 = T180 | T113;
  assign T180 = T181 | T116;
  assign T181 = T121 | T119;
  assign T182 = T184 & T183;
  assign T183 = last_grant < 3'h4;
  assign T184 = T185 ^ 1'h1;
  assign T185 = T186 | T113;
  assign T186 = T187 | T116;
  assign T187 = T121 | T119;
  assign T188 = lockIdx == 3'h4;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 3'h0;
    end else if(T11) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 3'h4;
    end else if(T27) begin
      lockIdx <= T19;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T35) begin
      locked <= 1'h0;
    end else if(T27) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R38 <= 2'h0;
    end else if(T29) begin
      R38 <= T37;
    end
  end
endmodule

module ClientUncachedTileLinkIOArbiter(input clk, input reset,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [25:0] io_in_4_acquire_bits_addr_block,
    input [2:0] io_in_4_acquire_bits_client_xact_id,
    input [1:0] io_in_4_acquire_bits_addr_beat,
    input  io_in_4_acquire_bits_is_builtin_type,
    input [2:0] io_in_4_acquire_bits_a_type,
    input [16:0] io_in_4_acquire_bits_union,
    input [3:0] io_in_4_acquire_bits_data,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_addr_beat,
    output[2:0] io_in_4_grant_bits_client_xact_id,
    output io_in_4_grant_bits_manager_xact_id,
    output io_in_4_grant_bits_is_builtin_type,
    output[3:0] io_in_4_grant_bits_g_type,
    output[3:0] io_in_4_grant_bits_data,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [25:0] io_in_3_acquire_bits_addr_block,
    input [2:0] io_in_3_acquire_bits_client_xact_id,
    input [1:0] io_in_3_acquire_bits_addr_beat,
    input  io_in_3_acquire_bits_is_builtin_type,
    input [2:0] io_in_3_acquire_bits_a_type,
    input [16:0] io_in_3_acquire_bits_union,
    input [3:0] io_in_3_acquire_bits_data,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_addr_beat,
    output[2:0] io_in_3_grant_bits_client_xact_id,
    output io_in_3_grant_bits_manager_xact_id,
    output io_in_3_grant_bits_is_builtin_type,
    output[3:0] io_in_3_grant_bits_g_type,
    output[3:0] io_in_3_grant_bits_data,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [25:0] io_in_2_acquire_bits_addr_block,
    input [2:0] io_in_2_acquire_bits_client_xact_id,
    input [1:0] io_in_2_acquire_bits_addr_beat,
    input  io_in_2_acquire_bits_is_builtin_type,
    input [2:0] io_in_2_acquire_bits_a_type,
    input [16:0] io_in_2_acquire_bits_union,
    input [3:0] io_in_2_acquire_bits_data,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_addr_beat,
    output[2:0] io_in_2_grant_bits_client_xact_id,
    output io_in_2_grant_bits_manager_xact_id,
    output io_in_2_grant_bits_is_builtin_type,
    output[3:0] io_in_2_grant_bits_g_type,
    output[3:0] io_in_2_grant_bits_data,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [25:0] io_in_1_acquire_bits_addr_block,
    input [2:0] io_in_1_acquire_bits_client_xact_id,
    input [1:0] io_in_1_acquire_bits_addr_beat,
    input  io_in_1_acquire_bits_is_builtin_type,
    input [2:0] io_in_1_acquire_bits_a_type,
    input [16:0] io_in_1_acquire_bits_union,
    input [3:0] io_in_1_acquire_bits_data,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_addr_beat,
    output[2:0] io_in_1_grant_bits_client_xact_id,
    output io_in_1_grant_bits_manager_xact_id,
    output io_in_1_grant_bits_is_builtin_type,
    output[3:0] io_in_1_grant_bits_g_type,
    output[3:0] io_in_1_grant_bits_data,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [25:0] io_in_0_acquire_bits_addr_block,
    input [2:0] io_in_0_acquire_bits_client_xact_id,
    input [1:0] io_in_0_acquire_bits_addr_beat,
    input  io_in_0_acquire_bits_is_builtin_type,
    input [2:0] io_in_0_acquire_bits_a_type,
    input [16:0] io_in_0_acquire_bits_union,
    input [3:0] io_in_0_acquire_bits_data,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_addr_beat,
    output[2:0] io_in_0_grant_bits_client_xact_id,
    output io_in_0_grant_bits_manager_xact_id,
    output io_in_0_grant_bits_is_builtin_type,
    output[3:0] io_in_0_grant_bits_g_type,
    output[3:0] io_in_0_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[3:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [3:0] io_out_grant_bits_data
);

  wire[2:0] T30;
  wire[5:0] T0;
  wire[2:0] T31;
  wire[5:0] T1;
  wire[2:0] T32;
  wire[5:0] T2;
  wire[2:0] T33;
  wire[5:0] T3;
  wire[2:0] T34;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire T21;
  wire T23;
  wire T25;
  wire T27;
  wire T29;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[25:0] LockingRRArbiter_io_out_bits_addr_block;
  wire[2:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[1:0] LockingRRArbiter_io_out_bits_addr_beat;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[2:0] LockingRRArbiter_io_out_bits_a_type;
  wire[16:0] LockingRRArbiter_io_out_bits_union;
  wire[3:0] LockingRRArbiter_io_out_bits_data;


  assign T30 = T0[2'h2:1'h0];
  assign T0 = {io_in_0_acquire_bits_client_xact_id, 3'h0};
  assign T31 = T1[2'h2:1'h0];
  assign T1 = {io_in_1_acquire_bits_client_xact_id, 3'h1};
  assign T32 = T2[2'h2:1'h0];
  assign T2 = {io_in_2_acquire_bits_client_xact_id, 3'h2};
  assign T33 = T3[2'h2:1'h0];
  assign T3 = {io_in_3_acquire_bits_client_xact_id, 3'h3};
  assign T34 = T4[2'h2:1'h0];
  assign T4 = {io_in_4_acquire_bits_client_xact_id, 3'h4};
  assign io_out_grant_ready = T5;
  assign T5 = T18 ? io_in_4_grant_ready : T6;
  assign T6 = T16 ? io_in_3_grant_ready : T7;
  assign T7 = T14 ? io_in_2_grant_ready : T8;
  assign T8 = T12 ? io_in_1_grant_ready : T9;
  assign T9 = T10 ? io_in_0_grant_ready : 1'h0;
  assign T10 = T11 == 3'h0;
  assign T11 = io_out_grant_bits_client_xact_id;
  assign T12 = T13 == 3'h1;
  assign T13 = io_out_grant_bits_client_xact_id;
  assign T14 = T15 == 3'h2;
  assign T15 = io_out_grant_bits_client_xact_id;
  assign T16 = T17 == 3'h3;
  assign T17 = io_out_grant_bits_client_xact_id;
  assign T18 = T19 == 3'h4;
  assign T19 = io_out_grant_bits_client_xact_id;
  assign io_out_acquire_bits_data = LockingRRArbiter_io_out_bits_data;
  assign io_out_acquire_bits_union = LockingRRArbiter_io_out_bits_union;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_io_out_bits_addr_block;
  assign io_out_acquire_valid = LockingRRArbiter_io_out_valid;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_client_xact_id = 3'h0;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_valid = T21;
  assign T21 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = LockingRRArbiter_io_in_0_ready;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_client_xact_id = 3'h0;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_valid = T23;
  assign T23 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = LockingRRArbiter_io_in_1_ready;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_client_xact_id = 3'h0;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_valid = T25;
  assign T25 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = LockingRRArbiter_io_in_2_ready;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_client_xact_id = 3'h0;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_valid = T27;
  assign T27 = T16 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = LockingRRArbiter_io_in_3_ready;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_client_xact_id = 3'h0;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_valid = T29;
  assign T29 = T18 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = LockingRRArbiter_io_in_4_ready;
  LockingRRArbiter_5 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_addr_block( io_in_4_acquire_bits_addr_block ),
       .io_in_4_bits_client_xact_id( T34 ),
       .io_in_4_bits_addr_beat( io_in_4_acquire_bits_addr_beat ),
       .io_in_4_bits_is_builtin_type( io_in_4_acquire_bits_is_builtin_type ),
       .io_in_4_bits_a_type( io_in_4_acquire_bits_a_type ),
       .io_in_4_bits_union( io_in_4_acquire_bits_union ),
       .io_in_4_bits_data( io_in_4_acquire_bits_data ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_addr_block( io_in_3_acquire_bits_addr_block ),
       .io_in_3_bits_client_xact_id( T33 ),
       .io_in_3_bits_addr_beat( io_in_3_acquire_bits_addr_beat ),
       .io_in_3_bits_is_builtin_type( io_in_3_acquire_bits_is_builtin_type ),
       .io_in_3_bits_a_type( io_in_3_acquire_bits_a_type ),
       .io_in_3_bits_union( io_in_3_acquire_bits_union ),
       .io_in_3_bits_data( io_in_3_acquire_bits_data ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_addr_block( io_in_2_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( T32 ),
       .io_in_2_bits_addr_beat( io_in_2_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( io_in_2_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( io_in_2_acquire_bits_a_type ),
       .io_in_2_bits_union( io_in_2_acquire_bits_union ),
       .io_in_2_bits_data( io_in_2_acquire_bits_data ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_addr_block( io_in_1_acquire_bits_addr_block ),
       .io_in_1_bits_client_xact_id( T31 ),
       .io_in_1_bits_addr_beat( io_in_1_acquire_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( io_in_1_acquire_bits_is_builtin_type ),
       .io_in_1_bits_a_type( io_in_1_acquire_bits_a_type ),
       .io_in_1_bits_union( io_in_1_acquire_bits_union ),
       .io_in_1_bits_data( io_in_1_acquire_bits_data ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_addr_block( io_in_0_acquire_bits_addr_block ),
       .io_in_0_bits_client_xact_id( T30 ),
       .io_in_0_bits_addr_beat( io_in_0_acquire_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( io_in_0_acquire_bits_is_builtin_type ),
       .io_in_0_bits_a_type( io_in_0_acquire_bits_a_type ),
       .io_in_0_bits_union( io_in_0_acquire_bits_union ),
       .io_in_0_bits_data( io_in_0_acquire_bits_data ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( LockingRRArbiter_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( LockingRRArbiter_io_out_bits_a_type ),
       .io_out_bits_union( LockingRRArbiter_io_out_bits_union ),
       .io_out_bits_data( LockingRRArbiter_io_out_bits_data )
       //.io_chosen(  )
  );
endmodule

module L2BroadcastHub(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [1:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input [1:0] io_inner_acquire_bits_client_id,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[1:0] io_inner_grant_bits_client_xact_id,
    output[2:0] io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    output[1:0] io_inner_grant_bits_client_id,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [2:0] io_inner_finish_bits_manager_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output[1:0] io_inner_probe_bits_client_id,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [1:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [127:0] io_inner_release_bits_data,
    input [1:0] io_inner_release_bits_client_id,
    input  io_incoherent_0,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[4:0] releaseMatches;
  wire[4:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[3:0] T224;
  wire[127:0] T225;
  wire[127:0] T226;
  wire[127:0] T227;
  wire[127:0] T228;
  wire[127:0] T229;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  reg [1:0] rel_data_cnt;
  wire[1:0] T230;
  wire[1:0] T14;
  wire[1:0] T15;
  wire vwbdq_enq;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T231;
  wire[2:0] T232;
  wire[2:0] T233;
  wire[2:0] T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  wire[1:0] T239;
  wire[1:0] T240;
  wire[1:0] T241;
  wire T242;
  wire[3:0] T31;
  reg [3:0] sdq_val;
  wire[3:0] T243;
  wire[3:0] T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[3:0] T244;
  wire sdq_enq;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[3:0] T56;
  wire[3:0] T245;
  wire free_sdq;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[3:0] T67;
  wire[1:0] T68;
  wire T69;
  wire T246;
  wire T247;
  wire T70;
  wire T71;
  wire[2:0] acquire_idx;
  wire[2:0] T248;
  wire[2:0] T249;
  wire[2:0] T250;
  wire[2:0] T251;
  wire T252;
  wire[4:0] acquireReadys;
  wire[4:0] T73;
  wire[2:0] T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire T253;
  wire T254;
  wire T255;
  wire[2:0] T256;
  wire[2:0] T257;
  wire[2:0] T258;
  wire[2:0] T259;
  wire T260;
  wire[4:0] acquireMatches;
  wire[4:0] T78;
  wire[2:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T261;
  wire T262;
  wire T263;
  wire T82;
  wire T83;
  wire T84;
  wire block_acquires;
  wire T85;
  wire sdq_rdy;
  wire T86;
  wire T87;
  wire[4:0] acquireConflicts;
  wire[4:0] T88;
  wire[2:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[3:0] T92;
  wire[3:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[3:0] T100;
  wire[3:0] T101;
  wire[1:0] T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[3:0] T116;
  wire[3:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire[3:0] T132;
  wire[3:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[3:0] T140;
  wire[3:0] T141;
  wire[1:0] T142;
  wire[1:0] T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire[3:0] T148;
  wire[3:0] T149;
  wire[1:0] T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire[127:0] T156;
  wire[127:0] T157;
  wire[127:0] T158;
  wire[127:0] T159;
  reg [127:0] vwbdq_0;
  wire[127:0] T160;
  wire T161;
  wire T162;
  wire[3:0] T163;
  wire[1:0] T164;
  reg [127:0] vwbdq_1;
  wire[127:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] T169;
  wire[127:0] T170;
  reg [127:0] vwbdq_2;
  wire[127:0] T171;
  wire T172;
  wire T173;
  reg [127:0] vwbdq_3;
  wire[127:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire[127:0] T180;
  wire[127:0] T181;
  reg [127:0] sdq_0;
  wire[127:0] T182;
  wire T183;
  wire T184;
  wire[3:0] T185;
  wire[1:0] T186;
  reg [127:0] sdq_1;
  wire[127:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire[1:0] T191;
  wire[127:0] T192;
  reg [127:0] sdq_2;
  wire[127:0] T193;
  wire T194;
  wire T195;
  reg [127:0] sdq_3;
  wire[127:0] T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[2:0] T205;
  wire[2:0] T206;
  wire T207;
  wire[4:0] releaseReadys;
  wire[4:0] T208;
  wire[2:0] T209;
  wire[1:0] T210;
  wire[1:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[2:0] T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_valid;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id;
  wire BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  wire BroadcastVoluntaryReleaseTracker_io_inner_probe_valid;
  wire BroadcastVoluntaryReleaseTracker_io_inner_release_ready;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data;
  wire BroadcastVoluntaryReleaseTracker_io_outer_grant_ready;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict;
  wire BroadcastVoluntaryReleaseTracker_io_has_acquire_match;
  wire BroadcastVoluntaryReleaseTracker_io_has_release_match;
  wire BroadcastAcquireTracker_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_finish_ready;
  wire BroadcastAcquireTracker_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_io_inner_release_ready;
  wire BroadcastAcquireTracker_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_io_outer_grant_ready;
  wire BroadcastAcquireTracker_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_io_has_acquire_match;
  wire BroadcastAcquireTracker_io_has_release_match;
  wire BroadcastAcquireTracker_1_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_1_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_1_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_finish_ready;
  wire BroadcastAcquireTracker_1_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_1_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_1_io_inner_release_ready;
  wire BroadcastAcquireTracker_1_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_1_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_1_io_outer_grant_ready;
  wire BroadcastAcquireTracker_1_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_1_io_has_acquire_match;
  wire BroadcastAcquireTracker_1_io_has_release_match;
  wire BroadcastAcquireTracker_2_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_2_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_2_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_finish_ready;
  wire BroadcastAcquireTracker_2_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_2_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_2_io_inner_release_ready;
  wire BroadcastAcquireTracker_2_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_2_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_2_io_outer_grant_ready;
  wire BroadcastAcquireTracker_2_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_2_io_has_acquire_match;
  wire BroadcastAcquireTracker_2_io_has_release_match;
  wire BroadcastAcquireTracker_3_io_inner_acquire_ready;
  wire BroadcastAcquireTracker_3_io_inner_grant_valid;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id;
  wire[2:0] BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id;
  wire BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_g_type;
  wire[3:0] BroadcastAcquireTracker_3_io_inner_grant_bits_data;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_grant_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_finish_ready;
  wire BroadcastAcquireTracker_3_io_inner_probe_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_p_type;
  wire[1:0] BroadcastAcquireTracker_3_io_inner_probe_bits_client_id;
  wire BroadcastAcquireTracker_3_io_inner_release_ready;
  wire BroadcastAcquireTracker_3_io_outer_acquire_valid;
  wire[25:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id;
  wire[1:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat;
  wire BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type;
  wire[16:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_union;
  wire[3:0] BroadcastAcquireTracker_3_io_outer_acquire_bits_data;
  wire BroadcastAcquireTracker_3_io_outer_grant_ready;
  wire BroadcastAcquireTracker_3_io_has_acquire_conflict;
  wire BroadcastAcquireTracker_3_io_has_acquire_match;
  wire BroadcastAcquireTracker_3_io_has_release_match;
  wire LockingRRArbiter_io_in_4_ready;
  wire LockingRRArbiter_io_in_3_ready;
  wire LockingRRArbiter_io_in_2_ready;
  wire LockingRRArbiter_io_in_1_ready;
  wire LockingRRArbiter_io_in_0_ready;
  wire LockingRRArbiter_io_out_valid;
  wire[1:0] LockingRRArbiter_io_out_bits_client_xact_id;
  wire[2:0] LockingRRArbiter_io_out_bits_manager_xact_id;
  wire LockingRRArbiter_io_out_bits_is_builtin_type;
  wire[3:0] LockingRRArbiter_io_out_bits_g_type;
  wire[1:0] LockingRRArbiter_io_out_bits_client_id;
  wire LockingRRArbiter_1_io_in_4_ready;
  wire LockingRRArbiter_1_io_in_3_ready;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire LockingRRArbiter_1_io_out_valid;
  wire[25:0] LockingRRArbiter_1_io_out_bits_addr_block;
  wire[1:0] LockingRRArbiter_1_io_out_bits_p_type;
  wire[1:0] LockingRRArbiter_1_io_out_bits_client_id;
  wire outer_arb_io_in_4_acquire_ready;
  wire outer_arb_io_in_4_grant_valid;
  wire[1:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire[2:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_4_grant_bits_data;
  wire outer_arb_io_in_3_acquire_ready;
  wire outer_arb_io_in_3_grant_valid;
  wire[1:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire[2:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_3_grant_bits_data;
  wire outer_arb_io_in_2_acquire_ready;
  wire outer_arb_io_in_2_grant_valid;
  wire[1:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire[2:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_2_grant_bits_data;
  wire outer_arb_io_in_1_acquire_ready;
  wire outer_arb_io_in_1_grant_valid;
  wire[1:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire[2:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_1_grant_bits_data;
  wire outer_arb_io_in_0_acquire_ready;
  wire outer_arb_io_in_0_grant_valid;
  wire[1:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire[2:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire[3:0] outer_arb_io_in_0_grant_bits_data;
  wire outer_arb_io_out_acquire_valid;
  wire[25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire[2:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire[1:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire outer_arb_io_out_acquire_bits_is_builtin_type;
  wire[2:0] outer_arb_io_out_acquire_bits_a_type;
  wire[16:0] outer_arb_io_out_acquire_bits_union;
  wire[3:0] outer_arb_io_out_acquire_bits_data;
  wire outer_arb_io_out_grant_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    rel_data_cnt = {1{$random}};
    sdq_val = {1{$random}};
    vwbdq_0 = {4{$random}};
    vwbdq_1 = {4{$random}};
    vwbdq_2 = {4{$random}};
    vwbdq_3 = {4{$random}};
    sdq_0 = {4{$random}};
    sdq_1 = {4{$random}};
    sdq_2 = {4{$random}};
    sdq_3 = {4{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_inner_release_valid & T4;
  assign T4 = T5 ^ 1'h1;
  assign T5 = releaseMatches != 5'h0;
  assign releaseMatches = T6;
  assign T6 = {T9, T7};
  assign T7 = {BroadcastAcquireTracker_1_io_has_release_match, T8};
  assign T8 = {BroadcastAcquireTracker_io_has_release_match, BroadcastVoluntaryReleaseTracker_io_has_release_match};
  assign T9 = {BroadcastAcquireTracker_3_io_has_release_match, BroadcastAcquireTracker_2_io_has_release_match};
  assign T224 = io_outer_grant_bits_data[2'h3:1'h0];
  assign T225 = {124'h0, BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data};
  assign T226 = {124'h0, BroadcastAcquireTracker_io_inner_grant_bits_data};
  assign T227 = {124'h0, BroadcastAcquireTracker_1_io_inner_grant_bits_data};
  assign T228 = {124'h0, BroadcastAcquireTracker_2_io_inner_grant_bits_data};
  assign T229 = {124'h0, BroadcastAcquireTracker_3_io_inner_grant_bits_data};
  assign T10 = T11;
  assign T11 = {T13, T12};
  assign T12 = 2'h2;
  assign T13 = rel_data_cnt;
  assign T230 = reset ? 2'h0 : T14;
  assign T14 = vwbdq_enq ? T15 : rel_data_cnt;
  assign T15 = rel_data_cnt + 2'h1;
  assign vwbdq_enq = T21 & T16;
  assign T16 = T18 | T17;
  assign T17 = 3'h2 == io_inner_release_bits_r_type;
  assign T18 = T20 | T19;
  assign T19 = 3'h1 == io_inner_release_bits_r_type;
  assign T20 = 3'h0 == io_inner_release_bits_r_type;
  assign T21 = T22 & io_inner_release_bits_voluntary;
  assign T22 = io_inner_release_ready & io_inner_release_valid;
  assign T23 = io_inner_release_valid & T24;
  assign T24 = T231 == 3'h4;
  assign T231 = T238 ? 1'h0 : T232;
  assign T232 = T237 ? 1'h1 : T233;
  assign T233 = T236 ? 2'h2 : T234;
  assign T234 = T235 ? 2'h3 : 3'h4;
  assign T235 = releaseMatches[2'h3:2'h3];
  assign T236 = releaseMatches[2'h2:2'h2];
  assign T237 = releaseMatches[1'h1:1'h1];
  assign T238 = releaseMatches[1'h0:1'h0];
  assign T25 = io_inner_finish_valid & T26;
  assign T26 = io_inner_finish_bits_manager_xact_id == 3'h4;
  assign T27 = T28;
  assign T28 = {T30, T29};
  assign T29 = 2'h0;
  assign T30 = T239;
  assign T239 = T247 ? 1'h0 : T240;
  assign T240 = T246 ? 1'h1 : T241;
  assign T241 = T242 ? 2'h2 : 2'h3;
  assign T242 = T31[2'h2:2'h2];
  assign T31 = ~ sdq_val;
  assign T243 = reset ? 4'h0 : T32;
  assign T32 = T69 ? T33 : sdq_val;
  assign T33 = T53 | T34;
  assign T34 = T43 & T35;
  assign T35 = 4'h0 - T244;
  assign T244 = {3'h0, sdq_enq};
  assign sdq_enq = T42 & T36;
  assign T36 = io_inner_acquire_bits_is_builtin_type & T37;
  assign T37 = T39 | T38;
  assign T38 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T39 = T41 | T40;
  assign T40 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T41 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T42 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T43 = T52 ? 4'h1 : T44;
  assign T44 = T51 ? 4'h2 : T45;
  assign T45 = T50 ? 4'h4 : T46;
  assign T46 = T47 ? 4'h8 : 4'h0;
  assign T47 = T48[2'h3:2'h3];
  assign T48 = ~ T49;
  assign T49 = sdq_val[2'h3:1'h0];
  assign T50 = T48[2'h2:2'h2];
  assign T51 = T48[1'h1:1'h1];
  assign T52 = T48[1'h0:1'h0];
  assign T53 = sdq_val & T54;
  assign T54 = ~ T55;
  assign T55 = T67 & T56;
  assign T56 = 4'h0 - T245;
  assign T245 = {3'h0, free_sdq};
  assign free_sdq = T59 & T57;
  assign T57 = T58 == 2'h0;
  assign T58 = outer_arb_io_out_acquire_bits_data[1'h1:1'h0];
  assign T59 = T66 & T60;
  assign T60 = io_outer_acquire_bits_is_builtin_type & T61;
  assign T61 = T63 | T62;
  assign T62 = 3'h4 == io_outer_acquire_bits_a_type;
  assign T63 = T65 | T64;
  assign T64 = 3'h3 == io_outer_acquire_bits_a_type;
  assign T65 = 3'h2 == io_outer_acquire_bits_a_type;
  assign T66 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T67 = 1'h1 << T68;
  assign T68 = outer_arb_io_out_acquire_bits_data[2'h3:2'h2];
  assign T69 = io_outer_acquire_valid | sdq_enq;
  assign T246 = T31[1'h1:1'h1];
  assign T247 = T31[1'h0:1'h0];
  assign T70 = T83 & T71;
  assign T71 = acquire_idx == 3'h4;
  assign acquire_idx = T82 ? T256 : T248;
  assign T248 = T255 ? 1'h0 : T249;
  assign T249 = T254 ? 1'h1 : T250;
  assign T250 = T253 ? 2'h2 : T251;
  assign T251 = T252 ? 2'h3 : 3'h4;
  assign T252 = acquireReadys[2'h3:2'h3];
  assign acquireReadys = T73;
  assign T73 = {T76, T74};
  assign T74 = {BroadcastAcquireTracker_1_io_inner_acquire_ready, T75};
  assign T75 = {BroadcastAcquireTracker_io_inner_acquire_ready, BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready};
  assign T76 = {BroadcastAcquireTracker_3_io_inner_acquire_ready, BroadcastAcquireTracker_2_io_inner_acquire_ready};
  assign T253 = acquireReadys[2'h2:2'h2];
  assign T254 = acquireReadys[1'h1:1'h1];
  assign T255 = acquireReadys[1'h0:1'h0];
  assign T256 = T263 ? 1'h0 : T257;
  assign T257 = T262 ? 1'h1 : T258;
  assign T258 = T261 ? 2'h2 : T259;
  assign T259 = T260 ? 2'h3 : 3'h4;
  assign T260 = acquireMatches[2'h3:2'h3];
  assign acquireMatches = T78;
  assign T78 = {T81, T79};
  assign T79 = {BroadcastAcquireTracker_1_io_has_acquire_match, T80};
  assign T80 = {BroadcastAcquireTracker_io_has_acquire_match, BroadcastVoluntaryReleaseTracker_io_has_acquire_match};
  assign T81 = {BroadcastAcquireTracker_3_io_has_acquire_match, BroadcastAcquireTracker_2_io_has_acquire_match};
  assign T261 = acquireMatches[2'h2:2'h2];
  assign T262 = acquireMatches[1'h1:1'h1];
  assign T263 = acquireMatches[1'h0:1'h0];
  assign T82 = acquireMatches != 5'h0;
  assign T83 = io_inner_acquire_valid & T84;
  assign T84 = block_acquires ^ 1'h1;
  assign block_acquires = T87 | T85;
  assign T85 = sdq_rdy ^ 1'h1;
  assign sdq_rdy = T86 ^ 1'h1;
  assign T86 = sdq_val == 4'hf;
  assign T87 = acquireConflicts != 5'h0;
  assign acquireConflicts = T88;
  assign T88 = {T91, T89};
  assign T89 = {BroadcastAcquireTracker_1_io_has_acquire_conflict, T90};
  assign T90 = {BroadcastAcquireTracker_io_has_acquire_conflict, BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict};
  assign T91 = {BroadcastAcquireTracker_3_io_has_acquire_conflict, BroadcastAcquireTracker_2_io_has_acquire_conflict};
  assign T92 = T93;
  assign T93 = {T95, T94};
  assign T94 = 2'h2;
  assign T95 = rel_data_cnt;
  assign T96 = io_inner_release_valid & T97;
  assign T97 = T231 == 3'h3;
  assign T98 = io_inner_finish_valid & T99;
  assign T99 = io_inner_finish_bits_manager_xact_id == 3'h3;
  assign T100 = T101;
  assign T101 = {T103, T102};
  assign T102 = 2'h0;
  assign T103 = T239;
  assign T104 = T106 & T105;
  assign T105 = acquire_idx == 3'h3;
  assign T106 = io_inner_acquire_valid & T107;
  assign T107 = block_acquires ^ 1'h1;
  assign T108 = T109;
  assign T109 = {T111, T110};
  assign T110 = 2'h2;
  assign T111 = rel_data_cnt;
  assign T112 = io_inner_release_valid & T113;
  assign T113 = T231 == 3'h2;
  assign T114 = io_inner_finish_valid & T115;
  assign T115 = io_inner_finish_bits_manager_xact_id == 3'h2;
  assign T116 = T117;
  assign T117 = {T119, T118};
  assign T118 = 2'h0;
  assign T119 = T239;
  assign T120 = T122 & T121;
  assign T121 = acquire_idx == 3'h2;
  assign T122 = io_inner_acquire_valid & T123;
  assign T123 = block_acquires ^ 1'h1;
  assign T124 = T125;
  assign T125 = {T127, T126};
  assign T126 = 2'h2;
  assign T127 = rel_data_cnt;
  assign T128 = io_inner_release_valid & T129;
  assign T129 = T231 == 3'h1;
  assign T130 = io_inner_finish_valid & T131;
  assign T131 = io_inner_finish_bits_manager_xact_id == 3'h1;
  assign T132 = T133;
  assign T133 = {T135, T134};
  assign T134 = 2'h0;
  assign T135 = T239;
  assign T136 = T138 & T137;
  assign T137 = acquire_idx == 3'h1;
  assign T138 = io_inner_acquire_valid & T139;
  assign T139 = block_acquires ^ 1'h1;
  assign T140 = T141;
  assign T141 = {T143, T142};
  assign T142 = 2'h1;
  assign T143 = rel_data_cnt;
  assign T144 = io_inner_release_valid & T145;
  assign T145 = T231 == 3'h0;
  assign T146 = io_inner_finish_valid & T147;
  assign T147 = io_inner_finish_bits_manager_xact_id == 3'h0;
  assign T148 = T149;
  assign T149 = {T151, T150};
  assign T150 = 2'h0;
  assign T151 = T239;
  assign T152 = T154 & T153;
  assign T153 = acquire_idx == 3'h0;
  assign T154 = io_inner_acquire_valid & T155;
  assign T155 = block_acquires ^ 1'h1;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_data = T156;
  assign T156 = T201 ? T180 : T157;
  assign T157 = T179 ? T158 : io_inner_release_bits_data;
  assign T158 = T178 ? T170 : T159;
  assign T159 = T168 ? vwbdq_1 : vwbdq_0;
  assign T160 = T161 ? io_inner_release_bits_data : vwbdq_0;
  assign T161 = vwbdq_enq & T162;
  assign T162 = T163[1'h0:1'h0];
  assign T163 = 1'h1 << T164;
  assign T164 = rel_data_cnt;
  assign T165 = T166 ? io_inner_release_bits_data : vwbdq_1;
  assign T166 = vwbdq_enq & T167;
  assign T167 = T163[1'h1:1'h1];
  assign T168 = T169[1'h0:1'h0];
  assign T169 = T68;
  assign T170 = T177 ? vwbdq_3 : vwbdq_2;
  assign T171 = T172 ? io_inner_release_bits_data : vwbdq_2;
  assign T172 = vwbdq_enq & T173;
  assign T173 = T163[2'h2:2'h2];
  assign T174 = T175 ? io_inner_release_bits_data : vwbdq_3;
  assign T175 = vwbdq_enq & T176;
  assign T176 = T163[2'h3:2'h3];
  assign T177 = T169[1'h0:1'h0];
  assign T178 = T169[1'h1:1'h1];
  assign T179 = T58 == 2'h1;
  assign T180 = T200 ? T192 : T181;
  assign T181 = T190 ? sdq_1 : sdq_0;
  assign T182 = T183 ? io_inner_acquire_bits_data : sdq_0;
  assign T183 = sdq_enq & T184;
  assign T184 = T185[1'h0:1'h0];
  assign T185 = 1'h1 << T186;
  assign T186 = T239;
  assign T187 = T188 ? io_inner_acquire_bits_data : sdq_1;
  assign T188 = sdq_enq & T189;
  assign T189 = T185[1'h1:1'h1];
  assign T190 = T191[1'h0:1'h0];
  assign T191 = T68;
  assign T192 = T199 ? sdq_3 : sdq_2;
  assign T193 = T194 ? io_inner_acquire_bits_data : sdq_2;
  assign T194 = sdq_enq & T195;
  assign T195 = T185[2'h2:2'h2];
  assign T196 = T197 ? io_inner_acquire_bits_data : sdq_3;
  assign T197 = sdq_enq & T198;
  assign T198 = T185[2'h3:2'h3];
  assign T199 = T191[1'h0:1'h0];
  assign T200 = T191[1'h1:1'h1];
  assign T201 = T58 == 2'h0;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T202;
  assign T202 = T207 & T203;
  assign T203 = T204 - 1'h1;
  assign T204 = 1'h1 << T205;
  assign T205 = T206 + 3'h1;
  assign T206 = T231 - T231;
  assign T207 = releaseReadys >> T231;
  assign releaseReadys = T208;
  assign T208 = {T211, T209};
  assign T209 = {BroadcastAcquireTracker_1_io_inner_release_ready, T210};
  assign T210 = {BroadcastAcquireTracker_io_inner_release_ready, BroadcastVoluntaryReleaseTracker_io_inner_release_ready};
  assign T211 = {BroadcastAcquireTracker_3_io_inner_release_ready, BroadcastAcquireTracker_2_io_inner_release_ready};
  assign io_inner_probe_bits_client_id = LockingRRArbiter_1_io_out_bits_client_id;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_1_io_out_bits_p_type;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_1_io_out_bits_addr_block;
  assign io_inner_probe_valid = LockingRRArbiter_1_io_out_valid;
  assign io_inner_finish_ready = T212;
  assign T212 = T220 ? BroadcastAcquireTracker_3_io_inner_finish_ready : T213;
  assign T213 = T219 ? T217 : T214;
  assign T214 = T215 ? BroadcastAcquireTracker_io_inner_finish_ready : BroadcastVoluntaryReleaseTracker_io_inner_finish_ready;
  assign T215 = T216[1'h0:1'h0];
  assign T216 = io_inner_finish_bits_manager_xact_id;
  assign T217 = T218 ? BroadcastAcquireTracker_2_io_inner_finish_ready : BroadcastAcquireTracker_1_io_inner_finish_ready;
  assign T218 = T216[1'h0:1'h0];
  assign T219 = T216[1'h1:1'h1];
  assign T220 = T216[2'h2:2'h2];
  assign io_inner_grant_bits_client_id = LockingRRArbiter_io_out_bits_client_id;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_io_out_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = LockingRRArbiter_io_out_valid;
  assign io_inner_acquire_ready = T221;
  assign T221 = T223 & T222;
  assign T222 = block_acquires ^ 1'h1;
  assign T223 = acquireReadys != 5'h0;
  BroadcastVoluntaryReleaseTracker BroadcastVoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastVoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T152 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T148 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_0_ready ),
       .io_inner_grant_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastVoluntaryReleaseTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T146 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_inner_probe_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_addr_block(  )
       //.io_inner_probe_bits_p_type(  )
       //.io_inner_probe_bits_client_id(  )
       .io_inner_release_ready( BroadcastVoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T144 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T140 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastVoluntaryReleaseTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastVoluntaryReleaseTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastVoluntaryReleaseTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_0 BroadcastAcquireTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T136 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T132 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_1_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_io_inner_finish_ready ),
       .io_inner_finish_valid( T130 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_io_inner_release_ready ),
       .io_inner_release_valid( T128 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T124 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_io_has_release_match )
  );
  BroadcastAcquireTracker_1 BroadcastAcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T120 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T116 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_2_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_1_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_1_io_inner_finish_ready ),
       .io_inner_finish_valid( T114 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T112 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T108 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_1_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_1_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_1_io_has_release_match )
  );
  BroadcastAcquireTracker_2 BroadcastAcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T104 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T100 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_3_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_2_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_2_io_inner_finish_ready ),
       .io_inner_finish_valid( T98 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T96 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T92 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_2_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_2_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_2_io_has_release_match )
  );
  BroadcastAcquireTracker_3 BroadcastAcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( BroadcastAcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( T70 ),
       .io_inner_acquire_bits_addr_block( io_inner_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( io_inner_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( io_inner_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( io_inner_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( io_inner_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( io_inner_acquire_bits_union ),
       .io_inner_acquire_bits_data( T27 ),
       .io_inner_acquire_bits_client_id( io_inner_acquire_bits_client_id ),
       .io_inner_grant_ready( LockingRRArbiter_io_in_4_ready ),
       .io_inner_grant_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( BroadcastAcquireTracker_3_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( BroadcastAcquireTracker_3_io_inner_finish_ready ),
       .io_inner_finish_valid( T25 ),
       .io_inner_finish_bits_manager_xact_id( io_inner_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_inner_probe_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( BroadcastAcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T23 ),
       .io_inner_release_bits_addr_beat( io_inner_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( io_inner_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( io_inner_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( io_inner_release_bits_voluntary ),
       .io_inner_release_bits_r_type( io_inner_release_bits_r_type ),
       .io_inner_release_bits_data( T10 ),
       .io_inner_release_bits_client_id( io_inner_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_outer_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_has_acquire_conflict( BroadcastAcquireTracker_3_io_has_acquire_conflict ),
       .io_has_acquire_match( BroadcastAcquireTracker_3_io_has_acquire_match ),
       .io_has_release_match( BroadcastAcquireTracker_3_io_has_release_match )
  );
  LockingRRArbiter_2 LockingRRArbiter(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_addr_beat( BroadcastAcquireTracker_3_io_inner_grant_bits_addr_beat ),
       .io_in_4_bits_client_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_xact_id ),
       .io_in_4_bits_manager_xact_id( BroadcastAcquireTracker_3_io_inner_grant_bits_manager_xact_id ),
       .io_in_4_bits_is_builtin_type( BroadcastAcquireTracker_3_io_inner_grant_bits_is_builtin_type ),
       .io_in_4_bits_g_type( BroadcastAcquireTracker_3_io_inner_grant_bits_g_type ),
       .io_in_4_bits_data( T229 ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_grant_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_addr_beat( BroadcastAcquireTracker_2_io_inner_grant_bits_addr_beat ),
       .io_in_3_bits_client_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_xact_id ),
       .io_in_3_bits_manager_xact_id( BroadcastAcquireTracker_2_io_inner_grant_bits_manager_xact_id ),
       .io_in_3_bits_is_builtin_type( BroadcastAcquireTracker_2_io_inner_grant_bits_is_builtin_type ),
       .io_in_3_bits_g_type( BroadcastAcquireTracker_2_io_inner_grant_bits_g_type ),
       .io_in_3_bits_data( T228 ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_grant_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_addr_beat( BroadcastAcquireTracker_1_io_inner_grant_bits_addr_beat ),
       .io_in_2_bits_client_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_xact_id ),
       .io_in_2_bits_manager_xact_id( BroadcastAcquireTracker_1_io_inner_grant_bits_manager_xact_id ),
       .io_in_2_bits_is_builtin_type( BroadcastAcquireTracker_1_io_inner_grant_bits_is_builtin_type ),
       .io_in_2_bits_g_type( BroadcastAcquireTracker_1_io_inner_grant_bits_g_type ),
       .io_in_2_bits_data( T227 ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_grant_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_grant_valid ),
       .io_in_1_bits_addr_beat( BroadcastAcquireTracker_io_inner_grant_bits_addr_beat ),
       .io_in_1_bits_client_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_1_bits_manager_xact_id( BroadcastAcquireTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_1_bits_is_builtin_type( BroadcastAcquireTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_1_bits_g_type( BroadcastAcquireTracker_io_inner_grant_bits_g_type ),
       .io_in_1_bits_data( T226 ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_grant_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_addr_beat ),
       .io_in_0_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_xact_id ),
       .io_in_0_bits_manager_xact_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_manager_xact_id ),
       .io_in_0_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_is_builtin_type ),
       .io_in_0_bits_g_type( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_g_type ),
       .io_in_0_bits_data( T225 ),
       .io_in_0_bits_client_id( BroadcastVoluntaryReleaseTracker_io_inner_grant_bits_client_id ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( LockingRRArbiter_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       .io_out_bits_client_xact_id( LockingRRArbiter_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( LockingRRArbiter_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( LockingRRArbiter_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( LockingRRArbiter_io_out_bits_g_type ),
       //.io_out_bits_data(  )
       .io_out_bits_client_id( LockingRRArbiter_io_out_bits_client_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_4_ready( LockingRRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( BroadcastAcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_addr_block( BroadcastAcquireTracker_3_io_inner_probe_bits_addr_block ),
       .io_in_4_bits_p_type( BroadcastAcquireTracker_3_io_inner_probe_bits_p_type ),
       .io_in_4_bits_client_id( BroadcastAcquireTracker_3_io_inner_probe_bits_client_id ),
       .io_in_3_ready( LockingRRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( BroadcastAcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_addr_block( BroadcastAcquireTracker_2_io_inner_probe_bits_addr_block ),
       .io_in_3_bits_p_type( BroadcastAcquireTracker_2_io_inner_probe_bits_p_type ),
       .io_in_3_bits_client_id( BroadcastAcquireTracker_2_io_inner_probe_bits_client_id ),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( BroadcastAcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_addr_block( BroadcastAcquireTracker_1_io_inner_probe_bits_addr_block ),
       .io_in_2_bits_p_type( BroadcastAcquireTracker_1_io_inner_probe_bits_p_type ),
       .io_in_2_bits_client_id( BroadcastAcquireTracker_1_io_inner_probe_bits_client_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( BroadcastAcquireTracker_io_inner_probe_valid ),
       .io_in_1_bits_addr_block( BroadcastAcquireTracker_io_inner_probe_bits_addr_block ),
       .io_in_1_bits_p_type( BroadcastAcquireTracker_io_inner_probe_bits_p_type ),
       .io_in_1_bits_client_id( BroadcastAcquireTracker_io_inner_probe_bits_client_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( BroadcastVoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_addr_block(  )
       //.io_in_0_bits_p_type(  )
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_addr_block( LockingRRArbiter_1_io_out_bits_addr_block ),
       .io_out_bits_p_type( LockingRRArbiter_1_io_out_bits_p_type ),
       .io_out_bits_client_id( LockingRRArbiter_1_io_out_bits_client_id )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign LockingRRArbiter_1.io_in_0_bits_addr_block = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_p_type = {1{$random}};
    assign LockingRRArbiter_1.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif
  ClientUncachedTileLinkIOArbiter outer_arb(.clk(clk), .reset(reset),
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( BroadcastAcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_addr_block( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_block ),
       .io_in_4_acquire_bits_client_xact_id( BroadcastAcquireTracker_3_io_outer_acquire_bits_client_xact_id ),
       .io_in_4_acquire_bits_addr_beat( BroadcastAcquireTracker_3_io_outer_acquire_bits_addr_beat ),
       .io_in_4_acquire_bits_is_builtin_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_is_builtin_type ),
       .io_in_4_acquire_bits_a_type( BroadcastAcquireTracker_3_io_outer_acquire_bits_a_type ),
       .io_in_4_acquire_bits_union( BroadcastAcquireTracker_3_io_outer_acquire_bits_union ),
       .io_in_4_acquire_bits_data( BroadcastAcquireTracker_3_io_outer_acquire_bits_data ),
       .io_in_4_grant_ready( BroadcastAcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_addr_beat( outer_arb_io_in_4_grant_bits_addr_beat ),
       .io_in_4_grant_bits_client_xact_id( outer_arb_io_in_4_grant_bits_client_xact_id ),
       .io_in_4_grant_bits_manager_xact_id( outer_arb_io_in_4_grant_bits_manager_xact_id ),
       .io_in_4_grant_bits_is_builtin_type( outer_arb_io_in_4_grant_bits_is_builtin_type ),
       .io_in_4_grant_bits_g_type( outer_arb_io_in_4_grant_bits_g_type ),
       .io_in_4_grant_bits_data( outer_arb_io_in_4_grant_bits_data ),
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( BroadcastAcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_addr_block( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_block ),
       .io_in_3_acquire_bits_client_xact_id( BroadcastAcquireTracker_2_io_outer_acquire_bits_client_xact_id ),
       .io_in_3_acquire_bits_addr_beat( BroadcastAcquireTracker_2_io_outer_acquire_bits_addr_beat ),
       .io_in_3_acquire_bits_is_builtin_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_is_builtin_type ),
       .io_in_3_acquire_bits_a_type( BroadcastAcquireTracker_2_io_outer_acquire_bits_a_type ),
       .io_in_3_acquire_bits_union( BroadcastAcquireTracker_2_io_outer_acquire_bits_union ),
       .io_in_3_acquire_bits_data( BroadcastAcquireTracker_2_io_outer_acquire_bits_data ),
       .io_in_3_grant_ready( BroadcastAcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_addr_beat( outer_arb_io_in_3_grant_bits_addr_beat ),
       .io_in_3_grant_bits_client_xact_id( outer_arb_io_in_3_grant_bits_client_xact_id ),
       .io_in_3_grant_bits_manager_xact_id( outer_arb_io_in_3_grant_bits_manager_xact_id ),
       .io_in_3_grant_bits_is_builtin_type( outer_arb_io_in_3_grant_bits_is_builtin_type ),
       .io_in_3_grant_bits_g_type( outer_arb_io_in_3_grant_bits_g_type ),
       .io_in_3_grant_bits_data( outer_arb_io_in_3_grant_bits_data ),
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( BroadcastAcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_addr_block( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_block ),
       .io_in_2_acquire_bits_client_xact_id( BroadcastAcquireTracker_1_io_outer_acquire_bits_client_xact_id ),
       .io_in_2_acquire_bits_addr_beat( BroadcastAcquireTracker_1_io_outer_acquire_bits_addr_beat ),
       .io_in_2_acquire_bits_is_builtin_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_is_builtin_type ),
       .io_in_2_acquire_bits_a_type( BroadcastAcquireTracker_1_io_outer_acquire_bits_a_type ),
       .io_in_2_acquire_bits_union( BroadcastAcquireTracker_1_io_outer_acquire_bits_union ),
       .io_in_2_acquire_bits_data( BroadcastAcquireTracker_1_io_outer_acquire_bits_data ),
       .io_in_2_grant_ready( BroadcastAcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_addr_beat( outer_arb_io_in_2_grant_bits_addr_beat ),
       .io_in_2_grant_bits_client_xact_id( outer_arb_io_in_2_grant_bits_client_xact_id ),
       .io_in_2_grant_bits_manager_xact_id( outer_arb_io_in_2_grant_bits_manager_xact_id ),
       .io_in_2_grant_bits_is_builtin_type( outer_arb_io_in_2_grant_bits_is_builtin_type ),
       .io_in_2_grant_bits_g_type( outer_arb_io_in_2_grant_bits_g_type ),
       .io_in_2_grant_bits_data( outer_arb_io_in_2_grant_bits_data ),
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( BroadcastAcquireTracker_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_addr_block( BroadcastAcquireTracker_io_outer_acquire_bits_addr_block ),
       .io_in_1_acquire_bits_client_xact_id( BroadcastAcquireTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_1_acquire_bits_addr_beat( BroadcastAcquireTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_1_acquire_bits_is_builtin_type( BroadcastAcquireTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_1_acquire_bits_a_type( BroadcastAcquireTracker_io_outer_acquire_bits_a_type ),
       .io_in_1_acquire_bits_union( BroadcastAcquireTracker_io_outer_acquire_bits_union ),
       .io_in_1_acquire_bits_data( BroadcastAcquireTracker_io_outer_acquire_bits_data ),
       .io_in_1_grant_ready( BroadcastAcquireTracker_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_addr_beat( outer_arb_io_in_1_grant_bits_addr_beat ),
       .io_in_1_grant_bits_client_xact_id( outer_arb_io_in_1_grant_bits_client_xact_id ),
       .io_in_1_grant_bits_manager_xact_id( outer_arb_io_in_1_grant_bits_manager_xact_id ),
       .io_in_1_grant_bits_is_builtin_type( outer_arb_io_in_1_grant_bits_is_builtin_type ),
       .io_in_1_grant_bits_g_type( outer_arb_io_in_1_grant_bits_g_type ),
       .io_in_1_grant_bits_data( outer_arb_io_in_1_grant_bits_data ),
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( BroadcastVoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_addr_block( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_block ),
       .io_in_0_acquire_bits_client_xact_id( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_client_xact_id ),
       .io_in_0_acquire_bits_addr_beat( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_addr_beat ),
       .io_in_0_acquire_bits_is_builtin_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_is_builtin_type ),
       .io_in_0_acquire_bits_a_type( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_a_type ),
       .io_in_0_acquire_bits_union( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_union ),
       .io_in_0_acquire_bits_data( BroadcastVoluntaryReleaseTracker_io_outer_acquire_bits_data ),
       .io_in_0_grant_ready( BroadcastVoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_addr_beat( outer_arb_io_in_0_grant_bits_addr_beat ),
       .io_in_0_grant_bits_client_xact_id( outer_arb_io_in_0_grant_bits_client_xact_id ),
       .io_in_0_grant_bits_manager_xact_id( outer_arb_io_in_0_grant_bits_manager_xact_id ),
       .io_in_0_grant_bits_is_builtin_type( outer_arb_io_in_0_grant_bits_is_builtin_type ),
       .io_in_0_grant_bits_g_type( outer_arb_io_in_0_grant_bits_g_type ),
       .io_in_0_grant_bits_data( outer_arb_io_in_0_grant_bits_data ),
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( outer_arb_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( outer_arb_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( outer_arb_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( outer_arb_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( outer_arb_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( outer_arb_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( outer_arb_io_out_acquire_bits_data ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_addr_beat( io_outer_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( io_outer_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( io_outer_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( io_outer_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( io_outer_grant_bits_g_type ),
       .io_out_grant_bits_data( T224 )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Non-voluntary release should always have a Tracker waiting for it.");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      rel_data_cnt <= 2'h0;
    end else if(vwbdq_enq) begin
      rel_data_cnt <= T15;
    end
    if(reset) begin
      sdq_val <= 4'h0;
    end else if(T69) begin
      sdq_val <= T33;
    end
    if(T161) begin
      vwbdq_0 <= io_inner_release_bits_data;
    end
    if(T166) begin
      vwbdq_1 <= io_inner_release_bits_data;
    end
    if(T172) begin
      vwbdq_2 <= io_inner_release_bits_data;
    end
    if(T175) begin
      vwbdq_3 <= io_inner_release_bits_data;
    end
    if(T183) begin
      sdq_0 <= io_inner_acquire_bits_data;
    end
    if(T188) begin
      sdq_1 <= io_inner_acquire_bits_data;
    end
    if(T194) begin
      sdq_2 <= io_inner_acquire_bits_data;
    end
    if(T197) begin
      sdq_3 <= io_inner_acquire_bits_data;
    end
  end
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_len,
    input [2:0] io_enq_bits_size,
    input [1:0] io_enq_bits_burst,
    input  io_enq_bits_lock,
    input [3:0] io_enq_bits_cache,
    input [2:0] io_enq_bits_prot,
    input [3:0] io_enq_bits_qos,
    input [3:0] io_enq_bits_region,
    input [3:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_len,
    output[2:0] io_deq_bits_size,
    output[1:0] io_deq_bits_burst,
    output io_deq_bits_lock,
    output[3:0] io_deq_bits_cache,
    output[2:0] io_deq_bits_prot,
    output[3:0] io_deq_bits_qos,
    output[3:0] io_deq_bits_region,
    output[3:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T37;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T38;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T39;
  wire T8;
  wire T9;
  wire T10;
  wire[65:0] T11;
  reg [65:0] ram [1:0];
  wire[65:0] T12;
  wire[65:0] T13;
  wire[65:0] T14;
  wire[19:0] T15;
  wire[8:0] T16;
  wire[4:0] T17;
  wire[10:0] T18;
  wire[6:0] T19;
  wire[45:0] T20;
  wire[5:0] T21;
  wire[2:0] T22;
  wire[39:0] T23;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[2:0] T27;
  wire[3:0] T28;
  wire T29;
  wire[1:0] T30;
  wire[2:0] T31;
  wire[7:0] T32;
  wire[31:0] T33;
  wire T34;
  wire empty;
  wire T35;
  wire T36;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T37 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T38 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T39 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T20, T15};
  assign T15 = {T18, T16};
  assign T16 = {io_enq_bits_region, T17};
  assign T17 = {io_enq_bits_id, io_enq_bits_user};
  assign T18 = {io_enq_bits_cache, T19};
  assign T19 = {io_enq_bits_prot, io_enq_bits_qos};
  assign T20 = {T23, T21};
  assign T21 = {io_enq_bits_size, T22};
  assign T22 = {io_enq_bits_burst, io_enq_bits_lock};
  assign T23 = {io_enq_bits_addr, io_enq_bits_len};
  assign io_deq_bits_id = T24;
  assign T24 = T11[3'h4:1'h1];
  assign io_deq_bits_region = T25;
  assign T25 = T11[4'h8:3'h5];
  assign io_deq_bits_qos = T26;
  assign T26 = T11[4'hc:4'h9];
  assign io_deq_bits_prot = T27;
  assign T27 = T11[4'hf:4'hd];
  assign io_deq_bits_cache = T28;
  assign T28 = T11[5'h13:5'h10];
  assign io_deq_bits_lock = T29;
  assign T29 = T11[5'h14:5'h14];
  assign io_deq_bits_burst = T30;
  assign T30 = T11[5'h16:5'h15];
  assign io_deq_bits_size = T31;
  assign T31 = T11[5'h19:5'h17];
  assign io_deq_bits_len = T32;
  assign T32 = T11[6'h21:5'h1a];
  assign io_deq_bits_addr = T33;
  assign T33 = T11[7'h41:6'h22];
  assign io_deq_valid = T34;
  assign T34 = empty ^ 1'h1;
  assign empty = ptr_match & T35;
  assign T35 = maybe_full ^ 1'h1;
  assign io_enq_ready = T36;
  assign T36 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [3:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[3:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[3:0] T10;
  reg [3:0] ram [1:0];
  wire[3:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module NastiErrorSlave(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [3:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[3:0] io_b_bits_id,
    //output io_b_bits_user
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [3:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[3:0] io_r_bits_id
    //output io_r_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[31:0] T3;
  wire[247:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire[239:0] T9;
  wire T10;
  wire T11;
  reg  draining;
  wire T39;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg [7:0] beats_left;
  wire[7:0] T40;
  wire[7:0] T22;
  wire[7:0] T23;
  wire T24;
  wire T25;
  reg  responding;
  wire T41;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[7:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire r_queue_io_enq_ready;
  wire r_queue_io_deq_valid;
  wire[7:0] r_queue_io_deq_bits_len;
  wire[3:0] r_queue_io_deq_bits_id;
  wire b_queue_io_enq_ready;
  wire b_queue_io_deq_valid;
  wire[3:0] b_queue_io_deq_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    draining = {1{$random}};
    beats_left = {1{$random}};
    responding = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_r_bits_user = {1{$random}};
//  assign io_b_bits_user = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T2 & T1;
  assign T1 = reset ^ 1'h1;
  assign T2 = io_aw_ready & io_aw_valid;
  assign T3 = io_aw_bits_addr;
  assign T5 = T7 & T6;
  assign T6 = reset ^ 1'h1;
  assign T7 = io_ar_ready & io_ar_valid;
  assign T8 = io_ar_bits_addr;
  assign T10 = io_b_ready & T11;
  assign T11 = draining ^ 1'h1;
  assign T39 = reset ? 1'h0 : T12;
  assign T12 = T15 ? 1'h0 : T13;
  assign T13 = T14 ? 1'h1 : draining;
  assign T14 = io_aw_ready & io_aw_valid;
  assign T15 = T16 & io_w_bits_last;
  assign T16 = io_w_ready & io_w_valid;
  assign T17 = io_aw_valid & T18;
  assign T18 = draining ^ 1'h1;
  assign T19 = T20 & io_r_bits_last;
  assign T20 = io_r_ready & io_r_valid;
  assign io_r_bits_id = r_queue_io_deq_bits_id;
  assign io_r_bits_last = T21;
  assign T21 = beats_left == 8'h0;
  assign T40 = reset ? 8'h0 : T22;
  assign T22 = T32 ? T31 : T23;
  assign T23 = T24 ? r_queue_io_deq_bits_len : beats_left;
  assign T24 = T25 & r_queue_io_deq_valid;
  assign T25 = responding ^ 1'h1;
  assign T41 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h0 : T27;
  assign T27 = T24 ? 1'h1 : responding;
  assign T28 = T30 & T29;
  assign T29 = beats_left == 8'h0;
  assign T30 = io_r_ready & io_r_valid;
  assign T31 = beats_left - 8'h1;
  assign T32 = T30 & T33;
  assign T33 = T29 ^ 1'h1;
  assign io_r_bits_data = 64'h0;
  assign io_r_bits_resp = 2'h3;
  assign io_r_valid = T34;
  assign T34 = r_queue_io_deq_valid & responding;
  assign io_ar_ready = r_queue_io_enq_ready;
  assign io_b_bits_id = b_queue_io_deq_bits;
  assign io_b_bits_resp = 2'h3;
  assign io_b_valid = T35;
  assign T35 = b_queue_io_deq_valid & T36;
  assign T36 = draining ^ 1'h1;
  assign io_w_ready = draining;
  assign io_aw_ready = T37;
  assign T37 = b_queue_io_enq_ready & T38;
  assign T38 = draining ^ 1'h1;
  Queue_2 r_queue(.clk(clk), .reset(reset),
       .io_enq_ready( r_queue_io_enq_ready ),
       .io_enq_valid( io_ar_valid ),
       .io_enq_bits_addr( io_ar_bits_addr ),
       .io_enq_bits_len( io_ar_bits_len ),
       .io_enq_bits_size( io_ar_bits_size ),
       .io_enq_bits_burst( io_ar_bits_burst ),
       .io_enq_bits_lock( io_ar_bits_lock ),
       .io_enq_bits_cache( io_ar_bits_cache ),
       .io_enq_bits_prot( io_ar_bits_prot ),
       .io_enq_bits_qos( io_ar_bits_qos ),
       .io_enq_bits_region( io_ar_bits_region ),
       .io_enq_bits_id( io_ar_bits_id ),
       .io_enq_bits_user( io_ar_bits_user ),
       .io_deq_ready( T19 ),
       .io_deq_valid( r_queue_io_deq_valid ),
       //.io_deq_bits_addr(  )
       .io_deq_bits_len( r_queue_io_deq_bits_len ),
       //.io_deq_bits_size(  )
       //.io_deq_bits_burst(  )
       //.io_deq_bits_lock(  )
       //.io_deq_bits_cache(  )
       //.io_deq_bits_prot(  )
       //.io_deq_bits_qos(  )
       //.io_deq_bits_region(  )
       .io_deq_bits_id( r_queue_io_deq_bits_id )
       //.io_deq_bits_user(  )
       //.io_count(  )
  );
  Queue_6 b_queue(.clk(clk), .reset(reset),
       .io_enq_ready( b_queue_io_enq_ready ),
       .io_enq_valid( T17 ),
       .io_enq_bits( io_aw_bits_id ),
       .io_deq_ready( T10 ),
       .io_deq_valid( b_queue_io_deq_valid ),
       .io_deq_bits( b_queue_io_deq_bits )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      draining <= 1'h0;
    end else if(T15) begin
      draining <= 1'h0;
    end else if(T14) begin
      draining <= 1'h1;
    end
    if(reset) begin
      beats_left <= 8'h0;
    end else if(T32) begin
      beats_left <= T31;
    end else if(T24) begin
      beats_left <= r_queue_io_deq_bits_len;
    end
    if(reset) begin
      responding <= 1'h0;
    end else if(T28) begin
      responding <= 1'h0;
    end else if(T24) begin
      responding <= 1'h1;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T5)
        $fwrite(32'h80000002, "Invalid read address %h\n", T8);
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "Invalid write address %h\n", T3);
// synthesis translate_on
`endif
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [3:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [3:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [3:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [3:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[3:0] io_out_bits_id,
    output io_out_bits_user,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  reg [1:0] last_grant;
  wire[1:0] T89;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[3:0] T23;
  wire T24;
  wire T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T11 ? 2'h1 : T0;
  assign T0 = T9 ? 2'h2 : T1;
  assign T1 = T5 ? 2'h3 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : T4;
  assign T4 = io_in_2_valid ? 2'h2 : 2'h3;
  assign T5 = io_in_3_valid & T6;
  assign T6 = last_grant < 2'h3;
  assign T89 = reset ? 2'h0 : T7;
  assign T7 = T8 ? chosen : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_2_valid & T10;
  assign T10 = last_grant < 2'h2;
  assign T11 = io_in_1_valid & T12;
  assign T12 = last_grant < 2'h1;
  assign io_out_bits_user = T13;
  assign T13 = T19 ? T17 : T14;
  assign T14 = T15 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T15 = T16[1'h0:1'h0];
  assign T16 = chosen;
  assign T17 = T18 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T18 = T16[1'h0:1'h0];
  assign T19 = T16[1'h1:1'h1];
  assign io_out_bits_id = T20;
  assign T20 = T25 ? T23 : T21;
  assign T21 = T22 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T22 = T16[1'h0:1'h0];
  assign T23 = T24 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T24 = T16[1'h0:1'h0];
  assign T25 = T16[1'h1:1'h1];
  assign io_out_bits_resp = T26;
  assign T26 = T31 ? T29 : T27;
  assign T27 = T28 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T28 = T16[1'h0:1'h0];
  assign T29 = T30 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T30 = T16[1'h0:1'h0];
  assign T31 = T16[1'h1:1'h1];
  assign io_out_valid = T32;
  assign T32 = T37 ? T35 : T33;
  assign T33 = T34 ? io_in_1_valid : io_in_0_valid;
  assign T34 = T16[1'h0:1'h0];
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T16[1'h0:1'h0];
  assign T37 = T16[1'h1:1'h1];
  assign io_in_0_ready = T38;
  assign T38 = T39 & io_out_ready;
  assign T39 = T52 | T40;
  assign T40 = T41 ^ 1'h1;
  assign T41 = T44 | T42;
  assign T42 = io_in_3_valid & T43;
  assign T43 = last_grant < 2'h3;
  assign T44 = T47 | T45;
  assign T45 = io_in_2_valid & T46;
  assign T46 = last_grant < 2'h2;
  assign T47 = T50 | T48;
  assign T48 = io_in_1_valid & T49;
  assign T49 = last_grant < 2'h1;
  assign T50 = io_in_0_valid & T51;
  assign T51 = last_grant < 2'h0;
  assign T52 = last_grant < 2'h0;
  assign io_in_1_ready = T53;
  assign T53 = T54 & io_out_ready;
  assign T54 = T60 | T55;
  assign T55 = T56 ^ 1'h1;
  assign T56 = T57 | io_in_0_valid;
  assign T57 = T58 | T42;
  assign T58 = T59 | T45;
  assign T59 = T50 | T48;
  assign T60 = T62 & T61;
  assign T61 = last_grant < 2'h1;
  assign T62 = T50 ^ 1'h1;
  assign io_in_2_ready = T63;
  assign T63 = T64 & io_out_ready;
  assign T64 = T71 | T65;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_1_valid;
  assign T67 = T68 | io_in_0_valid;
  assign T68 = T69 | T42;
  assign T69 = T70 | T45;
  assign T70 = T50 | T48;
  assign T71 = T73 & T72;
  assign T72 = last_grant < 2'h2;
  assign T73 = T74 ^ 1'h1;
  assign T74 = T50 | T48;
  assign io_in_3_ready = T75;
  assign T75 = T76 & io_out_ready;
  assign T76 = T84 | T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T79 | io_in_2_valid;
  assign T79 = T80 | io_in_1_valid;
  assign T80 = T81 | io_in_0_valid;
  assign T81 = T82 | T42;
  assign T82 = T83 | T45;
  assign T83 = T50 | T48;
  assign T84 = T86 & T85;
  assign T85 = last_grant < 2'h3;
  assign T86 = T87 ^ 1'h1;
  assign T87 = T88 | T45;
  assign T88 = T50 | T48;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= chosen;
    end
  end
endmodule

module JunctionsPeekingArbiter(input clk, input reset,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_resp,
    input [63:0] io_in_3_bits_data,
    input  io_in_3_bits_last,
    input [3:0] io_in_3_bits_id,
    input  io_in_3_bits_user,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_resp,
    input [63:0] io_in_2_bits_data,
    input  io_in_2_bits_last,
    input [3:0] io_in_2_bits_id,
    input  io_in_2_bits_user,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_resp,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_last,
    input [3:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_resp,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_last,
    input [3:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_resp,
    output[63:0] io_out_bits_data,
    output io_out_bits_last,
    output[3:0] io_out_bits_id,
    output io_out_bits_user
);

  wire T0;
  wire T1;
  wire T2;
  wire[1:0] T3;
  wire[1:0] chosen;
  wire[1:0] choice;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  reg [1:0] T7;
  wire[1:0] T9;
  wire[1:0] T10;
  reg [1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  reg [1:0] T15;
  wire[1:0] T16;
  reg [1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[1:0] T39;
  reg [1:0] T40;
  wire[1:0] T41;
  reg [1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  reg [1:0] T64;
  wire[1:0] T135;
  wire[2:0] T65;
  wire[2:0] T136;
  reg [1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[2:0] T137;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[1:0] T138;
  wire[2:0] T74;
  wire[2:0] T139;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[2:0] T140;
  reg [1:0] lockIdx;
  wire[1:0] T141;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire T90;
  reg  locked;
  wire T142;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire T99;
  wire[3:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire[63:0] T109;
  wire[63:0] T110;
  wire T111;
  wire[63:0] T112;
  wire T113;
  wire T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_bits_user = T0;
  assign T0 = T96 ? T94 : T1;
  assign T1 = T2 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T2 = T3[1'h0:1'h0];
  assign T3 = chosen;
  assign chosen = locked ? lockIdx : choice;
  assign choice = T69 ? T63 : T4;
  assign T4 = T45 ? T39 : T5;
  assign T5 = T20 ? T14 : T6;
  assign T6 = T13 ? T11 : T7;
  always @(*) case (T9)
    0: T7 = 2'h0;
    1: T7 = 2'h1;
    2: T7 = 2'h2;
    3: T7 = 2'h3;
    default: begin
      T7 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T7 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T9 = T10 - 2'h1;
  assign T10 = lockIdx + 2'h1;
  always @(*) case (T12)
    0: T11 = 2'h0;
    1: T11 = 2'h1;
    2: T11 = 2'h2;
    3: T11 = 2'h3;
    default: begin
      T11 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T11 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T12 = 2'h3 + T10;
  assign T13 = T10 < 2'h1;
  assign T14 = T19 ? T17 : T15;
  always @(*) case (T16)
    0: T15 = 2'h0;
    1: T15 = 2'h1;
    2: T15 = 2'h2;
    3: T15 = 2'h3;
    default: begin
      T15 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T15 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T16 = T10 - 2'h2;
  always @(*) case (T18)
    0: T17 = 2'h0;
    1: T17 = 2'h1;
    2: T17 = 2'h2;
    3: T17 = 2'h3;
    default: begin
      T17 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T17 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T18 = 2'h2 + T10;
  assign T19 = T10 < 2'h2;
  assign T20 = T38 ? T30 : T21;
  assign T21 = T29 ? T27 : T22;
  assign T22 = T23 ? io_in_1_valid : io_in_0_valid;
  assign T23 = T24[1'h0:1'h0];
  assign T24 = T25;
  assign T25 = T26 - 2'h2;
  assign T26 = lockIdx + 2'h1;
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T24[1'h0:1'h0];
  assign T29 = T24[1'h1:1'h1];
  assign T30 = T37 ? T35 : T31;
  assign T31 = T32 ? io_in_1_valid : io_in_0_valid;
  assign T32 = T33[1'h0:1'h0];
  assign T33 = T34;
  assign T34 = 2'h2 + T26;
  assign T35 = T36 ? io_in_3_valid : io_in_2_valid;
  assign T36 = T33[1'h0:1'h0];
  assign T37 = T33[1'h1:1'h1];
  assign T38 = T26 < 2'h2;
  assign T39 = T44 ? T42 : T40;
  always @(*) case (T41)
    0: T40 = 2'h0;
    1: T40 = 2'h1;
    2: T40 = 2'h2;
    3: T40 = 2'h3;
    default: begin
      T40 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T40 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T41 = T10 - 2'h3;
  always @(*) case (T43)
    0: T42 = 2'h0;
    1: T42 = 2'h1;
    2: T42 = 2'h2;
    3: T42 = 2'h3;
    default: begin
      T42 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T42 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T43 = 2'h1 + T10;
  assign T44 = T10 < 2'h3;
  assign T45 = T62 ? T54 : T46;
  assign T46 = T53 ? T51 : T47;
  assign T47 = T48 ? io_in_1_valid : io_in_0_valid;
  assign T48 = T49[1'h0:1'h0];
  assign T49 = T50;
  assign T50 = T26 - 2'h3;
  assign T51 = T52 ? io_in_3_valid : io_in_2_valid;
  assign T52 = T49[1'h0:1'h0];
  assign T53 = T49[1'h1:1'h1];
  assign T54 = T61 ? T59 : T55;
  assign T55 = T56 ? io_in_1_valid : io_in_0_valid;
  assign T56 = T57[1'h0:1'h0];
  assign T57 = T58;
  assign T58 = 2'h1 + T26;
  assign T59 = T60 ? io_in_3_valid : io_in_2_valid;
  assign T60 = T57[1'h0:1'h0];
  assign T61 = T57[1'h1:1'h1];
  assign T62 = T26 < 2'h3;
  assign T63 = T68 ? T66 : T64;
  always @(*) case (T135)
    0: T64 = 2'h0;
    1: T64 = 2'h1;
    2: T64 = 2'h2;
    3: T64 = 2'h3;
    default: begin
      T64 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T64 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T135 = T65[1'h1:1'h0];
  assign T65 = T136 - 3'h4;
  assign T136 = {1'h0, T10};
  always @(*) case (T67)
    0: T66 = 2'h0;
    1: T66 = 2'h1;
    2: T66 = 2'h2;
    3: T66 = 2'h3;
    default: begin
      T66 = 2'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T66 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T67 = 2'h0 + T10;
  assign T68 = T137 < 3'h4;
  assign T137 = {1'h0, T10};
  assign T69 = T86 ? T78 : T70;
  assign T70 = T77 ? T75 : T71;
  assign T71 = T72 ? io_in_1_valid : io_in_0_valid;
  assign T72 = T73[1'h0:1'h0];
  assign T73 = T138;
  assign T138 = T74[1'h1:1'h0];
  assign T74 = T139 - 3'h4;
  assign T139 = {1'h0, T26};
  assign T75 = T76 ? io_in_3_valid : io_in_2_valid;
  assign T76 = T73[1'h0:1'h0];
  assign T77 = T73[1'h1:1'h1];
  assign T78 = T85 ? T83 : T79;
  assign T79 = T80 ? io_in_1_valid : io_in_0_valid;
  assign T80 = T81[1'h0:1'h0];
  assign T81 = T82;
  assign T82 = 2'h0 + T26;
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T81[1'h0:1'h0];
  assign T85 = T81[1'h1:1'h1];
  assign T86 = T140 < 3'h4;
  assign T140 = {1'h0, T26};
  assign T141 = reset ? 2'h0 : T87;
  assign T87 = T88 ? choice : lockIdx;
  assign T88 = T90 & T89;
  assign T89 = locked ^ 1'h1;
  assign T90 = io_out_ready & io_out_valid;
  assign T142 = reset ? 1'h0 : T91;
  assign T91 = T93 ? 1'h0 : T92;
  assign T92 = T88 ? 1'h1 : locked;
  assign T93 = T90 & io_out_bits_last;
  assign T94 = T95 ? io_in_3_bits_user : io_in_2_bits_user;
  assign T95 = T3[1'h0:1'h0];
  assign T96 = T3[1'h1:1'h1];
  assign io_out_bits_id = T97;
  assign T97 = T102 ? T100 : T98;
  assign T98 = T99 ? io_in_1_bits_id : io_in_0_bits_id;
  assign T99 = T3[1'h0:1'h0];
  assign T100 = T101 ? io_in_3_bits_id : io_in_2_bits_id;
  assign T101 = T3[1'h0:1'h0];
  assign T102 = T3[1'h1:1'h1];
  assign io_out_bits_last = T103;
  assign T103 = T108 ? T106 : T104;
  assign T104 = T105 ? io_in_1_bits_last : io_in_0_bits_last;
  assign T105 = T3[1'h0:1'h0];
  assign T106 = T107 ? io_in_3_bits_last : io_in_2_bits_last;
  assign T107 = T3[1'h0:1'h0];
  assign T108 = T3[1'h1:1'h1];
  assign io_out_bits_data = T109;
  assign T109 = T114 ? T112 : T110;
  assign T110 = T111 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T111 = T3[1'h0:1'h0];
  assign T112 = T113 ? io_in_3_bits_data : io_in_2_bits_data;
  assign T113 = T3[1'h0:1'h0];
  assign T114 = T3[1'h1:1'h1];
  assign io_out_bits_resp = T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? io_in_1_bits_resp : io_in_0_bits_resp;
  assign T117 = T3[1'h0:1'h0];
  assign T118 = T119 ? io_in_3_bits_resp : io_in_2_bits_resp;
  assign T119 = T3[1'h0:1'h0];
  assign T120 = T3[1'h1:1'h1];
  assign io_out_valid = T121;
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? io_in_1_valid : io_in_0_valid;
  assign T123 = T3[1'h0:1'h0];
  assign T124 = T125 ? io_in_3_valid : io_in_2_valid;
  assign T125 = T3[1'h0:1'h0];
  assign T126 = T3[1'h1:1'h1];
  assign io_in_0_ready = T127;
  assign T127 = io_out_ready & T128;
  assign T128 = chosen == 2'h0;
  assign io_in_1_ready = T129;
  assign T129 = io_out_ready & T130;
  assign T130 = chosen == 2'h1;
  assign io_in_2_ready = T131;
  assign T131 = io_out_ready & T132;
  assign T132 = chosen == 2'h2;
  assign io_in_3_ready = T133;
  assign T133 = io_out_ready & T134;
  assign T134 = chosen == 2'h3;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h0;
    end else if(T88) begin
      lockIdx <= choice;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T93) begin
      locked <= 1'h0;
    end else if(T88) begin
      locked <= 1'h1;
    end
  end
endmodule

module NastiRouter_0(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [3:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[3:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [3:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[3:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_2_aw_ready,
    output io_slave_2_aw_valid,
    output[31:0] io_slave_2_aw_bits_addr,
    output[7:0] io_slave_2_aw_bits_len,
    output[2:0] io_slave_2_aw_bits_size,
    output[1:0] io_slave_2_aw_bits_burst,
    output io_slave_2_aw_bits_lock,
    output[3:0] io_slave_2_aw_bits_cache,
    output[2:0] io_slave_2_aw_bits_prot,
    output[3:0] io_slave_2_aw_bits_qos,
    output[3:0] io_slave_2_aw_bits_region,
    output[3:0] io_slave_2_aw_bits_id,
    output io_slave_2_aw_bits_user,
    input  io_slave_2_w_ready,
    output io_slave_2_w_valid,
    output[63:0] io_slave_2_w_bits_data,
    output io_slave_2_w_bits_last,
    output[7:0] io_slave_2_w_bits_strb,
    output io_slave_2_w_bits_user,
    output io_slave_2_b_ready,
    input  io_slave_2_b_valid,
    input [1:0] io_slave_2_b_bits_resp,
    input [3:0] io_slave_2_b_bits_id,
    input  io_slave_2_b_bits_user,
    input  io_slave_2_ar_ready,
    output io_slave_2_ar_valid,
    output[31:0] io_slave_2_ar_bits_addr,
    output[7:0] io_slave_2_ar_bits_len,
    output[2:0] io_slave_2_ar_bits_size,
    output[1:0] io_slave_2_ar_bits_burst,
    output io_slave_2_ar_bits_lock,
    output[3:0] io_slave_2_ar_bits_cache,
    output[2:0] io_slave_2_ar_bits_prot,
    output[3:0] io_slave_2_ar_bits_qos,
    output[3:0] io_slave_2_ar_bits_region,
    output[3:0] io_slave_2_ar_bits_id,
    output io_slave_2_ar_bits_user,
    output io_slave_2_r_ready,
    input  io_slave_2_r_valid,
    input [1:0] io_slave_2_r_bits_resp,
    input [63:0] io_slave_2_r_bits_data,
    input  io_slave_2_r_bits_last,
    input [3:0] io_slave_2_r_bits_id,
    input  io_slave_2_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[3:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [3:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[3:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [3:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[3:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [3:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[3:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [3:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[2:0] ar_route;
  wire[2:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[32:0] T82;
  wire T12;
  wire T13;
  wire w_invalid;
  wire T14;
  wire[2:0] aw_route;
  wire[2:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[32:0] T83;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T84;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg  R40;
  wire T85;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  R51;
  wire T86;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire ar_ready;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire w_ready;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire aw_ready;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire b_arb_io_in_3_ready;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[3:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_3_ready;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[3:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[3:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[3:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R29 = {1{$random}};
    R40 = {1{$random}};
    R51 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 3'h0;
  assign ar_route = T2;
  assign T2 = {T10, T3};
  assign T3 = {T7, T4};
  assign T4 = T6 & T5;
  assign T5 = io_master_ar_bits_addr < 32'h40000000;
  assign T6 = 32'h0 <= io_master_ar_bits_addr;
  assign T7 = T9 & T8;
  assign T8 = io_master_ar_bits_addr < 32'h80000000;
  assign T9 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T10 = T12 & T11;
  assign T11 = T82 < 33'h100000000;
  assign T82 = {1'h0, io_master_ar_bits_addr};
  assign T12 = 32'h80000000 <= io_master_ar_bits_addr;
  assign T13 = w_invalid & io_master_aw_valid;
  assign w_invalid = T14 ^ 1'h1;
  assign T14 = aw_route != 3'h0;
  assign aw_route = T15;
  assign T15 = {T23, T16};
  assign T16 = {T20, T17};
  assign T17 = T19 & T18;
  assign T18 = io_master_aw_bits_addr < 32'h40000000;
  assign T19 = 32'h0 <= io_master_aw_bits_addr;
  assign T20 = T22 & T21;
  assign T21 = io_master_aw_bits_addr < 32'h80000000;
  assign T22 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T23 = T25 & T24;
  assign T24 = T83 < 33'h100000000;
  assign T83 = {1'h0, io_master_aw_bits_addr};
  assign T25 = 32'h80000000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T26;
  assign T26 = io_master_ar_valid & T27;
  assign T27 = ar_route[1'h0:1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T28;
  assign T28 = io_master_w_valid & R29;
  assign T84 = reset ? 1'h0 : T30;
  assign T30 = T33 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : R29;
  assign T32 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T33 = T34 & io_slave_0_w_bits_last;
  assign T34 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T35;
  assign T35 = io_master_aw_valid & T36;
  assign T36 = aw_route[1'h0:1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T37;
  assign T37 = io_master_ar_valid & T38;
  assign T38 = ar_route[1'h1:1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T39;
  assign T39 = io_master_w_valid & R40;
  assign T85 = reset ? 1'h0 : T41;
  assign T41 = T44 ? 1'h0 : T42;
  assign T42 = T43 ? 1'h1 : R40;
  assign T43 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T44 = T45 & io_slave_1_w_bits_last;
  assign T45 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T46;
  assign T46 = io_master_aw_valid & T47;
  assign T47 = aw_route[1'h1:1'h1];
  assign io_slave_2_r_ready = r_arb_io_in_2_ready;
  assign io_slave_2_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_2_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_2_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_2_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_2_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_2_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_2_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_2_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_2_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_2_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_2_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_2_ar_valid = T48;
  assign T48 = io_master_ar_valid & T49;
  assign T49 = ar_route[2'h2:2'h2];
  assign io_slave_2_b_ready = b_arb_io_in_2_ready;
  assign io_slave_2_w_bits_user = io_master_w_bits_user;
  assign io_slave_2_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_2_w_bits_last = io_master_w_bits_last;
  assign io_slave_2_w_bits_data = io_master_w_bits_data;
  assign io_slave_2_w_valid = T50;
  assign T50 = io_master_w_valid & R51;
  assign T86 = reset ? 1'h0 : T52;
  assign T52 = T55 ? 1'h0 : T53;
  assign T53 = T54 ? 1'h1 : R51;
  assign T54 = io_slave_2_aw_ready & io_slave_2_aw_valid;
  assign T55 = T56 & io_slave_2_w_bits_last;
  assign T56 = io_slave_2_w_ready & io_slave_2_w_valid;
  assign io_slave_2_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_2_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_2_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_2_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_2_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_2_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_2_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_2_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_2_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_2_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_2_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_2_aw_valid = T57;
  assign T57 = io_master_aw_valid & T58;
  assign T58 = aw_route[2'h2:2'h2];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T59;
  assign T59 = ar_ready | T60;
  assign T60 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T63 | T61;
  assign T61 = io_slave_2_ar_ready & T62;
  assign T62 = ar_route[2'h2:2'h2];
  assign T63 = T66 | T64;
  assign T64 = io_slave_1_ar_ready & T65;
  assign T65 = ar_route[1'h1:1'h1];
  assign T66 = io_slave_0_ar_ready & T67;
  assign T67 = ar_route[1'h0:1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T68;
  assign T68 = w_ready | err_slave_io_w_ready;
  assign w_ready = T70 | T69;
  assign T69 = io_slave_2_w_ready & R51;
  assign T70 = T72 | T71;
  assign T71 = io_slave_1_w_ready & R40;
  assign T72 = io_slave_0_w_ready & R29;
  assign io_master_aw_ready = T73;
  assign T73 = aw_ready | T74;
  assign T74 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T77 | T75;
  assign T75 = io_slave_2_aw_ready & T76;
  assign T76 = aw_route[2'h2:2'h2];
  assign T77 = T80 | T78;
  assign T78 = io_slave_1_aw_ready & T79;
  assign T79 = aw_route[1'h1:1'h1];
  assign T80 = io_slave_0_aw_ready & T81;
  assign T81 = aw_route[1'h0:1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T13 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_3_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_3_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_4 b_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( b_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_b_valid ),
       .io_in_3_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_3_bits_id( err_slave_io_b_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_b_valid ),
       .io_in_2_bits_resp( io_slave_2_b_bits_resp ),
       .io_in_2_bits_id( io_slave_2_b_bits_id ),
       .io_in_2_bits_user( io_slave_2_b_bits_user ),
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter r_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( r_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_r_valid ),
       .io_in_3_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_3_bits_data( err_slave_io_r_bits_data ),
       .io_in_3_bits_last( err_slave_io_r_bits_last ),
       .io_in_3_bits_id( err_slave_io_r_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_r_valid ),
       .io_in_2_bits_resp( io_slave_2_r_bits_resp ),
       .io_in_2_bits_data( io_slave_2_r_bits_data ),
       .io_in_2_bits_last( io_slave_2_r_bits_last ),
       .io_in_2_bits_id( io_slave_2_r_bits_id ),
       .io_in_2_bits_user( io_slave_2_r_bits_user ),
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R29 <= 1'h0;
    end else if(T33) begin
      R29 <= 1'h0;
    end else if(T32) begin
      R29 <= 1'h1;
    end
    if(reset) begin
      R40 <= 1'h0;
    end else if(T44) begin
      R40 <= 1'h0;
    end else if(T43) begin
      R40 <= 1'h1;
    end
    if(reset) begin
      R51 <= 1'h0;
    end else if(T55) begin
      R51 <= 1'h0;
    end else if(T54) begin
      R51 <= 1'h1;
    end
  end
endmodule

module RRArbiter_5(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [31:0] io_in_1_bits_addr,
    input [7:0] io_in_1_bits_len,
    input [2:0] io_in_1_bits_size,
    input [1:0] io_in_1_bits_burst,
    input  io_in_1_bits_lock,
    input [3:0] io_in_1_bits_cache,
    input [2:0] io_in_1_bits_prot,
    input [3:0] io_in_1_bits_qos,
    input [3:0] io_in_1_bits_region,
    input [3:0] io_in_1_bits_id,
    input  io_in_1_bits_user,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [31:0] io_in_0_bits_addr,
    input [7:0] io_in_0_bits_len,
    input [2:0] io_in_0_bits_size,
    input [1:0] io_in_0_bits_burst,
    input  io_in_0_bits_lock,
    input [3:0] io_in_0_bits_cache,
    input [2:0] io_in_0_bits_prot,
    input [3:0] io_in_0_bits_qos,
    input [3:0] io_in_0_bits_region,
    input [3:0] io_in_0_bits_id,
    input  io_in_0_bits_user,
    input  io_out_ready,
    output io_out_valid,
    output[31:0] io_out_bits_addr,
    output[7:0] io_out_bits_len,
    output[2:0] io_out_bits_size,
    output[1:0] io_out_bits_burst,
    output io_out_bits_lock,
    output[3:0] io_out_bits_cache,
    output[2:0] io_out_bits_prot,
    output[3:0] io_out_bits_qos,
    output[3:0] io_out_bits_region,
    output[3:0] io_out_bits_id,
    output io_out_bits_user,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T35;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[2:0] T10;
  wire[3:0] T11;
  wire T12;
  wire[1:0] T13;
  wire[2:0] T14;
  wire[7:0] T15;
  wire[31:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T35 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_user = T5;
  assign T5 = T6 ? io_in_1_bits_user : io_in_0_bits_user;
  assign T6 = chosen;
  assign io_out_bits_id = T7;
  assign T7 = T6 ? io_in_1_bits_id : io_in_0_bits_id;
  assign io_out_bits_region = T8;
  assign T8 = T6 ? io_in_1_bits_region : io_in_0_bits_region;
  assign io_out_bits_qos = T9;
  assign T9 = T6 ? io_in_1_bits_qos : io_in_0_bits_qos;
  assign io_out_bits_prot = T10;
  assign T10 = T6 ? io_in_1_bits_prot : io_in_0_bits_prot;
  assign io_out_bits_cache = T11;
  assign T11 = T6 ? io_in_1_bits_cache : io_in_0_bits_cache;
  assign io_out_bits_lock = T12;
  assign T12 = T6 ? io_in_1_bits_lock : io_in_0_bits_lock;
  assign io_out_bits_burst = T13;
  assign T13 = T6 ? io_in_1_bits_burst : io_in_0_bits_burst;
  assign io_out_bits_size = T14;
  assign T14 = T6 ? io_in_1_bits_size : io_in_0_bits_size;
  assign io_out_bits_len = T15;
  assign T15 = T6 ? io_in_1_bits_len : io_in_0_bits_len;
  assign io_out_bits_addr = T16;
  assign T16 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T17;
  assign T17 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T18;
  assign T18 = T19 & io_out_ready;
  assign T19 = T26 | T20;
  assign T20 = T21 ^ 1'h1;
  assign T21 = T24 | T22;
  assign T22 = io_in_1_valid & T23;
  assign T23 = last_grant < 1'h1;
  assign T24 = io_in_0_valid & T25;
  assign T25 = last_grant < 1'h0;
  assign T26 = last_grant < 1'h0;
  assign io_in_1_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T32 | T29;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_0_valid;
  assign T31 = T24 | T22;
  assign T32 = T34 & T33;
  assign T33 = last_grant < 1'h1;
  assign T34 = T24 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module NastiArbiter(input clk, input reset,
    output io_master_1_aw_ready,
    input  io_master_1_aw_valid,
    input [31:0] io_master_1_aw_bits_addr,
    input [7:0] io_master_1_aw_bits_len,
    input [2:0] io_master_1_aw_bits_size,
    input [1:0] io_master_1_aw_bits_burst,
    input  io_master_1_aw_bits_lock,
    input [3:0] io_master_1_aw_bits_cache,
    input [2:0] io_master_1_aw_bits_prot,
    input [3:0] io_master_1_aw_bits_qos,
    input [3:0] io_master_1_aw_bits_region,
    input [3:0] io_master_1_aw_bits_id,
    input  io_master_1_aw_bits_user,
    output io_master_1_w_ready,
    input  io_master_1_w_valid,
    input [63:0] io_master_1_w_bits_data,
    input  io_master_1_w_bits_last,
    input [7:0] io_master_1_w_bits_strb,
    input  io_master_1_w_bits_user,
    input  io_master_1_b_ready,
    output io_master_1_b_valid,
    output[1:0] io_master_1_b_bits_resp,
    output[3:0] io_master_1_b_bits_id,
    output io_master_1_b_bits_user,
    output io_master_1_ar_ready,
    input  io_master_1_ar_valid,
    input [31:0] io_master_1_ar_bits_addr,
    input [7:0] io_master_1_ar_bits_len,
    input [2:0] io_master_1_ar_bits_size,
    input [1:0] io_master_1_ar_bits_burst,
    input  io_master_1_ar_bits_lock,
    input [3:0] io_master_1_ar_bits_cache,
    input [2:0] io_master_1_ar_bits_prot,
    input [3:0] io_master_1_ar_bits_qos,
    input [3:0] io_master_1_ar_bits_region,
    input [3:0] io_master_1_ar_bits_id,
    input  io_master_1_ar_bits_user,
    input  io_master_1_r_ready,
    output io_master_1_r_valid,
    output[1:0] io_master_1_r_bits_resp,
    output[63:0] io_master_1_r_bits_data,
    output io_master_1_r_bits_last,
    output[3:0] io_master_1_r_bits_id,
    output io_master_1_r_bits_user,
    output io_master_0_aw_ready,
    input  io_master_0_aw_valid,
    input [31:0] io_master_0_aw_bits_addr,
    input [7:0] io_master_0_aw_bits_len,
    input [2:0] io_master_0_aw_bits_size,
    input [1:0] io_master_0_aw_bits_burst,
    input  io_master_0_aw_bits_lock,
    input [3:0] io_master_0_aw_bits_cache,
    input [2:0] io_master_0_aw_bits_prot,
    input [3:0] io_master_0_aw_bits_qos,
    input [3:0] io_master_0_aw_bits_region,
    input [3:0] io_master_0_aw_bits_id,
    input  io_master_0_aw_bits_user,
    output io_master_0_w_ready,
    input  io_master_0_w_valid,
    input [63:0] io_master_0_w_bits_data,
    input  io_master_0_w_bits_last,
    input [7:0] io_master_0_w_bits_strb,
    input  io_master_0_w_bits_user,
    input  io_master_0_b_ready,
    output io_master_0_b_valid,
    output[1:0] io_master_0_b_bits_resp,
    output[3:0] io_master_0_b_bits_id,
    output io_master_0_b_bits_user,
    output io_master_0_ar_ready,
    input  io_master_0_ar_valid,
    input [31:0] io_master_0_ar_bits_addr,
    input [7:0] io_master_0_ar_bits_len,
    input [2:0] io_master_0_ar_bits_size,
    input [1:0] io_master_0_ar_bits_burst,
    input  io_master_0_ar_bits_lock,
    input [3:0] io_master_0_ar_bits_cache,
    input [2:0] io_master_0_ar_bits_prot,
    input [3:0] io_master_0_ar_bits_qos,
    input [3:0] io_master_0_ar_bits_region,
    input [3:0] io_master_0_ar_bits_id,
    input  io_master_0_ar_bits_user,
    input  io_master_0_r_ready,
    output io_master_0_r_valid,
    output[1:0] io_master_0_r_bits_resp,
    output[63:0] io_master_0_r_bits_data,
    output io_master_0_r_bits_last,
    output[3:0] io_master_0_r_bits_id,
    output io_master_0_r_bits_user,
    input  io_slave_aw_ready,
    output io_slave_aw_valid,
    output[31:0] io_slave_aw_bits_addr,
    output[7:0] io_slave_aw_bits_len,
    output[2:0] io_slave_aw_bits_size,
    output[1:0] io_slave_aw_bits_burst,
    output io_slave_aw_bits_lock,
    output[3:0] io_slave_aw_bits_cache,
    output[2:0] io_slave_aw_bits_prot,
    output[3:0] io_slave_aw_bits_qos,
    output[3:0] io_slave_aw_bits_region,
    output[3:0] io_slave_aw_bits_id,
    output io_slave_aw_bits_user,
    input  io_slave_w_ready,
    output io_slave_w_valid,
    output[63:0] io_slave_w_bits_data,
    output io_slave_w_bits_last,
    output[7:0] io_slave_w_bits_strb,
    output io_slave_w_bits_user,
    output io_slave_b_ready,
    input  io_slave_b_valid,
    input [1:0] io_slave_b_bits_resp,
    input [3:0] io_slave_b_bits_id,
    input  io_slave_b_bits_user,
    input  io_slave_ar_ready,
    output io_slave_ar_valid,
    output[31:0] io_slave_ar_bits_addr,
    output[7:0] io_slave_ar_bits_len,
    output[2:0] io_slave_ar_bits_size,
    output[1:0] io_slave_ar_bits_burst,
    output io_slave_ar_bits_lock,
    output[3:0] io_slave_ar_bits_cache,
    output[2:0] io_slave_ar_bits_prot,
    output[3:0] io_slave_ar_bits_qos,
    output[3:0] io_slave_ar_bits_region,
    output[3:0] io_slave_ar_bits_id,
    output io_slave_ar_bits_user,
    output io_slave_r_ready,
    input  io_slave_r_valid,
    input [1:0] io_slave_r_bits_resp,
    input [63:0] io_slave_r_bits_data,
    input  io_slave_r_bits_last,
    input [3:0] io_slave_r_bits_id,
    input  io_slave_r_bits_user
);

  wire T0;
  reg  R1;
  wire T48;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[3:0] T49;
  wire[4:0] T7;
  wire[3:0] T50;
  wire[4:0] T8;
  wire[3:0] T51;
  wire[4:0] T9;
  wire[3:0] T52;
  wire[4:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg  R19;
  wire T20;
  wire[7:0] T21;
  wire T22;
  wire[63:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[3:0] T53;
  wire[2:0] T28;
  wire T29;
  wire T30;
  wire[3:0] T54;
  wire[2:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[3:0] T55;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire[3:0] T56;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire RRArbiter_io_in_1_ready;
  wire RRArbiter_io_in_0_ready;
  wire RRArbiter_io_out_valid;
  wire[31:0] RRArbiter_io_out_bits_addr;
  wire[7:0] RRArbiter_io_out_bits_len;
  wire[2:0] RRArbiter_io_out_bits_size;
  wire[1:0] RRArbiter_io_out_bits_burst;
  wire RRArbiter_io_out_bits_lock;
  wire[3:0] RRArbiter_io_out_bits_cache;
  wire[2:0] RRArbiter_io_out_bits_prot;
  wire[3:0] RRArbiter_io_out_bits_qos;
  wire[3:0] RRArbiter_io_out_bits_region;
  wire[3:0] RRArbiter_io_out_bits_id;
  wire RRArbiter_io_out_bits_user;
  wire RRArbiter_1_io_in_1_ready;
  wire RRArbiter_1_io_in_0_ready;
  wire RRArbiter_1_io_out_valid;
  wire[31:0] RRArbiter_1_io_out_bits_addr;
  wire[7:0] RRArbiter_1_io_out_bits_len;
  wire[2:0] RRArbiter_1_io_out_bits_size;
  wire[1:0] RRArbiter_1_io_out_bits_burst;
  wire RRArbiter_1_io_out_bits_lock;
  wire[3:0] RRArbiter_1_io_out_bits_cache;
  wire[2:0] RRArbiter_1_io_out_bits_prot;
  wire[3:0] RRArbiter_1_io_out_bits_qos;
  wire[3:0] RRArbiter_1_io_out_bits_region;
  wire[3:0] RRArbiter_1_io_out_bits_id;
  wire RRArbiter_1_io_out_bits_user;
  wire RRArbiter_1_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R19 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_slave_aw_ready & R1;
  assign T48 = reset ? 1'h1 : T2;
  assign T2 = T5 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : R1;
  assign T4 = T0 & RRArbiter_1_io_out_valid;
  assign T5 = T6 & io_slave_w_bits_last;
  assign T6 = io_slave_w_ready & io_slave_w_valid;
  assign T49 = T7[2'h3:1'h0];
  assign T7 = {io_master_0_aw_bits_id, 1'h0};
  assign T50 = T8[2'h3:1'h0];
  assign T8 = {io_master_1_aw_bits_id, 1'h1};
  assign T51 = T9[2'h3:1'h0];
  assign T9 = {io_master_0_ar_bits_id, 1'h0};
  assign T52 = T10[2'h3:1'h0];
  assign T10 = {io_master_1_ar_bits_id, 1'h1};
  assign io_slave_r_ready = T11;
  assign T11 = T12 ? io_master_1_r_ready : io_master_0_r_ready;
  assign T12 = T13;
  assign T13 = io_slave_r_bits_id[1'h0:1'h0];
  assign io_slave_ar_bits_user = RRArbiter_io_out_bits_user;
  assign io_slave_ar_bits_id = RRArbiter_io_out_bits_id;
  assign io_slave_ar_bits_region = RRArbiter_io_out_bits_region;
  assign io_slave_ar_bits_qos = RRArbiter_io_out_bits_qos;
  assign io_slave_ar_bits_prot = RRArbiter_io_out_bits_prot;
  assign io_slave_ar_bits_cache = RRArbiter_io_out_bits_cache;
  assign io_slave_ar_bits_lock = RRArbiter_io_out_bits_lock;
  assign io_slave_ar_bits_burst = RRArbiter_io_out_bits_burst;
  assign io_slave_ar_bits_size = RRArbiter_io_out_bits_size;
  assign io_slave_ar_bits_len = RRArbiter_io_out_bits_len;
  assign io_slave_ar_bits_addr = RRArbiter_io_out_bits_addr;
  assign io_slave_ar_valid = RRArbiter_io_out_valid;
  assign io_slave_b_ready = T14;
  assign T14 = T15 ? io_master_1_b_ready : io_master_0_b_ready;
  assign T15 = T16;
  assign T16 = io_slave_b_bits_id[1'h0:1'h0];
  assign io_slave_w_bits_user = T17;
  assign T17 = T18 ? io_master_1_w_bits_user : io_master_0_w_bits_user;
  assign T18 = R19;
  assign T20 = T4 ? RRArbiter_1_io_chosen : R19;
  assign io_slave_w_bits_strb = T21;
  assign T21 = T18 ? io_master_1_w_bits_strb : io_master_0_w_bits_strb;
  assign io_slave_w_bits_last = T22;
  assign T22 = T18 ? io_master_1_w_bits_last : io_master_0_w_bits_last;
  assign io_slave_w_bits_data = T23;
  assign T23 = T18 ? io_master_1_w_bits_data : io_master_0_w_bits_data;
  assign io_slave_w_valid = T24;
  assign T24 = T26 & T25;
  assign T25 = R1 ^ 1'h1;
  assign T26 = T18 ? io_master_1_w_valid : io_master_0_w_valid;
  assign io_slave_aw_bits_user = RRArbiter_1_io_out_bits_user;
  assign io_slave_aw_bits_id = RRArbiter_1_io_out_bits_id;
  assign io_slave_aw_bits_region = RRArbiter_1_io_out_bits_region;
  assign io_slave_aw_bits_qos = RRArbiter_1_io_out_bits_qos;
  assign io_slave_aw_bits_prot = RRArbiter_1_io_out_bits_prot;
  assign io_slave_aw_bits_cache = RRArbiter_1_io_out_bits_cache;
  assign io_slave_aw_bits_lock = RRArbiter_1_io_out_bits_lock;
  assign io_slave_aw_bits_burst = RRArbiter_1_io_out_bits_burst;
  assign io_slave_aw_bits_size = RRArbiter_1_io_out_bits_size;
  assign io_slave_aw_bits_len = RRArbiter_1_io_out_bits_len;
  assign io_slave_aw_bits_addr = RRArbiter_1_io_out_bits_addr;
  assign io_slave_aw_valid = T27;
  assign T27 = RRArbiter_1_io_out_valid & R1;
  assign io_master_0_r_bits_user = io_slave_r_bits_user;
  assign io_master_0_r_bits_id = T53;
  assign T53 = {1'h0, T28};
  assign T28 = io_slave_r_bits_id >> 1'h1;
  assign io_master_0_r_bits_last = io_slave_r_bits_last;
  assign io_master_0_r_bits_data = io_slave_r_bits_data;
  assign io_master_0_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_0_r_valid = T29;
  assign T29 = io_slave_r_valid & T30;
  assign T30 = T13 == 1'h0;
  assign io_master_0_ar_ready = RRArbiter_io_in_0_ready;
  assign io_master_0_b_bits_user = io_slave_b_bits_user;
  assign io_master_0_b_bits_id = T54;
  assign T54 = {1'h0, T31};
  assign T31 = io_slave_b_bits_id >> 1'h1;
  assign io_master_0_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_0_b_valid = T32;
  assign T32 = io_slave_b_valid & T33;
  assign T33 = T16 == 1'h0;
  assign io_master_0_w_ready = T34;
  assign T34 = T36 & T35;
  assign T35 = R1 ^ 1'h1;
  assign T36 = io_slave_w_ready & T37;
  assign T37 = R19 == 1'h0;
  assign io_master_0_aw_ready = RRArbiter_1_io_in_0_ready;
  assign io_master_1_r_bits_user = io_slave_r_bits_user;
  assign io_master_1_r_bits_id = T55;
  assign T55 = {1'h0, T38};
  assign T38 = io_slave_r_bits_id >> 1'h1;
  assign io_master_1_r_bits_last = io_slave_r_bits_last;
  assign io_master_1_r_bits_data = io_slave_r_bits_data;
  assign io_master_1_r_bits_resp = io_slave_r_bits_resp;
  assign io_master_1_r_valid = T39;
  assign T39 = io_slave_r_valid & T40;
  assign T40 = T13 == 1'h1;
  assign io_master_1_ar_ready = RRArbiter_io_in_1_ready;
  assign io_master_1_b_bits_user = io_slave_b_bits_user;
  assign io_master_1_b_bits_id = T56;
  assign T56 = {1'h0, T41};
  assign T41 = io_slave_b_bits_id >> 1'h1;
  assign io_master_1_b_bits_resp = io_slave_b_bits_resp;
  assign io_master_1_b_valid = T42;
  assign T42 = io_slave_b_valid & T43;
  assign T43 = T16 == 1'h1;
  assign io_master_1_w_ready = T44;
  assign T44 = T46 & T45;
  assign T45 = R1 ^ 1'h1;
  assign T46 = io_slave_w_ready & T47;
  assign T47 = R19 == 1'h1;
  assign io_master_1_aw_ready = RRArbiter_1_io_in_1_ready;
  RRArbiter_5 RRArbiter(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_io_in_1_ready ),
       .io_in_1_valid( io_master_1_ar_valid ),
       .io_in_1_bits_addr( io_master_1_ar_bits_addr ),
       .io_in_1_bits_len( io_master_1_ar_bits_len ),
       .io_in_1_bits_size( io_master_1_ar_bits_size ),
       .io_in_1_bits_burst( io_master_1_ar_bits_burst ),
       .io_in_1_bits_lock( io_master_1_ar_bits_lock ),
       .io_in_1_bits_cache( io_master_1_ar_bits_cache ),
       .io_in_1_bits_prot( io_master_1_ar_bits_prot ),
       .io_in_1_bits_qos( io_master_1_ar_bits_qos ),
       .io_in_1_bits_region( io_master_1_ar_bits_region ),
       .io_in_1_bits_id( T52 ),
       .io_in_1_bits_user( io_master_1_ar_bits_user ),
       .io_in_0_ready( RRArbiter_io_in_0_ready ),
       .io_in_0_valid( io_master_0_ar_valid ),
       .io_in_0_bits_addr( io_master_0_ar_bits_addr ),
       .io_in_0_bits_len( io_master_0_ar_bits_len ),
       .io_in_0_bits_size( io_master_0_ar_bits_size ),
       .io_in_0_bits_burst( io_master_0_ar_bits_burst ),
       .io_in_0_bits_lock( io_master_0_ar_bits_lock ),
       .io_in_0_bits_cache( io_master_0_ar_bits_cache ),
       .io_in_0_bits_prot( io_master_0_ar_bits_prot ),
       .io_in_0_bits_qos( io_master_0_ar_bits_qos ),
       .io_in_0_bits_region( io_master_0_ar_bits_region ),
       .io_in_0_bits_id( T51 ),
       .io_in_0_bits_user( io_master_0_ar_bits_user ),
       .io_out_ready( io_slave_ar_ready ),
       .io_out_valid( RRArbiter_io_out_valid ),
       .io_out_bits_addr( RRArbiter_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_io_out_bits_user )
       //.io_chosen(  )
  );
  RRArbiter_5 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_master_1_aw_valid ),
       .io_in_1_bits_addr( io_master_1_aw_bits_addr ),
       .io_in_1_bits_len( io_master_1_aw_bits_len ),
       .io_in_1_bits_size( io_master_1_aw_bits_size ),
       .io_in_1_bits_burst( io_master_1_aw_bits_burst ),
       .io_in_1_bits_lock( io_master_1_aw_bits_lock ),
       .io_in_1_bits_cache( io_master_1_aw_bits_cache ),
       .io_in_1_bits_prot( io_master_1_aw_bits_prot ),
       .io_in_1_bits_qos( io_master_1_aw_bits_qos ),
       .io_in_1_bits_region( io_master_1_aw_bits_region ),
       .io_in_1_bits_id( T50 ),
       .io_in_1_bits_user( io_master_1_aw_bits_user ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_master_0_aw_valid ),
       .io_in_0_bits_addr( io_master_0_aw_bits_addr ),
       .io_in_0_bits_len( io_master_0_aw_bits_len ),
       .io_in_0_bits_size( io_master_0_aw_bits_size ),
       .io_in_0_bits_burst( io_master_0_aw_bits_burst ),
       .io_in_0_bits_lock( io_master_0_aw_bits_lock ),
       .io_in_0_bits_cache( io_master_0_aw_bits_cache ),
       .io_in_0_bits_prot( io_master_0_aw_bits_prot ),
       .io_in_0_bits_qos( io_master_0_aw_bits_qos ),
       .io_in_0_bits_region( io_master_0_aw_bits_region ),
       .io_in_0_bits_id( T49 ),
       .io_in_0_bits_user( io_master_0_aw_bits_user ),
       .io_out_ready( T0 ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_addr( RRArbiter_1_io_out_bits_addr ),
       .io_out_bits_len( RRArbiter_1_io_out_bits_len ),
       .io_out_bits_size( RRArbiter_1_io_out_bits_size ),
       .io_out_bits_burst( RRArbiter_1_io_out_bits_burst ),
       .io_out_bits_lock( RRArbiter_1_io_out_bits_lock ),
       .io_out_bits_cache( RRArbiter_1_io_out_bits_cache ),
       .io_out_bits_prot( RRArbiter_1_io_out_bits_prot ),
       .io_out_bits_qos( RRArbiter_1_io_out_bits_qos ),
       .io_out_bits_region( RRArbiter_1_io_out_bits_region ),
       .io_out_bits_id( RRArbiter_1_io_out_bits_id ),
       .io_out_bits_user( RRArbiter_1_io_out_bits_user ),
       .io_chosen( RRArbiter_1_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h1;
    end else if(T5) begin
      R1 <= 1'h1;
    end else if(T4) begin
      R1 <= 1'h0;
    end
    if(T4) begin
      R19 <= RRArbiter_1_io_chosen;
    end
  end
endmodule

module NastiCrossbar_0(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [3:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[3:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [3:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[3:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [3:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[3:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [3:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[3:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[3:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [3:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[3:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [3:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[3:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [3:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[3:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [3:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[3:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [3:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[3:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [3:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiArbiter_io_master_1_aw_ready;
  wire NastiArbiter_io_master_1_w_ready;
  wire NastiArbiter_io_master_1_b_valid;
  wire[1:0] NastiArbiter_io_master_1_b_bits_resp;
  wire[3:0] NastiArbiter_io_master_1_b_bits_id;
  wire NastiArbiter_io_master_1_b_bits_user;
  wire NastiArbiter_io_master_1_ar_ready;
  wire NastiArbiter_io_master_1_r_valid;
  wire[1:0] NastiArbiter_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_1_r_bits_data;
  wire NastiArbiter_io_master_1_r_bits_last;
  wire[3:0] NastiArbiter_io_master_1_r_bits_id;
  wire NastiArbiter_io_master_1_r_bits_user;
  wire NastiArbiter_io_master_0_aw_ready;
  wire NastiArbiter_io_master_0_w_ready;
  wire NastiArbiter_io_master_0_b_valid;
  wire[1:0] NastiArbiter_io_master_0_b_bits_resp;
  wire[3:0] NastiArbiter_io_master_0_b_bits_id;
  wire NastiArbiter_io_master_0_b_bits_user;
  wire NastiArbiter_io_master_0_ar_ready;
  wire NastiArbiter_io_master_0_r_valid;
  wire[1:0] NastiArbiter_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_io_master_0_r_bits_data;
  wire NastiArbiter_io_master_0_r_bits_last;
  wire[3:0] NastiArbiter_io_master_0_r_bits_id;
  wire NastiArbiter_io_master_0_r_bits_user;
  wire NastiArbiter_io_slave_aw_valid;
  wire[31:0] NastiArbiter_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_io_slave_aw_bits_burst;
  wire NastiArbiter_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_io_slave_aw_bits_region;
  wire[3:0] NastiArbiter_io_slave_aw_bits_id;
  wire NastiArbiter_io_slave_aw_bits_user;
  wire NastiArbiter_io_slave_w_valid;
  wire[63:0] NastiArbiter_io_slave_w_bits_data;
  wire NastiArbiter_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_io_slave_w_bits_strb;
  wire NastiArbiter_io_slave_w_bits_user;
  wire NastiArbiter_io_slave_b_ready;
  wire NastiArbiter_io_slave_ar_valid;
  wire[31:0] NastiArbiter_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_io_slave_ar_bits_burst;
  wire NastiArbiter_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_io_slave_ar_bits_region;
  wire[3:0] NastiArbiter_io_slave_ar_bits_id;
  wire NastiArbiter_io_slave_ar_bits_user;
  wire NastiArbiter_io_slave_r_ready;
  wire NastiArbiter_1_io_master_1_aw_ready;
  wire NastiArbiter_1_io_master_1_w_ready;
  wire NastiArbiter_1_io_master_1_b_valid;
  wire[1:0] NastiArbiter_1_io_master_1_b_bits_resp;
  wire[3:0] NastiArbiter_1_io_master_1_b_bits_id;
  wire NastiArbiter_1_io_master_1_b_bits_user;
  wire NastiArbiter_1_io_master_1_ar_ready;
  wire NastiArbiter_1_io_master_1_r_valid;
  wire[1:0] NastiArbiter_1_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_1_r_bits_data;
  wire NastiArbiter_1_io_master_1_r_bits_last;
  wire[3:0] NastiArbiter_1_io_master_1_r_bits_id;
  wire NastiArbiter_1_io_master_1_r_bits_user;
  wire NastiArbiter_1_io_master_0_aw_ready;
  wire NastiArbiter_1_io_master_0_w_ready;
  wire NastiArbiter_1_io_master_0_b_valid;
  wire[1:0] NastiArbiter_1_io_master_0_b_bits_resp;
  wire[3:0] NastiArbiter_1_io_master_0_b_bits_id;
  wire NastiArbiter_1_io_master_0_b_bits_user;
  wire NastiArbiter_1_io_master_0_ar_ready;
  wire NastiArbiter_1_io_master_0_r_valid;
  wire[1:0] NastiArbiter_1_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_1_io_master_0_r_bits_data;
  wire NastiArbiter_1_io_master_0_r_bits_last;
  wire[3:0] NastiArbiter_1_io_master_0_r_bits_id;
  wire NastiArbiter_1_io_master_0_r_bits_user;
  wire NastiArbiter_1_io_slave_aw_valid;
  wire[31:0] NastiArbiter_1_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_aw_bits_burst;
  wire NastiArbiter_1_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_region;
  wire[3:0] NastiArbiter_1_io_slave_aw_bits_id;
  wire NastiArbiter_1_io_slave_aw_bits_user;
  wire NastiArbiter_1_io_slave_w_valid;
  wire[63:0] NastiArbiter_1_io_slave_w_bits_data;
  wire NastiArbiter_1_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_1_io_slave_w_bits_strb;
  wire NastiArbiter_1_io_slave_w_bits_user;
  wire NastiArbiter_1_io_slave_b_ready;
  wire NastiArbiter_1_io_slave_ar_valid;
  wire[31:0] NastiArbiter_1_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_1_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_1_io_slave_ar_bits_burst;
  wire NastiArbiter_1_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_1_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_region;
  wire[3:0] NastiArbiter_1_io_slave_ar_bits_id;
  wire NastiArbiter_1_io_slave_ar_bits_user;
  wire NastiArbiter_1_io_slave_r_ready;
  wire NastiArbiter_2_io_master_1_aw_ready;
  wire NastiArbiter_2_io_master_1_w_ready;
  wire NastiArbiter_2_io_master_1_b_valid;
  wire[1:0] NastiArbiter_2_io_master_1_b_bits_resp;
  wire[3:0] NastiArbiter_2_io_master_1_b_bits_id;
  wire NastiArbiter_2_io_master_1_b_bits_user;
  wire NastiArbiter_2_io_master_1_ar_ready;
  wire NastiArbiter_2_io_master_1_r_valid;
  wire[1:0] NastiArbiter_2_io_master_1_r_bits_resp;
  wire[63:0] NastiArbiter_2_io_master_1_r_bits_data;
  wire NastiArbiter_2_io_master_1_r_bits_last;
  wire[3:0] NastiArbiter_2_io_master_1_r_bits_id;
  wire NastiArbiter_2_io_master_1_r_bits_user;
  wire NastiArbiter_2_io_master_0_aw_ready;
  wire NastiArbiter_2_io_master_0_w_ready;
  wire NastiArbiter_2_io_master_0_b_valid;
  wire[1:0] NastiArbiter_2_io_master_0_b_bits_resp;
  wire[3:0] NastiArbiter_2_io_master_0_b_bits_id;
  wire NastiArbiter_2_io_master_0_b_bits_user;
  wire NastiArbiter_2_io_master_0_ar_ready;
  wire NastiArbiter_2_io_master_0_r_valid;
  wire[1:0] NastiArbiter_2_io_master_0_r_bits_resp;
  wire[63:0] NastiArbiter_2_io_master_0_r_bits_data;
  wire NastiArbiter_2_io_master_0_r_bits_last;
  wire[3:0] NastiArbiter_2_io_master_0_r_bits_id;
  wire NastiArbiter_2_io_master_0_r_bits_user;
  wire NastiArbiter_2_io_slave_aw_valid;
  wire[31:0] NastiArbiter_2_io_slave_aw_bits_addr;
  wire[7:0] NastiArbiter_2_io_slave_aw_bits_len;
  wire[2:0] NastiArbiter_2_io_slave_aw_bits_size;
  wire[1:0] NastiArbiter_2_io_slave_aw_bits_burst;
  wire NastiArbiter_2_io_slave_aw_bits_lock;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_cache;
  wire[2:0] NastiArbiter_2_io_slave_aw_bits_prot;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_qos;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_region;
  wire[3:0] NastiArbiter_2_io_slave_aw_bits_id;
  wire NastiArbiter_2_io_slave_aw_bits_user;
  wire NastiArbiter_2_io_slave_w_valid;
  wire[63:0] NastiArbiter_2_io_slave_w_bits_data;
  wire NastiArbiter_2_io_slave_w_bits_last;
  wire[7:0] NastiArbiter_2_io_slave_w_bits_strb;
  wire NastiArbiter_2_io_slave_w_bits_user;
  wire NastiArbiter_2_io_slave_b_ready;
  wire NastiArbiter_2_io_slave_ar_valid;
  wire[31:0] NastiArbiter_2_io_slave_ar_bits_addr;
  wire[7:0] NastiArbiter_2_io_slave_ar_bits_len;
  wire[2:0] NastiArbiter_2_io_slave_ar_bits_size;
  wire[1:0] NastiArbiter_2_io_slave_ar_bits_burst;
  wire NastiArbiter_2_io_slave_ar_bits_lock;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_cache;
  wire[2:0] NastiArbiter_2_io_slave_ar_bits_prot;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_qos;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_region;
  wire[3:0] NastiArbiter_2_io_slave_ar_bits_id;
  wire NastiArbiter_2_io_slave_ar_bits_user;
  wire NastiArbiter_2_io_slave_r_ready;
  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[3:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[3:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_2_aw_bits_burst;
  wire NastiRouter_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_id;
  wire NastiRouter_io_slave_2_aw_bits_user;
  wire NastiRouter_io_slave_2_w_valid;
  wire[63:0] NastiRouter_io_slave_2_w_bits_data;
  wire NastiRouter_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_io_slave_2_w_bits_strb;
  wire NastiRouter_io_slave_2_w_bits_user;
  wire NastiRouter_io_slave_2_b_ready;
  wire NastiRouter_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_2_ar_bits_burst;
  wire NastiRouter_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_id;
  wire NastiRouter_io_slave_2_ar_bits_user;
  wire NastiRouter_io_slave_2_r_ready;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;
  wire NastiRouter_1_io_master_aw_ready;
  wire NastiRouter_1_io_master_w_ready;
  wire NastiRouter_1_io_master_b_valid;
  wire[1:0] NastiRouter_1_io_master_b_bits_resp;
  wire[3:0] NastiRouter_1_io_master_b_bits_id;
  wire NastiRouter_1_io_master_b_bits_user;
  wire NastiRouter_1_io_master_ar_ready;
  wire NastiRouter_1_io_master_r_valid;
  wire[1:0] NastiRouter_1_io_master_r_bits_resp;
  wire[63:0] NastiRouter_1_io_master_r_bits_data;
  wire NastiRouter_1_io_master_r_bits_last;
  wire[3:0] NastiRouter_1_io_master_r_bits_id;
  wire NastiRouter_1_io_master_r_bits_user;
  wire NastiRouter_1_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_2_aw_bits_burst;
  wire NastiRouter_1_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_region;
  wire[3:0] NastiRouter_1_io_slave_2_aw_bits_id;
  wire NastiRouter_1_io_slave_2_aw_bits_user;
  wire NastiRouter_1_io_slave_2_w_valid;
  wire[63:0] NastiRouter_1_io_slave_2_w_bits_data;
  wire NastiRouter_1_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_2_w_bits_strb;
  wire NastiRouter_1_io_slave_2_w_bits_user;
  wire NastiRouter_1_io_slave_2_b_ready;
  wire NastiRouter_1_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_2_ar_bits_burst;
  wire NastiRouter_1_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_region;
  wire[3:0] NastiRouter_1_io_slave_2_ar_bits_id;
  wire NastiRouter_1_io_slave_2_ar_bits_user;
  wire NastiRouter_1_io_slave_2_r_ready;
  wire NastiRouter_1_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_aw_bits_burst;
  wire NastiRouter_1_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_region;
  wire[3:0] NastiRouter_1_io_slave_1_aw_bits_id;
  wire NastiRouter_1_io_slave_1_aw_bits_user;
  wire NastiRouter_1_io_slave_1_w_valid;
  wire[63:0] NastiRouter_1_io_slave_1_w_bits_data;
  wire NastiRouter_1_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_1_w_bits_strb;
  wire NastiRouter_1_io_slave_1_w_bits_user;
  wire NastiRouter_1_io_slave_1_b_ready;
  wire NastiRouter_1_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_1_ar_bits_burst;
  wire NastiRouter_1_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_region;
  wire[3:0] NastiRouter_1_io_slave_1_ar_bits_id;
  wire NastiRouter_1_io_slave_1_ar_bits_user;
  wire NastiRouter_1_io_slave_1_r_ready;
  wire NastiRouter_1_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_1_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_aw_bits_burst;
  wire NastiRouter_1_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_region;
  wire[3:0] NastiRouter_1_io_slave_0_aw_bits_id;
  wire NastiRouter_1_io_slave_0_aw_bits_user;
  wire NastiRouter_1_io_slave_0_w_valid;
  wire[63:0] NastiRouter_1_io_slave_0_w_bits_data;
  wire NastiRouter_1_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_1_io_slave_0_w_bits_strb;
  wire NastiRouter_1_io_slave_0_w_bits_user;
  wire NastiRouter_1_io_slave_0_b_ready;
  wire NastiRouter_1_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_1_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_1_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_1_io_slave_0_ar_bits_burst;
  wire NastiRouter_1_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_1_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_region;
  wire[3:0] NastiRouter_1_io_slave_0_ar_bits_id;
  wire NastiRouter_1_io_slave_0_ar_bits_user;
  wire NastiRouter_1_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiArbiter_io_slave_r_ready;
  assign io_slaves_0_ar_bits_user = NastiArbiter_io_slave_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiArbiter_io_slave_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiArbiter_io_slave_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiArbiter_io_slave_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiArbiter_io_slave_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiArbiter_io_slave_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiArbiter_io_slave_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiArbiter_io_slave_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiArbiter_io_slave_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiArbiter_io_slave_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiArbiter_io_slave_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiArbiter_io_slave_ar_valid;
  assign io_slaves_0_b_ready = NastiArbiter_io_slave_b_ready;
  assign io_slaves_0_w_bits_user = NastiArbiter_io_slave_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiArbiter_io_slave_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiArbiter_io_slave_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiArbiter_io_slave_w_bits_data;
  assign io_slaves_0_w_valid = NastiArbiter_io_slave_w_valid;
  assign io_slaves_0_aw_bits_user = NastiArbiter_io_slave_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiArbiter_io_slave_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiArbiter_io_slave_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiArbiter_io_slave_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiArbiter_io_slave_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiArbiter_io_slave_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiArbiter_io_slave_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiArbiter_io_slave_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiArbiter_io_slave_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiArbiter_io_slave_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiArbiter_io_slave_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiArbiter_io_slave_aw_valid;
  assign io_slaves_1_r_ready = NastiArbiter_1_io_slave_r_ready;
  assign io_slaves_1_ar_bits_user = NastiArbiter_1_io_slave_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiArbiter_1_io_slave_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiArbiter_1_io_slave_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiArbiter_1_io_slave_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiArbiter_1_io_slave_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiArbiter_1_io_slave_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiArbiter_1_io_slave_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiArbiter_1_io_slave_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiArbiter_1_io_slave_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiArbiter_1_io_slave_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiArbiter_1_io_slave_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiArbiter_1_io_slave_ar_valid;
  assign io_slaves_1_b_ready = NastiArbiter_1_io_slave_b_ready;
  assign io_slaves_1_w_bits_user = NastiArbiter_1_io_slave_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiArbiter_1_io_slave_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiArbiter_1_io_slave_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiArbiter_1_io_slave_w_bits_data;
  assign io_slaves_1_w_valid = NastiArbiter_1_io_slave_w_valid;
  assign io_slaves_1_aw_bits_user = NastiArbiter_1_io_slave_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiArbiter_1_io_slave_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiArbiter_1_io_slave_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiArbiter_1_io_slave_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiArbiter_1_io_slave_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiArbiter_1_io_slave_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiArbiter_1_io_slave_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiArbiter_1_io_slave_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiArbiter_1_io_slave_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiArbiter_1_io_slave_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiArbiter_1_io_slave_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiArbiter_1_io_slave_aw_valid;
  assign io_slaves_2_r_ready = NastiArbiter_2_io_slave_r_ready;
  assign io_slaves_2_ar_bits_user = NastiArbiter_2_io_slave_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiArbiter_2_io_slave_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiArbiter_2_io_slave_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiArbiter_2_io_slave_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiArbiter_2_io_slave_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiArbiter_2_io_slave_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiArbiter_2_io_slave_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiArbiter_2_io_slave_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiArbiter_2_io_slave_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiArbiter_2_io_slave_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiArbiter_2_io_slave_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiArbiter_2_io_slave_ar_valid;
  assign io_slaves_2_b_ready = NastiArbiter_2_io_slave_b_ready;
  assign io_slaves_2_w_bits_user = NastiArbiter_2_io_slave_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiArbiter_2_io_slave_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiArbiter_2_io_slave_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiArbiter_2_io_slave_w_bits_data;
  assign io_slaves_2_w_valid = NastiArbiter_2_io_slave_w_valid;
  assign io_slaves_2_aw_bits_user = NastiArbiter_2_io_slave_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiArbiter_2_io_slave_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiArbiter_2_io_slave_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiArbiter_2_io_slave_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiArbiter_2_io_slave_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiArbiter_2_io_slave_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiArbiter_2_io_slave_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiArbiter_2_io_slave_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiArbiter_2_io_slave_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiArbiter_2_io_slave_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiArbiter_2_io_slave_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiArbiter_2_io_slave_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  assign io_masters_1_r_bits_user = NastiRouter_1_io_master_r_bits_user;
  assign io_masters_1_r_bits_id = NastiRouter_1_io_master_r_bits_id;
  assign io_masters_1_r_bits_last = NastiRouter_1_io_master_r_bits_last;
  assign io_masters_1_r_bits_data = NastiRouter_1_io_master_r_bits_data;
  assign io_masters_1_r_bits_resp = NastiRouter_1_io_master_r_bits_resp;
  assign io_masters_1_r_valid = NastiRouter_1_io_master_r_valid;
  assign io_masters_1_ar_ready = NastiRouter_1_io_master_ar_ready;
  assign io_masters_1_b_bits_user = NastiRouter_1_io_master_b_bits_user;
  assign io_masters_1_b_bits_id = NastiRouter_1_io_master_b_bits_id;
  assign io_masters_1_b_bits_resp = NastiRouter_1_io_master_b_bits_resp;
  assign io_masters_1_b_valid = NastiRouter_1_io_master_b_valid;
  assign io_masters_1_w_ready = NastiRouter_1_io_master_w_ready;
  assign io_masters_1_aw_ready = NastiRouter_1_io_master_aw_ready;
  NastiRouter_0 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_2_aw_ready( NastiArbiter_2_io_master_0_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( NastiArbiter_2_io_master_0_w_ready ),
       .io_slave_2_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_slave_2_b_valid( NastiArbiter_2_io_master_0_b_valid ),
       .io_slave_2_b_bits_resp( NastiArbiter_2_io_master_0_b_bits_resp ),
       .io_slave_2_b_bits_id( NastiArbiter_2_io_master_0_b_bits_id ),
       .io_slave_2_b_bits_user( NastiArbiter_2_io_master_0_b_bits_user ),
       .io_slave_2_ar_ready( NastiArbiter_2_io_master_0_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_slave_2_r_valid( NastiArbiter_2_io_master_0_r_valid ),
       .io_slave_2_r_bits_resp( NastiArbiter_2_io_master_0_r_bits_resp ),
       .io_slave_2_r_bits_data( NastiArbiter_2_io_master_0_r_bits_data ),
       .io_slave_2_r_bits_last( NastiArbiter_2_io_master_0_r_bits_last ),
       .io_slave_2_r_bits_id( NastiArbiter_2_io_master_0_r_bits_id ),
       .io_slave_2_r_bits_user( NastiArbiter_2_io_master_0_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user )
  );
  NastiRouter_0 NastiRouter_1(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_1_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_1_aw_valid ),
       .io_master_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_master_w_ready( NastiRouter_1_io_master_w_ready ),
       .io_master_w_valid( io_masters_1_w_valid ),
       .io_master_w_bits_data( io_masters_1_w_bits_data ),
       .io_master_w_bits_last( io_masters_1_w_bits_last ),
       .io_master_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_master_w_bits_user( io_masters_1_w_bits_user ),
       .io_master_b_ready( io_masters_1_b_ready ),
       .io_master_b_valid( NastiRouter_1_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_1_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_1_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_1_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_1_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_1_ar_valid ),
       .io_master_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_master_r_ready( io_masters_1_r_ready ),
       .io_master_r_valid( NastiRouter_1_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_1_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_1_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_1_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_1_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_1_io_master_r_bits_user ),
       .io_slave_2_aw_ready( NastiArbiter_2_io_master_1_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_1_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_1_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_1_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_1_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_1_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_1_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_1_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_1_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_1_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_1_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_1_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_1_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( NastiArbiter_2_io_master_1_w_ready ),
       .io_slave_2_w_valid( NastiRouter_1_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_1_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_1_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_1_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_1_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_1_io_slave_2_b_ready ),
       .io_slave_2_b_valid( NastiArbiter_2_io_master_1_b_valid ),
       .io_slave_2_b_bits_resp( NastiArbiter_2_io_master_1_b_bits_resp ),
       .io_slave_2_b_bits_id( NastiArbiter_2_io_master_1_b_bits_id ),
       .io_slave_2_b_bits_user( NastiArbiter_2_io_master_1_b_bits_user ),
       .io_slave_2_ar_ready( NastiArbiter_2_io_master_1_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_1_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_1_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_1_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_1_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_1_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_1_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_1_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_1_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_1_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_1_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_1_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_1_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_1_io_slave_2_r_ready ),
       .io_slave_2_r_valid( NastiArbiter_2_io_master_1_r_valid ),
       .io_slave_2_r_bits_resp( NastiArbiter_2_io_master_1_r_bits_resp ),
       .io_slave_2_r_bits_data( NastiArbiter_2_io_master_1_r_bits_data ),
       .io_slave_2_r_bits_last( NastiArbiter_2_io_master_1_r_bits_last ),
       .io_slave_2_r_bits_id( NastiArbiter_2_io_master_1_r_bits_id ),
       .io_slave_2_r_bits_user( NastiArbiter_2_io_master_1_r_bits_user ),
       .io_slave_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_slave_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_slave_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_slave_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_slave_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_slave_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_slave_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_slave_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_slave_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_slave_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_slave_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_slave_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_slave_0_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_slave_0_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_slave_0_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_slave_0_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_slave_0_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_slave_0_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_slave_0_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_slave_0_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_slave_0_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_slave_0_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_slave_0_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_slave_0_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_slave_0_r_bits_user( NastiArbiter_io_master_1_r_bits_user )
  );
  NastiArbiter NastiArbiter(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_0_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_0_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_0_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_0_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_0_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_0_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_0_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_0_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_0_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_0_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_0_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_0_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_0_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_0_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_0_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_0_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_0_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_0_b_ready ),
       .io_master_1_b_valid( NastiArbiter_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_0_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_0_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_0_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_0_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_0_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_0_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_0_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_0_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_0_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_0_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_0_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_0_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_0_r_ready ),
       .io_master_1_r_valid( NastiArbiter_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_master_0_b_valid( NastiArbiter_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_master_0_r_valid( NastiArbiter_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_0_w_ready ),
       .io_slave_w_valid( NastiArbiter_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_0_b_valid ),
       .io_slave_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_0_r_valid ),
       .io_slave_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiArbiter NastiArbiter_1(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_1_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_1_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_1_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_1_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_1_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_1_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_1_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_1_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_1_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_1_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_1_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_1_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_1_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_1_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_1_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_1_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_1_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_1_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_1_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_1_b_ready ),
       .io_master_1_b_valid( NastiArbiter_1_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_1_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_1_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_1_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_1_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_1_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_1_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_1_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_1_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_1_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_1_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_1_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_1_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_1_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_1_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_1_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_1_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_1_r_ready ),
       .io_master_1_r_valid( NastiArbiter_1_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_1_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_1_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_1_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_1_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_1_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_1_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_1_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_master_0_b_valid( NastiArbiter_1_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_1_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_1_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_1_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_1_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_master_0_r_valid( NastiArbiter_1_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_1_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_1_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_1_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_1_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_1_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_1_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_1_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_1_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_1_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_1_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_1_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_1_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_1_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_1_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_1_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_1_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_1_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_1_w_ready ),
       .io_slave_w_valid( NastiArbiter_1_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_1_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_1_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_1_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_1_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_1_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_1_b_valid ),
       .io_slave_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_1_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_1_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_1_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_1_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_1_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_1_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_1_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_1_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_1_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_1_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_1_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_1_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_1_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_1_r_valid ),
       .io_slave_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_1_r_bits_user )
  );
  NastiArbiter NastiArbiter_2(.clk(clk), .reset(reset),
       .io_master_1_aw_ready( NastiArbiter_2_io_master_1_aw_ready ),
       .io_master_1_aw_valid( NastiRouter_1_io_slave_2_aw_valid ),
       .io_master_1_aw_bits_addr( NastiRouter_1_io_slave_2_aw_bits_addr ),
       .io_master_1_aw_bits_len( NastiRouter_1_io_slave_2_aw_bits_len ),
       .io_master_1_aw_bits_size( NastiRouter_1_io_slave_2_aw_bits_size ),
       .io_master_1_aw_bits_burst( NastiRouter_1_io_slave_2_aw_bits_burst ),
       .io_master_1_aw_bits_lock( NastiRouter_1_io_slave_2_aw_bits_lock ),
       .io_master_1_aw_bits_cache( NastiRouter_1_io_slave_2_aw_bits_cache ),
       .io_master_1_aw_bits_prot( NastiRouter_1_io_slave_2_aw_bits_prot ),
       .io_master_1_aw_bits_qos( NastiRouter_1_io_slave_2_aw_bits_qos ),
       .io_master_1_aw_bits_region( NastiRouter_1_io_slave_2_aw_bits_region ),
       .io_master_1_aw_bits_id( NastiRouter_1_io_slave_2_aw_bits_id ),
       .io_master_1_aw_bits_user( NastiRouter_1_io_slave_2_aw_bits_user ),
       .io_master_1_w_ready( NastiArbiter_2_io_master_1_w_ready ),
       .io_master_1_w_valid( NastiRouter_1_io_slave_2_w_valid ),
       .io_master_1_w_bits_data( NastiRouter_1_io_slave_2_w_bits_data ),
       .io_master_1_w_bits_last( NastiRouter_1_io_slave_2_w_bits_last ),
       .io_master_1_w_bits_strb( NastiRouter_1_io_slave_2_w_bits_strb ),
       .io_master_1_w_bits_user( NastiRouter_1_io_slave_2_w_bits_user ),
       .io_master_1_b_ready( NastiRouter_1_io_slave_2_b_ready ),
       .io_master_1_b_valid( NastiArbiter_2_io_master_1_b_valid ),
       .io_master_1_b_bits_resp( NastiArbiter_2_io_master_1_b_bits_resp ),
       .io_master_1_b_bits_id( NastiArbiter_2_io_master_1_b_bits_id ),
       .io_master_1_b_bits_user( NastiArbiter_2_io_master_1_b_bits_user ),
       .io_master_1_ar_ready( NastiArbiter_2_io_master_1_ar_ready ),
       .io_master_1_ar_valid( NastiRouter_1_io_slave_2_ar_valid ),
       .io_master_1_ar_bits_addr( NastiRouter_1_io_slave_2_ar_bits_addr ),
       .io_master_1_ar_bits_len( NastiRouter_1_io_slave_2_ar_bits_len ),
       .io_master_1_ar_bits_size( NastiRouter_1_io_slave_2_ar_bits_size ),
       .io_master_1_ar_bits_burst( NastiRouter_1_io_slave_2_ar_bits_burst ),
       .io_master_1_ar_bits_lock( NastiRouter_1_io_slave_2_ar_bits_lock ),
       .io_master_1_ar_bits_cache( NastiRouter_1_io_slave_2_ar_bits_cache ),
       .io_master_1_ar_bits_prot( NastiRouter_1_io_slave_2_ar_bits_prot ),
       .io_master_1_ar_bits_qos( NastiRouter_1_io_slave_2_ar_bits_qos ),
       .io_master_1_ar_bits_region( NastiRouter_1_io_slave_2_ar_bits_region ),
       .io_master_1_ar_bits_id( NastiRouter_1_io_slave_2_ar_bits_id ),
       .io_master_1_ar_bits_user( NastiRouter_1_io_slave_2_ar_bits_user ),
       .io_master_1_r_ready( NastiRouter_1_io_slave_2_r_ready ),
       .io_master_1_r_valid( NastiArbiter_2_io_master_1_r_valid ),
       .io_master_1_r_bits_resp( NastiArbiter_2_io_master_1_r_bits_resp ),
       .io_master_1_r_bits_data( NastiArbiter_2_io_master_1_r_bits_data ),
       .io_master_1_r_bits_last( NastiArbiter_2_io_master_1_r_bits_last ),
       .io_master_1_r_bits_id( NastiArbiter_2_io_master_1_r_bits_id ),
       .io_master_1_r_bits_user( NastiArbiter_2_io_master_1_r_bits_user ),
       .io_master_0_aw_ready( NastiArbiter_2_io_master_0_aw_ready ),
       .io_master_0_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_master_0_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_master_0_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_master_0_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_master_0_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_master_0_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_master_0_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_master_0_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_master_0_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_master_0_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_master_0_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_master_0_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_master_0_w_ready( NastiArbiter_2_io_master_0_w_ready ),
       .io_master_0_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_master_0_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_master_0_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_master_0_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_master_0_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_master_0_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_master_0_b_valid( NastiArbiter_2_io_master_0_b_valid ),
       .io_master_0_b_bits_resp( NastiArbiter_2_io_master_0_b_bits_resp ),
       .io_master_0_b_bits_id( NastiArbiter_2_io_master_0_b_bits_id ),
       .io_master_0_b_bits_user( NastiArbiter_2_io_master_0_b_bits_user ),
       .io_master_0_ar_ready( NastiArbiter_2_io_master_0_ar_ready ),
       .io_master_0_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_master_0_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_master_0_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_master_0_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_master_0_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_master_0_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_master_0_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_master_0_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_master_0_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_master_0_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_master_0_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_master_0_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_master_0_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_master_0_r_valid( NastiArbiter_2_io_master_0_r_valid ),
       .io_master_0_r_bits_resp( NastiArbiter_2_io_master_0_r_bits_resp ),
       .io_master_0_r_bits_data( NastiArbiter_2_io_master_0_r_bits_data ),
       .io_master_0_r_bits_last( NastiArbiter_2_io_master_0_r_bits_last ),
       .io_master_0_r_bits_id( NastiArbiter_2_io_master_0_r_bits_id ),
       .io_master_0_r_bits_user( NastiArbiter_2_io_master_0_r_bits_user ),
       .io_slave_aw_ready( io_slaves_2_aw_ready ),
       .io_slave_aw_valid( NastiArbiter_2_io_slave_aw_valid ),
       .io_slave_aw_bits_addr( NastiArbiter_2_io_slave_aw_bits_addr ),
       .io_slave_aw_bits_len( NastiArbiter_2_io_slave_aw_bits_len ),
       .io_slave_aw_bits_size( NastiArbiter_2_io_slave_aw_bits_size ),
       .io_slave_aw_bits_burst( NastiArbiter_2_io_slave_aw_bits_burst ),
       .io_slave_aw_bits_lock( NastiArbiter_2_io_slave_aw_bits_lock ),
       .io_slave_aw_bits_cache( NastiArbiter_2_io_slave_aw_bits_cache ),
       .io_slave_aw_bits_prot( NastiArbiter_2_io_slave_aw_bits_prot ),
       .io_slave_aw_bits_qos( NastiArbiter_2_io_slave_aw_bits_qos ),
       .io_slave_aw_bits_region( NastiArbiter_2_io_slave_aw_bits_region ),
       .io_slave_aw_bits_id( NastiArbiter_2_io_slave_aw_bits_id ),
       .io_slave_aw_bits_user( NastiArbiter_2_io_slave_aw_bits_user ),
       .io_slave_w_ready( io_slaves_2_w_ready ),
       .io_slave_w_valid( NastiArbiter_2_io_slave_w_valid ),
       .io_slave_w_bits_data( NastiArbiter_2_io_slave_w_bits_data ),
       .io_slave_w_bits_last( NastiArbiter_2_io_slave_w_bits_last ),
       .io_slave_w_bits_strb( NastiArbiter_2_io_slave_w_bits_strb ),
       .io_slave_w_bits_user( NastiArbiter_2_io_slave_w_bits_user ),
       .io_slave_b_ready( NastiArbiter_2_io_slave_b_ready ),
       .io_slave_b_valid( io_slaves_2_b_valid ),
       .io_slave_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slave_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slave_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slave_ar_ready( io_slaves_2_ar_ready ),
       .io_slave_ar_valid( NastiArbiter_2_io_slave_ar_valid ),
       .io_slave_ar_bits_addr( NastiArbiter_2_io_slave_ar_bits_addr ),
       .io_slave_ar_bits_len( NastiArbiter_2_io_slave_ar_bits_len ),
       .io_slave_ar_bits_size( NastiArbiter_2_io_slave_ar_bits_size ),
       .io_slave_ar_bits_burst( NastiArbiter_2_io_slave_ar_bits_burst ),
       .io_slave_ar_bits_lock( NastiArbiter_2_io_slave_ar_bits_lock ),
       .io_slave_ar_bits_cache( NastiArbiter_2_io_slave_ar_bits_cache ),
       .io_slave_ar_bits_prot( NastiArbiter_2_io_slave_ar_bits_prot ),
       .io_slave_ar_bits_qos( NastiArbiter_2_io_slave_ar_bits_qos ),
       .io_slave_ar_bits_region( NastiArbiter_2_io_slave_ar_bits_region ),
       .io_slave_ar_bits_id( NastiArbiter_2_io_slave_ar_bits_id ),
       .io_slave_ar_bits_user( NastiArbiter_2_io_slave_ar_bits_user ),
       .io_slave_r_ready( NastiArbiter_2_io_slave_r_ready ),
       .io_slave_r_valid( io_slaves_2_r_valid ),
       .io_slave_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slave_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slave_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slave_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slave_r_bits_user( io_slaves_2_r_bits_user )
  );
endmodule

module NastiRouter_1(input clk, input reset,
    output io_master_aw_ready,
    input  io_master_aw_valid,
    input [31:0] io_master_aw_bits_addr,
    input [7:0] io_master_aw_bits_len,
    input [2:0] io_master_aw_bits_size,
    input [1:0] io_master_aw_bits_burst,
    input  io_master_aw_bits_lock,
    input [3:0] io_master_aw_bits_cache,
    input [2:0] io_master_aw_bits_prot,
    input [3:0] io_master_aw_bits_qos,
    input [3:0] io_master_aw_bits_region,
    input [3:0] io_master_aw_bits_id,
    input  io_master_aw_bits_user,
    output io_master_w_ready,
    input  io_master_w_valid,
    input [63:0] io_master_w_bits_data,
    input  io_master_w_bits_last,
    input [7:0] io_master_w_bits_strb,
    input  io_master_w_bits_user,
    input  io_master_b_ready,
    output io_master_b_valid,
    output[1:0] io_master_b_bits_resp,
    output[3:0] io_master_b_bits_id,
    output io_master_b_bits_user,
    output io_master_ar_ready,
    input  io_master_ar_valid,
    input [31:0] io_master_ar_bits_addr,
    input [7:0] io_master_ar_bits_len,
    input [2:0] io_master_ar_bits_size,
    input [1:0] io_master_ar_bits_burst,
    input  io_master_ar_bits_lock,
    input [3:0] io_master_ar_bits_cache,
    input [2:0] io_master_ar_bits_prot,
    input [3:0] io_master_ar_bits_qos,
    input [3:0] io_master_ar_bits_region,
    input [3:0] io_master_ar_bits_id,
    input  io_master_ar_bits_user,
    input  io_master_r_ready,
    output io_master_r_valid,
    output[1:0] io_master_r_bits_resp,
    output[63:0] io_master_r_bits_data,
    output io_master_r_bits_last,
    output[3:0] io_master_r_bits_id,
    output io_master_r_bits_user,
    input  io_slave_2_aw_ready,
    output io_slave_2_aw_valid,
    output[31:0] io_slave_2_aw_bits_addr,
    output[7:0] io_slave_2_aw_bits_len,
    output[2:0] io_slave_2_aw_bits_size,
    output[1:0] io_slave_2_aw_bits_burst,
    output io_slave_2_aw_bits_lock,
    output[3:0] io_slave_2_aw_bits_cache,
    output[2:0] io_slave_2_aw_bits_prot,
    output[3:0] io_slave_2_aw_bits_qos,
    output[3:0] io_slave_2_aw_bits_region,
    output[3:0] io_slave_2_aw_bits_id,
    output io_slave_2_aw_bits_user,
    input  io_slave_2_w_ready,
    output io_slave_2_w_valid,
    output[63:0] io_slave_2_w_bits_data,
    output io_slave_2_w_bits_last,
    output[7:0] io_slave_2_w_bits_strb,
    output io_slave_2_w_bits_user,
    output io_slave_2_b_ready,
    input  io_slave_2_b_valid,
    input [1:0] io_slave_2_b_bits_resp,
    input [3:0] io_slave_2_b_bits_id,
    input  io_slave_2_b_bits_user,
    input  io_slave_2_ar_ready,
    output io_slave_2_ar_valid,
    output[31:0] io_slave_2_ar_bits_addr,
    output[7:0] io_slave_2_ar_bits_len,
    output[2:0] io_slave_2_ar_bits_size,
    output[1:0] io_slave_2_ar_bits_burst,
    output io_slave_2_ar_bits_lock,
    output[3:0] io_slave_2_ar_bits_cache,
    output[2:0] io_slave_2_ar_bits_prot,
    output[3:0] io_slave_2_ar_bits_qos,
    output[3:0] io_slave_2_ar_bits_region,
    output[3:0] io_slave_2_ar_bits_id,
    output io_slave_2_ar_bits_user,
    output io_slave_2_r_ready,
    input  io_slave_2_r_valid,
    input [1:0] io_slave_2_r_bits_resp,
    input [63:0] io_slave_2_r_bits_data,
    input  io_slave_2_r_bits_last,
    input [3:0] io_slave_2_r_bits_id,
    input  io_slave_2_r_bits_user,
    input  io_slave_1_aw_ready,
    output io_slave_1_aw_valid,
    output[31:0] io_slave_1_aw_bits_addr,
    output[7:0] io_slave_1_aw_bits_len,
    output[2:0] io_slave_1_aw_bits_size,
    output[1:0] io_slave_1_aw_bits_burst,
    output io_slave_1_aw_bits_lock,
    output[3:0] io_slave_1_aw_bits_cache,
    output[2:0] io_slave_1_aw_bits_prot,
    output[3:0] io_slave_1_aw_bits_qos,
    output[3:0] io_slave_1_aw_bits_region,
    output[3:0] io_slave_1_aw_bits_id,
    output io_slave_1_aw_bits_user,
    input  io_slave_1_w_ready,
    output io_slave_1_w_valid,
    output[63:0] io_slave_1_w_bits_data,
    output io_slave_1_w_bits_last,
    output[7:0] io_slave_1_w_bits_strb,
    output io_slave_1_w_bits_user,
    output io_slave_1_b_ready,
    input  io_slave_1_b_valid,
    input [1:0] io_slave_1_b_bits_resp,
    input [3:0] io_slave_1_b_bits_id,
    input  io_slave_1_b_bits_user,
    input  io_slave_1_ar_ready,
    output io_slave_1_ar_valid,
    output[31:0] io_slave_1_ar_bits_addr,
    output[7:0] io_slave_1_ar_bits_len,
    output[2:0] io_slave_1_ar_bits_size,
    output[1:0] io_slave_1_ar_bits_burst,
    output io_slave_1_ar_bits_lock,
    output[3:0] io_slave_1_ar_bits_cache,
    output[2:0] io_slave_1_ar_bits_prot,
    output[3:0] io_slave_1_ar_bits_qos,
    output[3:0] io_slave_1_ar_bits_region,
    output[3:0] io_slave_1_ar_bits_id,
    output io_slave_1_ar_bits_user,
    output io_slave_1_r_ready,
    input  io_slave_1_r_valid,
    input [1:0] io_slave_1_r_bits_resp,
    input [63:0] io_slave_1_r_bits_data,
    input  io_slave_1_r_bits_last,
    input [3:0] io_slave_1_r_bits_id,
    input  io_slave_1_r_bits_user,
    input  io_slave_0_aw_ready,
    output io_slave_0_aw_valid,
    output[31:0] io_slave_0_aw_bits_addr,
    output[7:0] io_slave_0_aw_bits_len,
    output[2:0] io_slave_0_aw_bits_size,
    output[1:0] io_slave_0_aw_bits_burst,
    output io_slave_0_aw_bits_lock,
    output[3:0] io_slave_0_aw_bits_cache,
    output[2:0] io_slave_0_aw_bits_prot,
    output[3:0] io_slave_0_aw_bits_qos,
    output[3:0] io_slave_0_aw_bits_region,
    output[3:0] io_slave_0_aw_bits_id,
    output io_slave_0_aw_bits_user,
    input  io_slave_0_w_ready,
    output io_slave_0_w_valid,
    output[63:0] io_slave_0_w_bits_data,
    output io_slave_0_w_bits_last,
    output[7:0] io_slave_0_w_bits_strb,
    output io_slave_0_w_bits_user,
    output io_slave_0_b_ready,
    input  io_slave_0_b_valid,
    input [1:0] io_slave_0_b_bits_resp,
    input [3:0] io_slave_0_b_bits_id,
    input  io_slave_0_b_bits_user,
    input  io_slave_0_ar_ready,
    output io_slave_0_ar_valid,
    output[31:0] io_slave_0_ar_bits_addr,
    output[7:0] io_slave_0_ar_bits_len,
    output[2:0] io_slave_0_ar_bits_size,
    output[1:0] io_slave_0_ar_bits_burst,
    output io_slave_0_ar_bits_lock,
    output[3:0] io_slave_0_ar_bits_cache,
    output[2:0] io_slave_0_ar_bits_prot,
    output[3:0] io_slave_0_ar_bits_qos,
    output[3:0] io_slave_0_ar_bits_region,
    output[3:0] io_slave_0_ar_bits_id,
    output io_slave_0_ar_bits_user,
    output io_slave_0_r_ready,
    input  io_slave_0_r_valid,
    input [1:0] io_slave_0_r_bits_resp,
    input [63:0] io_slave_0_r_bits_data,
    input  io_slave_0_r_bits_last,
    input [3:0] io_slave_0_r_bits_id,
    input  io_slave_0_r_bits_user
);

  wire T0;
  wire r_invalid;
  wire T1;
  wire[2:0] ar_route;
  wire[2:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire w_invalid;
  wire T14;
  wire[2:0] aw_route;
  wire[2:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  reg  R29;
  wire T82;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  reg  R40;
  wire T83;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  reg  R51;
  wire T84;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire ar_ready;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire w_ready;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire aw_ready;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire b_arb_io_in_3_ready;
  wire b_arb_io_in_2_ready;
  wire b_arb_io_in_1_ready;
  wire b_arb_io_in_0_ready;
  wire b_arb_io_out_valid;
  wire[1:0] b_arb_io_out_bits_resp;
  wire[3:0] b_arb_io_out_bits_id;
  wire b_arb_io_out_bits_user;
  wire r_arb_io_in_3_ready;
  wire r_arb_io_in_2_ready;
  wire r_arb_io_in_1_ready;
  wire r_arb_io_in_0_ready;
  wire r_arb_io_out_valid;
  wire[1:0] r_arb_io_out_bits_resp;
  wire[63:0] r_arb_io_out_bits_data;
  wire r_arb_io_out_bits_last;
  wire[3:0] r_arb_io_out_bits_id;
  wire r_arb_io_out_bits_user;
  wire err_slave_io_aw_ready;
  wire err_slave_io_w_ready;
  wire err_slave_io_b_valid;
  wire[1:0] err_slave_io_b_bits_resp;
  wire[3:0] err_slave_io_b_bits_id;
  wire err_slave_io_ar_ready;
  wire err_slave_io_r_valid;
  wire[1:0] err_slave_io_r_bits_resp;
  wire[63:0] err_slave_io_r_bits_data;
  wire err_slave_io_r_bits_last;
  wire[3:0] err_slave_io_r_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R29 = {1{$random}};
    R40 = {1{$random}};
    R51 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = r_invalid & io_master_ar_valid;
  assign r_invalid = T1 ^ 1'h1;
  assign T1 = ar_route != 3'h0;
  assign ar_route = T2;
  assign T2 = {T10, T3};
  assign T3 = {T7, T4};
  assign T4 = T6 & T5;
  assign T5 = io_master_ar_bits_addr < 32'h40008000;
  assign T6 = 32'h40000000 <= io_master_ar_bits_addr;
  assign T7 = T9 & T8;
  assign T8 = io_master_ar_bits_addr < 32'h40010000;
  assign T9 = 32'h40008000 <= io_master_ar_bits_addr;
  assign T10 = T12 & T11;
  assign T11 = io_master_ar_bits_addr < 32'h40010200;
  assign T12 = 32'h40010000 <= io_master_ar_bits_addr;
  assign T13 = w_invalid & io_master_aw_valid;
  assign w_invalid = T14 ^ 1'h1;
  assign T14 = aw_route != 3'h0;
  assign aw_route = T15;
  assign T15 = {T23, T16};
  assign T16 = {T20, T17};
  assign T17 = T19 & T18;
  assign T18 = io_master_aw_bits_addr < 32'h40008000;
  assign T19 = 32'h40000000 <= io_master_aw_bits_addr;
  assign T20 = T22 & T21;
  assign T21 = io_master_aw_bits_addr < 32'h40010000;
  assign T22 = 32'h40008000 <= io_master_aw_bits_addr;
  assign T23 = T25 & T24;
  assign T24 = io_master_aw_bits_addr < 32'h40010200;
  assign T25 = 32'h40010000 <= io_master_aw_bits_addr;
  assign io_slave_0_r_ready = r_arb_io_in_0_ready;
  assign io_slave_0_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_0_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_0_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_0_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_0_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_0_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_0_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_0_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_0_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_0_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_0_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_0_ar_valid = T26;
  assign T26 = io_master_ar_valid & T27;
  assign T27 = ar_route[1'h0:1'h0];
  assign io_slave_0_b_ready = b_arb_io_in_0_ready;
  assign io_slave_0_w_bits_user = io_master_w_bits_user;
  assign io_slave_0_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_0_w_bits_last = io_master_w_bits_last;
  assign io_slave_0_w_bits_data = io_master_w_bits_data;
  assign io_slave_0_w_valid = T28;
  assign T28 = io_master_w_valid & R29;
  assign T82 = reset ? 1'h0 : T30;
  assign T30 = T33 ? 1'h0 : T31;
  assign T31 = T32 ? 1'h1 : R29;
  assign T32 = io_slave_0_aw_ready & io_slave_0_aw_valid;
  assign T33 = T34 & io_slave_0_w_bits_last;
  assign T34 = io_slave_0_w_ready & io_slave_0_w_valid;
  assign io_slave_0_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_0_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_0_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_0_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_0_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_0_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_0_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_0_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_0_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_0_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_0_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_0_aw_valid = T35;
  assign T35 = io_master_aw_valid & T36;
  assign T36 = aw_route[1'h0:1'h0];
  assign io_slave_1_r_ready = r_arb_io_in_1_ready;
  assign io_slave_1_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_1_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_1_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_1_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_1_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_1_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_1_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_1_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_1_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_1_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_1_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_1_ar_valid = T37;
  assign T37 = io_master_ar_valid & T38;
  assign T38 = ar_route[1'h1:1'h1];
  assign io_slave_1_b_ready = b_arb_io_in_1_ready;
  assign io_slave_1_w_bits_user = io_master_w_bits_user;
  assign io_slave_1_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_1_w_bits_last = io_master_w_bits_last;
  assign io_slave_1_w_bits_data = io_master_w_bits_data;
  assign io_slave_1_w_valid = T39;
  assign T39 = io_master_w_valid & R40;
  assign T83 = reset ? 1'h0 : T41;
  assign T41 = T44 ? 1'h0 : T42;
  assign T42 = T43 ? 1'h1 : R40;
  assign T43 = io_slave_1_aw_ready & io_slave_1_aw_valid;
  assign T44 = T45 & io_slave_1_w_bits_last;
  assign T45 = io_slave_1_w_ready & io_slave_1_w_valid;
  assign io_slave_1_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_1_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_1_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_1_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_1_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_1_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_1_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_1_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_1_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_1_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_1_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_1_aw_valid = T46;
  assign T46 = io_master_aw_valid & T47;
  assign T47 = aw_route[1'h1:1'h1];
  assign io_slave_2_r_ready = r_arb_io_in_2_ready;
  assign io_slave_2_ar_bits_user = io_master_ar_bits_user;
  assign io_slave_2_ar_bits_id = io_master_ar_bits_id;
  assign io_slave_2_ar_bits_region = io_master_ar_bits_region;
  assign io_slave_2_ar_bits_qos = io_master_ar_bits_qos;
  assign io_slave_2_ar_bits_prot = io_master_ar_bits_prot;
  assign io_slave_2_ar_bits_cache = io_master_ar_bits_cache;
  assign io_slave_2_ar_bits_lock = io_master_ar_bits_lock;
  assign io_slave_2_ar_bits_burst = io_master_ar_bits_burst;
  assign io_slave_2_ar_bits_size = io_master_ar_bits_size;
  assign io_slave_2_ar_bits_len = io_master_ar_bits_len;
  assign io_slave_2_ar_bits_addr = io_master_ar_bits_addr;
  assign io_slave_2_ar_valid = T48;
  assign T48 = io_master_ar_valid & T49;
  assign T49 = ar_route[2'h2:2'h2];
  assign io_slave_2_b_ready = b_arb_io_in_2_ready;
  assign io_slave_2_w_bits_user = io_master_w_bits_user;
  assign io_slave_2_w_bits_strb = io_master_w_bits_strb;
  assign io_slave_2_w_bits_last = io_master_w_bits_last;
  assign io_slave_2_w_bits_data = io_master_w_bits_data;
  assign io_slave_2_w_valid = T50;
  assign T50 = io_master_w_valid & R51;
  assign T84 = reset ? 1'h0 : T52;
  assign T52 = T55 ? 1'h0 : T53;
  assign T53 = T54 ? 1'h1 : R51;
  assign T54 = io_slave_2_aw_ready & io_slave_2_aw_valid;
  assign T55 = T56 & io_slave_2_w_bits_last;
  assign T56 = io_slave_2_w_ready & io_slave_2_w_valid;
  assign io_slave_2_aw_bits_user = io_master_aw_bits_user;
  assign io_slave_2_aw_bits_id = io_master_aw_bits_id;
  assign io_slave_2_aw_bits_region = io_master_aw_bits_region;
  assign io_slave_2_aw_bits_qos = io_master_aw_bits_qos;
  assign io_slave_2_aw_bits_prot = io_master_aw_bits_prot;
  assign io_slave_2_aw_bits_cache = io_master_aw_bits_cache;
  assign io_slave_2_aw_bits_lock = io_master_aw_bits_lock;
  assign io_slave_2_aw_bits_burst = io_master_aw_bits_burst;
  assign io_slave_2_aw_bits_size = io_master_aw_bits_size;
  assign io_slave_2_aw_bits_len = io_master_aw_bits_len;
  assign io_slave_2_aw_bits_addr = io_master_aw_bits_addr;
  assign io_slave_2_aw_valid = T57;
  assign T57 = io_master_aw_valid & T58;
  assign T58 = aw_route[2'h2:2'h2];
  assign io_master_r_bits_user = r_arb_io_out_bits_user;
  assign io_master_r_bits_id = r_arb_io_out_bits_id;
  assign io_master_r_bits_last = r_arb_io_out_bits_last;
  assign io_master_r_bits_data = r_arb_io_out_bits_data;
  assign io_master_r_bits_resp = r_arb_io_out_bits_resp;
  assign io_master_r_valid = r_arb_io_out_valid;
  assign io_master_ar_ready = T59;
  assign T59 = ar_ready | T60;
  assign T60 = r_invalid & err_slave_io_ar_ready;
  assign ar_ready = T63 | T61;
  assign T61 = io_slave_2_ar_ready & T62;
  assign T62 = ar_route[2'h2:2'h2];
  assign T63 = T66 | T64;
  assign T64 = io_slave_1_ar_ready & T65;
  assign T65 = ar_route[1'h1:1'h1];
  assign T66 = io_slave_0_ar_ready & T67;
  assign T67 = ar_route[1'h0:1'h0];
  assign io_master_b_bits_user = b_arb_io_out_bits_user;
  assign io_master_b_bits_id = b_arb_io_out_bits_id;
  assign io_master_b_bits_resp = b_arb_io_out_bits_resp;
  assign io_master_b_valid = b_arb_io_out_valid;
  assign io_master_w_ready = T68;
  assign T68 = w_ready | err_slave_io_w_ready;
  assign w_ready = T70 | T69;
  assign T69 = io_slave_2_w_ready & R51;
  assign T70 = T72 | T71;
  assign T71 = io_slave_1_w_ready & R40;
  assign T72 = io_slave_0_w_ready & R29;
  assign io_master_aw_ready = T73;
  assign T73 = aw_ready | T74;
  assign T74 = w_invalid & err_slave_io_aw_ready;
  assign aw_ready = T77 | T75;
  assign T75 = io_slave_2_aw_ready & T76;
  assign T76 = aw_route[2'h2:2'h2];
  assign T77 = T80 | T78;
  assign T78 = io_slave_1_aw_ready & T79;
  assign T79 = aw_route[1'h1:1'h1];
  assign T80 = io_slave_0_aw_ready & T81;
  assign T81 = aw_route[1'h0:1'h0];
  NastiErrorSlave err_slave(.clk(clk), .reset(reset),
       .io_aw_ready( err_slave_io_aw_ready ),
       .io_aw_valid( T13 ),
       .io_aw_bits_addr( io_master_aw_bits_addr ),
       .io_aw_bits_len( io_master_aw_bits_len ),
       .io_aw_bits_size( io_master_aw_bits_size ),
       .io_aw_bits_burst( io_master_aw_bits_burst ),
       .io_aw_bits_lock( io_master_aw_bits_lock ),
       .io_aw_bits_cache( io_master_aw_bits_cache ),
       .io_aw_bits_prot( io_master_aw_bits_prot ),
       .io_aw_bits_qos( io_master_aw_bits_qos ),
       .io_aw_bits_region( io_master_aw_bits_region ),
       .io_aw_bits_id( io_master_aw_bits_id ),
       .io_aw_bits_user( io_master_aw_bits_user ),
       .io_w_ready( err_slave_io_w_ready ),
       .io_w_valid( io_master_w_valid ),
       .io_w_bits_data( io_master_w_bits_data ),
       .io_w_bits_last( io_master_w_bits_last ),
       .io_w_bits_strb( io_master_w_bits_strb ),
       .io_w_bits_user( io_master_w_bits_user ),
       .io_b_ready( b_arb_io_in_3_ready ),
       .io_b_valid( err_slave_io_b_valid ),
       .io_b_bits_resp( err_slave_io_b_bits_resp ),
       .io_b_bits_id( err_slave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( err_slave_io_ar_ready ),
       .io_ar_valid( T0 ),
       .io_ar_bits_addr( io_master_ar_bits_addr ),
       .io_ar_bits_len( io_master_ar_bits_len ),
       .io_ar_bits_size( io_master_ar_bits_size ),
       .io_ar_bits_burst( io_master_ar_bits_burst ),
       .io_ar_bits_lock( io_master_ar_bits_lock ),
       .io_ar_bits_cache( io_master_ar_bits_cache ),
       .io_ar_bits_prot( io_master_ar_bits_prot ),
       .io_ar_bits_qos( io_master_ar_bits_qos ),
       .io_ar_bits_region( io_master_ar_bits_region ),
       .io_ar_bits_id( io_master_ar_bits_id ),
       .io_ar_bits_user( io_master_ar_bits_user ),
       .io_r_ready( r_arb_io_in_3_ready ),
       .io_r_valid( err_slave_io_r_valid ),
       .io_r_bits_resp( err_slave_io_r_bits_resp ),
       .io_r_bits_data( err_slave_io_r_bits_data ),
       .io_r_bits_last( err_slave_io_r_bits_last ),
       .io_r_bits_id( err_slave_io_r_bits_id )
       //.io_r_bits_user(  )
  );
  RRArbiter_4 b_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( b_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_b_valid ),
       .io_in_3_bits_resp( err_slave_io_b_bits_resp ),
       .io_in_3_bits_id( err_slave_io_b_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( b_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_b_valid ),
       .io_in_2_bits_resp( io_slave_2_b_bits_resp ),
       .io_in_2_bits_id( io_slave_2_b_bits_id ),
       .io_in_2_bits_user( io_slave_2_b_bits_user ),
       .io_in_1_ready( b_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_b_valid ),
       .io_in_1_bits_resp( io_slave_1_b_bits_resp ),
       .io_in_1_bits_id( io_slave_1_b_bits_id ),
       .io_in_1_bits_user( io_slave_1_b_bits_user ),
       .io_in_0_ready( b_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_b_valid ),
       .io_in_0_bits_resp( io_slave_0_b_bits_resp ),
       .io_in_0_bits_id( io_slave_0_b_bits_id ),
       .io_in_0_bits_user( io_slave_0_b_bits_user ),
       .io_out_ready( io_master_b_ready ),
       .io_out_valid( b_arb_io_out_valid ),
       .io_out_bits_resp( b_arb_io_out_bits_resp ),
       .io_out_bits_id( b_arb_io_out_bits_id ),
       .io_out_bits_user( b_arb_io_out_bits_user )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign b_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif
  JunctionsPeekingArbiter r_arb(.clk(clk), .reset(reset),
       .io_in_3_ready( r_arb_io_in_3_ready ),
       .io_in_3_valid( err_slave_io_r_valid ),
       .io_in_3_bits_resp( err_slave_io_r_bits_resp ),
       .io_in_3_bits_data( err_slave_io_r_bits_data ),
       .io_in_3_bits_last( err_slave_io_r_bits_last ),
       .io_in_3_bits_id( err_slave_io_r_bits_id ),
       //.io_in_3_bits_user(  )
       .io_in_2_ready( r_arb_io_in_2_ready ),
       .io_in_2_valid( io_slave_2_r_valid ),
       .io_in_2_bits_resp( io_slave_2_r_bits_resp ),
       .io_in_2_bits_data( io_slave_2_r_bits_data ),
       .io_in_2_bits_last( io_slave_2_r_bits_last ),
       .io_in_2_bits_id( io_slave_2_r_bits_id ),
       .io_in_2_bits_user( io_slave_2_r_bits_user ),
       .io_in_1_ready( r_arb_io_in_1_ready ),
       .io_in_1_valid( io_slave_1_r_valid ),
       .io_in_1_bits_resp( io_slave_1_r_bits_resp ),
       .io_in_1_bits_data( io_slave_1_r_bits_data ),
       .io_in_1_bits_last( io_slave_1_r_bits_last ),
       .io_in_1_bits_id( io_slave_1_r_bits_id ),
       .io_in_1_bits_user( io_slave_1_r_bits_user ),
       .io_in_0_ready( r_arb_io_in_0_ready ),
       .io_in_0_valid( io_slave_0_r_valid ),
       .io_in_0_bits_resp( io_slave_0_r_bits_resp ),
       .io_in_0_bits_data( io_slave_0_r_bits_data ),
       .io_in_0_bits_last( io_slave_0_r_bits_last ),
       .io_in_0_bits_id( io_slave_0_r_bits_id ),
       .io_in_0_bits_user( io_slave_0_r_bits_user ),
       .io_out_ready( io_master_r_ready ),
       .io_out_valid( r_arb_io_out_valid ),
       .io_out_bits_resp( r_arb_io_out_bits_resp ),
       .io_out_bits_data( r_arb_io_out_bits_data ),
       .io_out_bits_last( r_arb_io_out_bits_last ),
       .io_out_bits_id( r_arb_io_out_bits_id ),
       .io_out_bits_user( r_arb_io_out_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign r_arb.io_in_3_bits_user = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(reset) begin
      R29 <= 1'h0;
    end else if(T33) begin
      R29 <= 1'h0;
    end else if(T32) begin
      R29 <= 1'h1;
    end
    if(reset) begin
      R40 <= 1'h0;
    end else if(T44) begin
      R40 <= 1'h0;
    end else if(T43) begin
      R40 <= 1'h1;
    end
    if(reset) begin
      R51 <= 1'h0;
    end else if(T55) begin
      R51 <= 1'h0;
    end else if(T54) begin
      R51 <= 1'h1;
    end
  end
endmodule

module NastiCrossbar_1(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [3:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[3:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [3:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[3:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[3:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [3:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[3:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [3:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[3:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [3:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[3:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [3:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[3:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [3:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[3:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [3:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire NastiRouter_io_master_aw_ready;
  wire NastiRouter_io_master_w_ready;
  wire NastiRouter_io_master_b_valid;
  wire[1:0] NastiRouter_io_master_b_bits_resp;
  wire[3:0] NastiRouter_io_master_b_bits_id;
  wire NastiRouter_io_master_b_bits_user;
  wire NastiRouter_io_master_ar_ready;
  wire NastiRouter_io_master_r_valid;
  wire[1:0] NastiRouter_io_master_r_bits_resp;
  wire[63:0] NastiRouter_io_master_r_bits_data;
  wire NastiRouter_io_master_r_bits_last;
  wire[3:0] NastiRouter_io_master_r_bits_id;
  wire NastiRouter_io_master_r_bits_user;
  wire NastiRouter_io_slave_2_aw_valid;
  wire[31:0] NastiRouter_io_slave_2_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_2_aw_bits_burst;
  wire NastiRouter_io_slave_2_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_2_aw_bits_id;
  wire NastiRouter_io_slave_2_aw_bits_user;
  wire NastiRouter_io_slave_2_w_valid;
  wire[63:0] NastiRouter_io_slave_2_w_bits_data;
  wire NastiRouter_io_slave_2_w_bits_last;
  wire[7:0] NastiRouter_io_slave_2_w_bits_strb;
  wire NastiRouter_io_slave_2_w_bits_user;
  wire NastiRouter_io_slave_2_b_ready;
  wire NastiRouter_io_slave_2_ar_valid;
  wire[31:0] NastiRouter_io_slave_2_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_2_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_2_ar_bits_burst;
  wire NastiRouter_io_slave_2_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_2_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_2_ar_bits_id;
  wire NastiRouter_io_slave_2_ar_bits_user;
  wire NastiRouter_io_slave_2_r_ready;
  wire NastiRouter_io_slave_1_aw_valid;
  wire[31:0] NastiRouter_io_slave_1_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_1_aw_bits_burst;
  wire NastiRouter_io_slave_1_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_1_aw_bits_id;
  wire NastiRouter_io_slave_1_aw_bits_user;
  wire NastiRouter_io_slave_1_w_valid;
  wire[63:0] NastiRouter_io_slave_1_w_bits_data;
  wire NastiRouter_io_slave_1_w_bits_last;
  wire[7:0] NastiRouter_io_slave_1_w_bits_strb;
  wire NastiRouter_io_slave_1_w_bits_user;
  wire NastiRouter_io_slave_1_b_ready;
  wire NastiRouter_io_slave_1_ar_valid;
  wire[31:0] NastiRouter_io_slave_1_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_1_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_1_ar_bits_burst;
  wire NastiRouter_io_slave_1_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_1_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_1_ar_bits_id;
  wire NastiRouter_io_slave_1_ar_bits_user;
  wire NastiRouter_io_slave_1_r_ready;
  wire NastiRouter_io_slave_0_aw_valid;
  wire[31:0] NastiRouter_io_slave_0_aw_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_aw_bits_len;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_size;
  wire[1:0] NastiRouter_io_slave_0_aw_bits_burst;
  wire NastiRouter_io_slave_0_aw_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_aw_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_region;
  wire[3:0] NastiRouter_io_slave_0_aw_bits_id;
  wire NastiRouter_io_slave_0_aw_bits_user;
  wire NastiRouter_io_slave_0_w_valid;
  wire[63:0] NastiRouter_io_slave_0_w_bits_data;
  wire NastiRouter_io_slave_0_w_bits_last;
  wire[7:0] NastiRouter_io_slave_0_w_bits_strb;
  wire NastiRouter_io_slave_0_w_bits_user;
  wire NastiRouter_io_slave_0_b_ready;
  wire NastiRouter_io_slave_0_ar_valid;
  wire[31:0] NastiRouter_io_slave_0_ar_bits_addr;
  wire[7:0] NastiRouter_io_slave_0_ar_bits_len;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_size;
  wire[1:0] NastiRouter_io_slave_0_ar_bits_burst;
  wire NastiRouter_io_slave_0_ar_bits_lock;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_cache;
  wire[2:0] NastiRouter_io_slave_0_ar_bits_prot;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_qos;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_region;
  wire[3:0] NastiRouter_io_slave_0_ar_bits_id;
  wire NastiRouter_io_slave_0_ar_bits_user;
  wire NastiRouter_io_slave_0_r_ready;


  assign io_slaves_0_r_ready = NastiRouter_io_slave_0_r_ready;
  assign io_slaves_0_ar_bits_user = NastiRouter_io_slave_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = NastiRouter_io_slave_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = NastiRouter_io_slave_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = NastiRouter_io_slave_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = NastiRouter_io_slave_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = NastiRouter_io_slave_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = NastiRouter_io_slave_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = NastiRouter_io_slave_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = NastiRouter_io_slave_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = NastiRouter_io_slave_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = NastiRouter_io_slave_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = NastiRouter_io_slave_0_ar_valid;
  assign io_slaves_0_b_ready = NastiRouter_io_slave_0_b_ready;
  assign io_slaves_0_w_bits_user = NastiRouter_io_slave_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = NastiRouter_io_slave_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = NastiRouter_io_slave_0_w_bits_last;
  assign io_slaves_0_w_bits_data = NastiRouter_io_slave_0_w_bits_data;
  assign io_slaves_0_w_valid = NastiRouter_io_slave_0_w_valid;
  assign io_slaves_0_aw_bits_user = NastiRouter_io_slave_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = NastiRouter_io_slave_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = NastiRouter_io_slave_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = NastiRouter_io_slave_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = NastiRouter_io_slave_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = NastiRouter_io_slave_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = NastiRouter_io_slave_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = NastiRouter_io_slave_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = NastiRouter_io_slave_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = NastiRouter_io_slave_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = NastiRouter_io_slave_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = NastiRouter_io_slave_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRouter_io_slave_1_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRouter_io_slave_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRouter_io_slave_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRouter_io_slave_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRouter_io_slave_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRouter_io_slave_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRouter_io_slave_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRouter_io_slave_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRouter_io_slave_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRouter_io_slave_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRouter_io_slave_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRouter_io_slave_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRouter_io_slave_1_ar_valid;
  assign io_slaves_1_b_ready = NastiRouter_io_slave_1_b_ready;
  assign io_slaves_1_w_bits_user = NastiRouter_io_slave_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRouter_io_slave_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRouter_io_slave_1_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRouter_io_slave_1_w_bits_data;
  assign io_slaves_1_w_valid = NastiRouter_io_slave_1_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRouter_io_slave_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRouter_io_slave_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRouter_io_slave_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRouter_io_slave_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRouter_io_slave_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRouter_io_slave_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRouter_io_slave_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRouter_io_slave_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRouter_io_slave_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRouter_io_slave_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRouter_io_slave_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRouter_io_slave_1_aw_valid;
  assign io_slaves_2_r_ready = NastiRouter_io_slave_2_r_ready;
  assign io_slaves_2_ar_bits_user = NastiRouter_io_slave_2_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiRouter_io_slave_2_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiRouter_io_slave_2_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiRouter_io_slave_2_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiRouter_io_slave_2_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiRouter_io_slave_2_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiRouter_io_slave_2_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiRouter_io_slave_2_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiRouter_io_slave_2_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiRouter_io_slave_2_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiRouter_io_slave_2_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiRouter_io_slave_2_ar_valid;
  assign io_slaves_2_b_ready = NastiRouter_io_slave_2_b_ready;
  assign io_slaves_2_w_bits_user = NastiRouter_io_slave_2_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiRouter_io_slave_2_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiRouter_io_slave_2_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiRouter_io_slave_2_w_bits_data;
  assign io_slaves_2_w_valid = NastiRouter_io_slave_2_w_valid;
  assign io_slaves_2_aw_bits_user = NastiRouter_io_slave_2_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiRouter_io_slave_2_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiRouter_io_slave_2_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiRouter_io_slave_2_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiRouter_io_slave_2_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiRouter_io_slave_2_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiRouter_io_slave_2_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiRouter_io_slave_2_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiRouter_io_slave_2_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiRouter_io_slave_2_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiRouter_io_slave_2_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiRouter_io_slave_2_aw_valid;
  assign io_masters_0_r_bits_user = NastiRouter_io_master_r_bits_user;
  assign io_masters_0_r_bits_id = NastiRouter_io_master_r_bits_id;
  assign io_masters_0_r_bits_last = NastiRouter_io_master_r_bits_last;
  assign io_masters_0_r_bits_data = NastiRouter_io_master_r_bits_data;
  assign io_masters_0_r_bits_resp = NastiRouter_io_master_r_bits_resp;
  assign io_masters_0_r_valid = NastiRouter_io_master_r_valid;
  assign io_masters_0_ar_ready = NastiRouter_io_master_ar_ready;
  assign io_masters_0_b_bits_user = NastiRouter_io_master_b_bits_user;
  assign io_masters_0_b_bits_id = NastiRouter_io_master_b_bits_id;
  assign io_masters_0_b_bits_resp = NastiRouter_io_master_b_bits_resp;
  assign io_masters_0_b_valid = NastiRouter_io_master_b_valid;
  assign io_masters_0_w_ready = NastiRouter_io_master_w_ready;
  assign io_masters_0_aw_ready = NastiRouter_io_master_aw_ready;
  NastiRouter_1 NastiRouter(.clk(clk), .reset(reset),
       .io_master_aw_ready( NastiRouter_io_master_aw_ready ),
       .io_master_aw_valid( io_masters_0_aw_valid ),
       .io_master_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_master_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_master_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_master_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_master_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_master_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_master_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_master_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_master_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_master_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_master_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_master_w_ready( NastiRouter_io_master_w_ready ),
       .io_master_w_valid( io_masters_0_w_valid ),
       .io_master_w_bits_data( io_masters_0_w_bits_data ),
       .io_master_w_bits_last( io_masters_0_w_bits_last ),
       .io_master_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_master_w_bits_user( io_masters_0_w_bits_user ),
       .io_master_b_ready( io_masters_0_b_ready ),
       .io_master_b_valid( NastiRouter_io_master_b_valid ),
       .io_master_b_bits_resp( NastiRouter_io_master_b_bits_resp ),
       .io_master_b_bits_id( NastiRouter_io_master_b_bits_id ),
       .io_master_b_bits_user( NastiRouter_io_master_b_bits_user ),
       .io_master_ar_ready( NastiRouter_io_master_ar_ready ),
       .io_master_ar_valid( io_masters_0_ar_valid ),
       .io_master_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_master_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_master_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_master_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_master_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_master_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_master_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_master_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_master_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_master_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_master_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_master_r_ready( io_masters_0_r_ready ),
       .io_master_r_valid( NastiRouter_io_master_r_valid ),
       .io_master_r_bits_resp( NastiRouter_io_master_r_bits_resp ),
       .io_master_r_bits_data( NastiRouter_io_master_r_bits_data ),
       .io_master_r_bits_last( NastiRouter_io_master_r_bits_last ),
       .io_master_r_bits_id( NastiRouter_io_master_r_bits_id ),
       .io_master_r_bits_user( NastiRouter_io_master_r_bits_user ),
       .io_slave_2_aw_ready( io_slaves_2_aw_ready ),
       .io_slave_2_aw_valid( NastiRouter_io_slave_2_aw_valid ),
       .io_slave_2_aw_bits_addr( NastiRouter_io_slave_2_aw_bits_addr ),
       .io_slave_2_aw_bits_len( NastiRouter_io_slave_2_aw_bits_len ),
       .io_slave_2_aw_bits_size( NastiRouter_io_slave_2_aw_bits_size ),
       .io_slave_2_aw_bits_burst( NastiRouter_io_slave_2_aw_bits_burst ),
       .io_slave_2_aw_bits_lock( NastiRouter_io_slave_2_aw_bits_lock ),
       .io_slave_2_aw_bits_cache( NastiRouter_io_slave_2_aw_bits_cache ),
       .io_slave_2_aw_bits_prot( NastiRouter_io_slave_2_aw_bits_prot ),
       .io_slave_2_aw_bits_qos( NastiRouter_io_slave_2_aw_bits_qos ),
       .io_slave_2_aw_bits_region( NastiRouter_io_slave_2_aw_bits_region ),
       .io_slave_2_aw_bits_id( NastiRouter_io_slave_2_aw_bits_id ),
       .io_slave_2_aw_bits_user( NastiRouter_io_slave_2_aw_bits_user ),
       .io_slave_2_w_ready( io_slaves_2_w_ready ),
       .io_slave_2_w_valid( NastiRouter_io_slave_2_w_valid ),
       .io_slave_2_w_bits_data( NastiRouter_io_slave_2_w_bits_data ),
       .io_slave_2_w_bits_last( NastiRouter_io_slave_2_w_bits_last ),
       .io_slave_2_w_bits_strb( NastiRouter_io_slave_2_w_bits_strb ),
       .io_slave_2_w_bits_user( NastiRouter_io_slave_2_w_bits_user ),
       .io_slave_2_b_ready( NastiRouter_io_slave_2_b_ready ),
       .io_slave_2_b_valid( io_slaves_2_b_valid ),
       .io_slave_2_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slave_2_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slave_2_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slave_2_ar_ready( io_slaves_2_ar_ready ),
       .io_slave_2_ar_valid( NastiRouter_io_slave_2_ar_valid ),
       .io_slave_2_ar_bits_addr( NastiRouter_io_slave_2_ar_bits_addr ),
       .io_slave_2_ar_bits_len( NastiRouter_io_slave_2_ar_bits_len ),
       .io_slave_2_ar_bits_size( NastiRouter_io_slave_2_ar_bits_size ),
       .io_slave_2_ar_bits_burst( NastiRouter_io_slave_2_ar_bits_burst ),
       .io_slave_2_ar_bits_lock( NastiRouter_io_slave_2_ar_bits_lock ),
       .io_slave_2_ar_bits_cache( NastiRouter_io_slave_2_ar_bits_cache ),
       .io_slave_2_ar_bits_prot( NastiRouter_io_slave_2_ar_bits_prot ),
       .io_slave_2_ar_bits_qos( NastiRouter_io_slave_2_ar_bits_qos ),
       .io_slave_2_ar_bits_region( NastiRouter_io_slave_2_ar_bits_region ),
       .io_slave_2_ar_bits_id( NastiRouter_io_slave_2_ar_bits_id ),
       .io_slave_2_ar_bits_user( NastiRouter_io_slave_2_ar_bits_user ),
       .io_slave_2_r_ready( NastiRouter_io_slave_2_r_ready ),
       .io_slave_2_r_valid( io_slaves_2_r_valid ),
       .io_slave_2_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slave_2_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slave_2_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slave_2_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slave_2_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slave_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slave_1_aw_valid( NastiRouter_io_slave_1_aw_valid ),
       .io_slave_1_aw_bits_addr( NastiRouter_io_slave_1_aw_bits_addr ),
       .io_slave_1_aw_bits_len( NastiRouter_io_slave_1_aw_bits_len ),
       .io_slave_1_aw_bits_size( NastiRouter_io_slave_1_aw_bits_size ),
       .io_slave_1_aw_bits_burst( NastiRouter_io_slave_1_aw_bits_burst ),
       .io_slave_1_aw_bits_lock( NastiRouter_io_slave_1_aw_bits_lock ),
       .io_slave_1_aw_bits_cache( NastiRouter_io_slave_1_aw_bits_cache ),
       .io_slave_1_aw_bits_prot( NastiRouter_io_slave_1_aw_bits_prot ),
       .io_slave_1_aw_bits_qos( NastiRouter_io_slave_1_aw_bits_qos ),
       .io_slave_1_aw_bits_region( NastiRouter_io_slave_1_aw_bits_region ),
       .io_slave_1_aw_bits_id( NastiRouter_io_slave_1_aw_bits_id ),
       .io_slave_1_aw_bits_user( NastiRouter_io_slave_1_aw_bits_user ),
       .io_slave_1_w_ready( io_slaves_1_w_ready ),
       .io_slave_1_w_valid( NastiRouter_io_slave_1_w_valid ),
       .io_slave_1_w_bits_data( NastiRouter_io_slave_1_w_bits_data ),
       .io_slave_1_w_bits_last( NastiRouter_io_slave_1_w_bits_last ),
       .io_slave_1_w_bits_strb( NastiRouter_io_slave_1_w_bits_strb ),
       .io_slave_1_w_bits_user( NastiRouter_io_slave_1_w_bits_user ),
       .io_slave_1_b_ready( NastiRouter_io_slave_1_b_ready ),
       .io_slave_1_b_valid( io_slaves_1_b_valid ),
       .io_slave_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slave_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slave_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slave_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slave_1_ar_valid( NastiRouter_io_slave_1_ar_valid ),
       .io_slave_1_ar_bits_addr( NastiRouter_io_slave_1_ar_bits_addr ),
       .io_slave_1_ar_bits_len( NastiRouter_io_slave_1_ar_bits_len ),
       .io_slave_1_ar_bits_size( NastiRouter_io_slave_1_ar_bits_size ),
       .io_slave_1_ar_bits_burst( NastiRouter_io_slave_1_ar_bits_burst ),
       .io_slave_1_ar_bits_lock( NastiRouter_io_slave_1_ar_bits_lock ),
       .io_slave_1_ar_bits_cache( NastiRouter_io_slave_1_ar_bits_cache ),
       .io_slave_1_ar_bits_prot( NastiRouter_io_slave_1_ar_bits_prot ),
       .io_slave_1_ar_bits_qos( NastiRouter_io_slave_1_ar_bits_qos ),
       .io_slave_1_ar_bits_region( NastiRouter_io_slave_1_ar_bits_region ),
       .io_slave_1_ar_bits_id( NastiRouter_io_slave_1_ar_bits_id ),
       .io_slave_1_ar_bits_user( NastiRouter_io_slave_1_ar_bits_user ),
       .io_slave_1_r_ready( NastiRouter_io_slave_1_r_ready ),
       .io_slave_1_r_valid( io_slaves_1_r_valid ),
       .io_slave_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slave_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slave_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slave_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slave_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slave_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slave_0_aw_valid( NastiRouter_io_slave_0_aw_valid ),
       .io_slave_0_aw_bits_addr( NastiRouter_io_slave_0_aw_bits_addr ),
       .io_slave_0_aw_bits_len( NastiRouter_io_slave_0_aw_bits_len ),
       .io_slave_0_aw_bits_size( NastiRouter_io_slave_0_aw_bits_size ),
       .io_slave_0_aw_bits_burst( NastiRouter_io_slave_0_aw_bits_burst ),
       .io_slave_0_aw_bits_lock( NastiRouter_io_slave_0_aw_bits_lock ),
       .io_slave_0_aw_bits_cache( NastiRouter_io_slave_0_aw_bits_cache ),
       .io_slave_0_aw_bits_prot( NastiRouter_io_slave_0_aw_bits_prot ),
       .io_slave_0_aw_bits_qos( NastiRouter_io_slave_0_aw_bits_qos ),
       .io_slave_0_aw_bits_region( NastiRouter_io_slave_0_aw_bits_region ),
       .io_slave_0_aw_bits_id( NastiRouter_io_slave_0_aw_bits_id ),
       .io_slave_0_aw_bits_user( NastiRouter_io_slave_0_aw_bits_user ),
       .io_slave_0_w_ready( io_slaves_0_w_ready ),
       .io_slave_0_w_valid( NastiRouter_io_slave_0_w_valid ),
       .io_slave_0_w_bits_data( NastiRouter_io_slave_0_w_bits_data ),
       .io_slave_0_w_bits_last( NastiRouter_io_slave_0_w_bits_last ),
       .io_slave_0_w_bits_strb( NastiRouter_io_slave_0_w_bits_strb ),
       .io_slave_0_w_bits_user( NastiRouter_io_slave_0_w_bits_user ),
       .io_slave_0_b_ready( NastiRouter_io_slave_0_b_ready ),
       .io_slave_0_b_valid( io_slaves_0_b_valid ),
       .io_slave_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slave_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slave_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slave_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slave_0_ar_valid( NastiRouter_io_slave_0_ar_valid ),
       .io_slave_0_ar_bits_addr( NastiRouter_io_slave_0_ar_bits_addr ),
       .io_slave_0_ar_bits_len( NastiRouter_io_slave_0_ar_bits_len ),
       .io_slave_0_ar_bits_size( NastiRouter_io_slave_0_ar_bits_size ),
       .io_slave_0_ar_bits_burst( NastiRouter_io_slave_0_ar_bits_burst ),
       .io_slave_0_ar_bits_lock( NastiRouter_io_slave_0_ar_bits_lock ),
       .io_slave_0_ar_bits_cache( NastiRouter_io_slave_0_ar_bits_cache ),
       .io_slave_0_ar_bits_prot( NastiRouter_io_slave_0_ar_bits_prot ),
       .io_slave_0_ar_bits_qos( NastiRouter_io_slave_0_ar_bits_qos ),
       .io_slave_0_ar_bits_region( NastiRouter_io_slave_0_ar_bits_region ),
       .io_slave_0_ar_bits_id( NastiRouter_io_slave_0_ar_bits_id ),
       .io_slave_0_ar_bits_user( NastiRouter_io_slave_0_ar_bits_user ),
       .io_slave_0_r_ready( NastiRouter_io_slave_0_r_ready ),
       .io_slave_0_r_valid( io_slaves_0_r_valid ),
       .io_slave_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slave_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slave_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slave_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slave_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect(input clk, input reset,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [3:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[3:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [3:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[3:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[3:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [3:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[3:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [3:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[3:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [3:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[3:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [3:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[3:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [3:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[3:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [3:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[3:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[3:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_2_aw_valid;
  wire[31:0] xbar_io_slaves_2_aw_bits_addr;
  wire[7:0] xbar_io_slaves_2_aw_bits_len;
  wire[2:0] xbar_io_slaves_2_aw_bits_size;
  wire[1:0] xbar_io_slaves_2_aw_bits_burst;
  wire xbar_io_slaves_2_aw_bits_lock;
  wire[3:0] xbar_io_slaves_2_aw_bits_cache;
  wire[2:0] xbar_io_slaves_2_aw_bits_prot;
  wire[3:0] xbar_io_slaves_2_aw_bits_qos;
  wire[3:0] xbar_io_slaves_2_aw_bits_region;
  wire[3:0] xbar_io_slaves_2_aw_bits_id;
  wire xbar_io_slaves_2_aw_bits_user;
  wire xbar_io_slaves_2_w_valid;
  wire[63:0] xbar_io_slaves_2_w_bits_data;
  wire xbar_io_slaves_2_w_bits_last;
  wire[7:0] xbar_io_slaves_2_w_bits_strb;
  wire xbar_io_slaves_2_w_bits_user;
  wire xbar_io_slaves_2_b_ready;
  wire xbar_io_slaves_2_ar_valid;
  wire[31:0] xbar_io_slaves_2_ar_bits_addr;
  wire[7:0] xbar_io_slaves_2_ar_bits_len;
  wire[2:0] xbar_io_slaves_2_ar_bits_size;
  wire[1:0] xbar_io_slaves_2_ar_bits_burst;
  wire xbar_io_slaves_2_ar_bits_lock;
  wire[3:0] xbar_io_slaves_2_ar_bits_cache;
  wire[2:0] xbar_io_slaves_2_ar_bits_prot;
  wire[3:0] xbar_io_slaves_2_ar_bits_qos;
  wire[3:0] xbar_io_slaves_2_ar_bits_region;
  wire[3:0] xbar_io_slaves_2_ar_bits_id;
  wire xbar_io_slaves_2_ar_bits_user;
  wire xbar_io_slaves_2_r_ready;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[3:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[3:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[3:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[3:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = xbar_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = xbar_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = xbar_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = xbar_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = xbar_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = xbar_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = xbar_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = xbar_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = xbar_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = xbar_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = xbar_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = xbar_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = xbar_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = xbar_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = xbar_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = xbar_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = xbar_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = xbar_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = xbar_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = xbar_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = xbar_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = xbar_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = xbar_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = xbar_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = xbar_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = xbar_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = xbar_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = xbar_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = xbar_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = xbar_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = xbar_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = xbar_io_slaves_1_r_ready;
  assign io_slaves_1_ar_bits_user = xbar_io_slaves_1_ar_bits_user;
  assign io_slaves_1_ar_bits_id = xbar_io_slaves_1_ar_bits_id;
  assign io_slaves_1_ar_bits_region = xbar_io_slaves_1_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = xbar_io_slaves_1_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = xbar_io_slaves_1_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = xbar_io_slaves_1_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = xbar_io_slaves_1_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = xbar_io_slaves_1_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = xbar_io_slaves_1_ar_bits_size;
  assign io_slaves_1_ar_bits_len = xbar_io_slaves_1_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = xbar_io_slaves_1_ar_bits_addr;
  assign io_slaves_1_ar_valid = xbar_io_slaves_1_ar_valid;
  assign io_slaves_1_b_ready = xbar_io_slaves_1_b_ready;
  assign io_slaves_1_w_bits_user = xbar_io_slaves_1_w_bits_user;
  assign io_slaves_1_w_bits_strb = xbar_io_slaves_1_w_bits_strb;
  assign io_slaves_1_w_bits_last = xbar_io_slaves_1_w_bits_last;
  assign io_slaves_1_w_bits_data = xbar_io_slaves_1_w_bits_data;
  assign io_slaves_1_w_valid = xbar_io_slaves_1_w_valid;
  assign io_slaves_1_aw_bits_user = xbar_io_slaves_1_aw_bits_user;
  assign io_slaves_1_aw_bits_id = xbar_io_slaves_1_aw_bits_id;
  assign io_slaves_1_aw_bits_region = xbar_io_slaves_1_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = xbar_io_slaves_1_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = xbar_io_slaves_1_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = xbar_io_slaves_1_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = xbar_io_slaves_1_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = xbar_io_slaves_1_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = xbar_io_slaves_1_aw_bits_size;
  assign io_slaves_1_aw_bits_len = xbar_io_slaves_1_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = xbar_io_slaves_1_aw_bits_addr;
  assign io_slaves_1_aw_valid = xbar_io_slaves_1_aw_valid;
  assign io_slaves_2_r_ready = xbar_io_slaves_2_r_ready;
  assign io_slaves_2_ar_bits_user = xbar_io_slaves_2_ar_bits_user;
  assign io_slaves_2_ar_bits_id = xbar_io_slaves_2_ar_bits_id;
  assign io_slaves_2_ar_bits_region = xbar_io_slaves_2_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = xbar_io_slaves_2_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = xbar_io_slaves_2_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = xbar_io_slaves_2_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = xbar_io_slaves_2_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = xbar_io_slaves_2_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = xbar_io_slaves_2_ar_bits_size;
  assign io_slaves_2_ar_bits_len = xbar_io_slaves_2_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = xbar_io_slaves_2_ar_bits_addr;
  assign io_slaves_2_ar_valid = xbar_io_slaves_2_ar_valid;
  assign io_slaves_2_b_ready = xbar_io_slaves_2_b_ready;
  assign io_slaves_2_w_bits_user = xbar_io_slaves_2_w_bits_user;
  assign io_slaves_2_w_bits_strb = xbar_io_slaves_2_w_bits_strb;
  assign io_slaves_2_w_bits_last = xbar_io_slaves_2_w_bits_last;
  assign io_slaves_2_w_bits_data = xbar_io_slaves_2_w_bits_data;
  assign io_slaves_2_w_valid = xbar_io_slaves_2_w_valid;
  assign io_slaves_2_aw_bits_user = xbar_io_slaves_2_aw_bits_user;
  assign io_slaves_2_aw_bits_id = xbar_io_slaves_2_aw_bits_id;
  assign io_slaves_2_aw_bits_region = xbar_io_slaves_2_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = xbar_io_slaves_2_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = xbar_io_slaves_2_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = xbar_io_slaves_2_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = xbar_io_slaves_2_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = xbar_io_slaves_2_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = xbar_io_slaves_2_aw_bits_size;
  assign io_slaves_2_aw_bits_len = xbar_io_slaves_2_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = xbar_io_slaves_2_aw_bits_addr;
  assign io_slaves_2_aw_valid = xbar_io_slaves_2_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  NastiCrossbar_1 xbar(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_2_aw_ready ),
       .io_slaves_2_aw_valid( xbar_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( xbar_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( xbar_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( xbar_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( xbar_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( xbar_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( xbar_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( xbar_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( xbar_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( xbar_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( xbar_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( xbar_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_2_w_ready ),
       .io_slaves_2_w_valid( xbar_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( xbar_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( xbar_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( xbar_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( xbar_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( xbar_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_2_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_2_ar_ready ),
       .io_slaves_2_ar_valid( xbar_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( xbar_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( xbar_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( xbar_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( xbar_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( xbar_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( xbar_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( xbar_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( xbar_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( xbar_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( xbar_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( xbar_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( xbar_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_2_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_1_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_1_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_1_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_1_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
endmodule

module NastiRecursiveInterconnect_1(input clk, input reset,
    output io_masters_1_aw_ready,
    input  io_masters_1_aw_valid,
    input [31:0] io_masters_1_aw_bits_addr,
    input [7:0] io_masters_1_aw_bits_len,
    input [2:0] io_masters_1_aw_bits_size,
    input [1:0] io_masters_1_aw_bits_burst,
    input  io_masters_1_aw_bits_lock,
    input [3:0] io_masters_1_aw_bits_cache,
    input [2:0] io_masters_1_aw_bits_prot,
    input [3:0] io_masters_1_aw_bits_qos,
    input [3:0] io_masters_1_aw_bits_region,
    input [3:0] io_masters_1_aw_bits_id,
    input  io_masters_1_aw_bits_user,
    output io_masters_1_w_ready,
    input  io_masters_1_w_valid,
    input [63:0] io_masters_1_w_bits_data,
    input  io_masters_1_w_bits_last,
    input [7:0] io_masters_1_w_bits_strb,
    input  io_masters_1_w_bits_user,
    input  io_masters_1_b_ready,
    output io_masters_1_b_valid,
    output[1:0] io_masters_1_b_bits_resp,
    output[3:0] io_masters_1_b_bits_id,
    output io_masters_1_b_bits_user,
    output io_masters_1_ar_ready,
    input  io_masters_1_ar_valid,
    input [31:0] io_masters_1_ar_bits_addr,
    input [7:0] io_masters_1_ar_bits_len,
    input [2:0] io_masters_1_ar_bits_size,
    input [1:0] io_masters_1_ar_bits_burst,
    input  io_masters_1_ar_bits_lock,
    input [3:0] io_masters_1_ar_bits_cache,
    input [2:0] io_masters_1_ar_bits_prot,
    input [3:0] io_masters_1_ar_bits_qos,
    input [3:0] io_masters_1_ar_bits_region,
    input [3:0] io_masters_1_ar_bits_id,
    input  io_masters_1_ar_bits_user,
    input  io_masters_1_r_ready,
    output io_masters_1_r_valid,
    output[1:0] io_masters_1_r_bits_resp,
    output[63:0] io_masters_1_r_bits_data,
    output io_masters_1_r_bits_last,
    output[3:0] io_masters_1_r_bits_id,
    output io_masters_1_r_bits_user,
    output io_masters_0_aw_ready,
    input  io_masters_0_aw_valid,
    input [31:0] io_masters_0_aw_bits_addr,
    input [7:0] io_masters_0_aw_bits_len,
    input [2:0] io_masters_0_aw_bits_size,
    input [1:0] io_masters_0_aw_bits_burst,
    input  io_masters_0_aw_bits_lock,
    input [3:0] io_masters_0_aw_bits_cache,
    input [2:0] io_masters_0_aw_bits_prot,
    input [3:0] io_masters_0_aw_bits_qos,
    input [3:0] io_masters_0_aw_bits_region,
    input [3:0] io_masters_0_aw_bits_id,
    input  io_masters_0_aw_bits_user,
    output io_masters_0_w_ready,
    input  io_masters_0_w_valid,
    input [63:0] io_masters_0_w_bits_data,
    input  io_masters_0_w_bits_last,
    input [7:0] io_masters_0_w_bits_strb,
    input  io_masters_0_w_bits_user,
    input  io_masters_0_b_ready,
    output io_masters_0_b_valid,
    output[1:0] io_masters_0_b_bits_resp,
    output[3:0] io_masters_0_b_bits_id,
    output io_masters_0_b_bits_user,
    output io_masters_0_ar_ready,
    input  io_masters_0_ar_valid,
    input [31:0] io_masters_0_ar_bits_addr,
    input [7:0] io_masters_0_ar_bits_len,
    input [2:0] io_masters_0_ar_bits_size,
    input [1:0] io_masters_0_ar_bits_burst,
    input  io_masters_0_ar_bits_lock,
    input [3:0] io_masters_0_ar_bits_cache,
    input [2:0] io_masters_0_ar_bits_prot,
    input [3:0] io_masters_0_ar_bits_qos,
    input [3:0] io_masters_0_ar_bits_region,
    input [3:0] io_masters_0_ar_bits_id,
    input  io_masters_0_ar_bits_user,
    input  io_masters_0_r_ready,
    output io_masters_0_r_valid,
    output[1:0] io_masters_0_r_bits_resp,
    output[63:0] io_masters_0_r_bits_data,
    output io_masters_0_r_bits_last,
    output[3:0] io_masters_0_r_bits_id,
    output io_masters_0_r_bits_user,
    input  io_slaves_4_aw_ready,
    output io_slaves_4_aw_valid,
    output[31:0] io_slaves_4_aw_bits_addr,
    output[7:0] io_slaves_4_aw_bits_len,
    output[2:0] io_slaves_4_aw_bits_size,
    output[1:0] io_slaves_4_aw_bits_burst,
    output io_slaves_4_aw_bits_lock,
    output[3:0] io_slaves_4_aw_bits_cache,
    output[2:0] io_slaves_4_aw_bits_prot,
    output[3:0] io_slaves_4_aw_bits_qos,
    output[3:0] io_slaves_4_aw_bits_region,
    output[3:0] io_slaves_4_aw_bits_id,
    output io_slaves_4_aw_bits_user,
    input  io_slaves_4_w_ready,
    output io_slaves_4_w_valid,
    output[63:0] io_slaves_4_w_bits_data,
    output io_slaves_4_w_bits_last,
    output[7:0] io_slaves_4_w_bits_strb,
    output io_slaves_4_w_bits_user,
    output io_slaves_4_b_ready,
    input  io_slaves_4_b_valid,
    input [1:0] io_slaves_4_b_bits_resp,
    input [3:0] io_slaves_4_b_bits_id,
    input  io_slaves_4_b_bits_user,
    input  io_slaves_4_ar_ready,
    output io_slaves_4_ar_valid,
    output[31:0] io_slaves_4_ar_bits_addr,
    output[7:0] io_slaves_4_ar_bits_len,
    output[2:0] io_slaves_4_ar_bits_size,
    output[1:0] io_slaves_4_ar_bits_burst,
    output io_slaves_4_ar_bits_lock,
    output[3:0] io_slaves_4_ar_bits_cache,
    output[2:0] io_slaves_4_ar_bits_prot,
    output[3:0] io_slaves_4_ar_bits_qos,
    output[3:0] io_slaves_4_ar_bits_region,
    output[3:0] io_slaves_4_ar_bits_id,
    output io_slaves_4_ar_bits_user,
    output io_slaves_4_r_ready,
    input  io_slaves_4_r_valid,
    input [1:0] io_slaves_4_r_bits_resp,
    input [63:0] io_slaves_4_r_bits_data,
    input  io_slaves_4_r_bits_last,
    input [3:0] io_slaves_4_r_bits_id,
    input  io_slaves_4_r_bits_user,
    input  io_slaves_3_aw_ready,
    output io_slaves_3_aw_valid,
    output[31:0] io_slaves_3_aw_bits_addr,
    output[7:0] io_slaves_3_aw_bits_len,
    output[2:0] io_slaves_3_aw_bits_size,
    output[1:0] io_slaves_3_aw_bits_burst,
    output io_slaves_3_aw_bits_lock,
    output[3:0] io_slaves_3_aw_bits_cache,
    output[2:0] io_slaves_3_aw_bits_prot,
    output[3:0] io_slaves_3_aw_bits_qos,
    output[3:0] io_slaves_3_aw_bits_region,
    output[3:0] io_slaves_3_aw_bits_id,
    output io_slaves_3_aw_bits_user,
    input  io_slaves_3_w_ready,
    output io_slaves_3_w_valid,
    output[63:0] io_slaves_3_w_bits_data,
    output io_slaves_3_w_bits_last,
    output[7:0] io_slaves_3_w_bits_strb,
    output io_slaves_3_w_bits_user,
    output io_slaves_3_b_ready,
    input  io_slaves_3_b_valid,
    input [1:0] io_slaves_3_b_bits_resp,
    input [3:0] io_slaves_3_b_bits_id,
    input  io_slaves_3_b_bits_user,
    input  io_slaves_3_ar_ready,
    output io_slaves_3_ar_valid,
    output[31:0] io_slaves_3_ar_bits_addr,
    output[7:0] io_slaves_3_ar_bits_len,
    output[2:0] io_slaves_3_ar_bits_size,
    output[1:0] io_slaves_3_ar_bits_burst,
    output io_slaves_3_ar_bits_lock,
    output[3:0] io_slaves_3_ar_bits_cache,
    output[2:0] io_slaves_3_ar_bits_prot,
    output[3:0] io_slaves_3_ar_bits_qos,
    output[3:0] io_slaves_3_ar_bits_region,
    output[3:0] io_slaves_3_ar_bits_id,
    output io_slaves_3_ar_bits_user,
    output io_slaves_3_r_ready,
    input  io_slaves_3_r_valid,
    input [1:0] io_slaves_3_r_bits_resp,
    input [63:0] io_slaves_3_r_bits_data,
    input  io_slaves_3_r_bits_last,
    input [3:0] io_slaves_3_r_bits_id,
    input  io_slaves_3_r_bits_user,
    input  io_slaves_2_aw_ready,
    output io_slaves_2_aw_valid,
    output[31:0] io_slaves_2_aw_bits_addr,
    output[7:0] io_slaves_2_aw_bits_len,
    output[2:0] io_slaves_2_aw_bits_size,
    output[1:0] io_slaves_2_aw_bits_burst,
    output io_slaves_2_aw_bits_lock,
    output[3:0] io_slaves_2_aw_bits_cache,
    output[2:0] io_slaves_2_aw_bits_prot,
    output[3:0] io_slaves_2_aw_bits_qos,
    output[3:0] io_slaves_2_aw_bits_region,
    output[3:0] io_slaves_2_aw_bits_id,
    output io_slaves_2_aw_bits_user,
    input  io_slaves_2_w_ready,
    output io_slaves_2_w_valid,
    output[63:0] io_slaves_2_w_bits_data,
    output io_slaves_2_w_bits_last,
    output[7:0] io_slaves_2_w_bits_strb,
    output io_slaves_2_w_bits_user,
    output io_slaves_2_b_ready,
    input  io_slaves_2_b_valid,
    input [1:0] io_slaves_2_b_bits_resp,
    input [3:0] io_slaves_2_b_bits_id,
    input  io_slaves_2_b_bits_user,
    input  io_slaves_2_ar_ready,
    output io_slaves_2_ar_valid,
    output[31:0] io_slaves_2_ar_bits_addr,
    output[7:0] io_slaves_2_ar_bits_len,
    output[2:0] io_slaves_2_ar_bits_size,
    output[1:0] io_slaves_2_ar_bits_burst,
    output io_slaves_2_ar_bits_lock,
    output[3:0] io_slaves_2_ar_bits_cache,
    output[2:0] io_slaves_2_ar_bits_prot,
    output[3:0] io_slaves_2_ar_bits_qos,
    output[3:0] io_slaves_2_ar_bits_region,
    output[3:0] io_slaves_2_ar_bits_id,
    output io_slaves_2_ar_bits_user,
    output io_slaves_2_r_ready,
    input  io_slaves_2_r_valid,
    input [1:0] io_slaves_2_r_bits_resp,
    input [63:0] io_slaves_2_r_bits_data,
    input  io_slaves_2_r_bits_last,
    input [3:0] io_slaves_2_r_bits_id,
    input  io_slaves_2_r_bits_user,
    input  io_slaves_1_aw_ready,
    output io_slaves_1_aw_valid,
    output[31:0] io_slaves_1_aw_bits_addr,
    output[7:0] io_slaves_1_aw_bits_len,
    output[2:0] io_slaves_1_aw_bits_size,
    output[1:0] io_slaves_1_aw_bits_burst,
    output io_slaves_1_aw_bits_lock,
    output[3:0] io_slaves_1_aw_bits_cache,
    output[2:0] io_slaves_1_aw_bits_prot,
    output[3:0] io_slaves_1_aw_bits_qos,
    output[3:0] io_slaves_1_aw_bits_region,
    output[3:0] io_slaves_1_aw_bits_id,
    output io_slaves_1_aw_bits_user,
    input  io_slaves_1_w_ready,
    output io_slaves_1_w_valid,
    output[63:0] io_slaves_1_w_bits_data,
    output io_slaves_1_w_bits_last,
    output[7:0] io_slaves_1_w_bits_strb,
    output io_slaves_1_w_bits_user,
    output io_slaves_1_b_ready,
    input  io_slaves_1_b_valid,
    input [1:0] io_slaves_1_b_bits_resp,
    input [3:0] io_slaves_1_b_bits_id,
    input  io_slaves_1_b_bits_user,
    input  io_slaves_1_ar_ready,
    output io_slaves_1_ar_valid,
    output[31:0] io_slaves_1_ar_bits_addr,
    output[7:0] io_slaves_1_ar_bits_len,
    output[2:0] io_slaves_1_ar_bits_size,
    output[1:0] io_slaves_1_ar_bits_burst,
    output io_slaves_1_ar_bits_lock,
    output[3:0] io_slaves_1_ar_bits_cache,
    output[2:0] io_slaves_1_ar_bits_prot,
    output[3:0] io_slaves_1_ar_bits_qos,
    output[3:0] io_slaves_1_ar_bits_region,
    output[3:0] io_slaves_1_ar_bits_id,
    output io_slaves_1_ar_bits_user,
    output io_slaves_1_r_ready,
    input  io_slaves_1_r_valid,
    input [1:0] io_slaves_1_r_bits_resp,
    input [63:0] io_slaves_1_r_bits_data,
    input  io_slaves_1_r_bits_last,
    input [3:0] io_slaves_1_r_bits_id,
    input  io_slaves_1_r_bits_user,
    input  io_slaves_0_aw_ready,
    output io_slaves_0_aw_valid,
    output[31:0] io_slaves_0_aw_bits_addr,
    output[7:0] io_slaves_0_aw_bits_len,
    output[2:0] io_slaves_0_aw_bits_size,
    output[1:0] io_slaves_0_aw_bits_burst,
    output io_slaves_0_aw_bits_lock,
    output[3:0] io_slaves_0_aw_bits_cache,
    output[2:0] io_slaves_0_aw_bits_prot,
    output[3:0] io_slaves_0_aw_bits_qos,
    output[3:0] io_slaves_0_aw_bits_region,
    output[3:0] io_slaves_0_aw_bits_id,
    output io_slaves_0_aw_bits_user,
    input  io_slaves_0_w_ready,
    output io_slaves_0_w_valid,
    output[63:0] io_slaves_0_w_bits_data,
    output io_slaves_0_w_bits_last,
    output[7:0] io_slaves_0_w_bits_strb,
    output io_slaves_0_w_bits_user,
    output io_slaves_0_b_ready,
    input  io_slaves_0_b_valid,
    input [1:0] io_slaves_0_b_bits_resp,
    input [3:0] io_slaves_0_b_bits_id,
    input  io_slaves_0_b_bits_user,
    input  io_slaves_0_ar_ready,
    output io_slaves_0_ar_valid,
    output[31:0] io_slaves_0_ar_bits_addr,
    output[7:0] io_slaves_0_ar_bits_len,
    output[2:0] io_slaves_0_ar_bits_size,
    output[1:0] io_slaves_0_ar_bits_burst,
    output io_slaves_0_ar_bits_lock,
    output[3:0] io_slaves_0_ar_bits_cache,
    output[2:0] io_slaves_0_ar_bits_prot,
    output[3:0] io_slaves_0_ar_bits_qos,
    output[3:0] io_slaves_0_ar_bits_region,
    output[3:0] io_slaves_0_ar_bits_id,
    output io_slaves_0_ar_bits_user,
    output io_slaves_0_r_ready,
    input  io_slaves_0_r_valid,
    input [1:0] io_slaves_0_r_bits_resp,
    input [63:0] io_slaves_0_r_bits_data,
    input  io_slaves_0_r_bits_last,
    input [3:0] io_slaves_0_r_bits_id,
    input  io_slaves_0_r_bits_user
);

  wire xbar_io_masters_1_aw_ready;
  wire xbar_io_masters_1_w_ready;
  wire xbar_io_masters_1_b_valid;
  wire[1:0] xbar_io_masters_1_b_bits_resp;
  wire[3:0] xbar_io_masters_1_b_bits_id;
  wire xbar_io_masters_1_b_bits_user;
  wire xbar_io_masters_1_ar_ready;
  wire xbar_io_masters_1_r_valid;
  wire[1:0] xbar_io_masters_1_r_bits_resp;
  wire[63:0] xbar_io_masters_1_r_bits_data;
  wire xbar_io_masters_1_r_bits_last;
  wire[3:0] xbar_io_masters_1_r_bits_id;
  wire xbar_io_masters_1_r_bits_user;
  wire xbar_io_masters_0_aw_ready;
  wire xbar_io_masters_0_w_ready;
  wire xbar_io_masters_0_b_valid;
  wire[1:0] xbar_io_masters_0_b_bits_resp;
  wire[3:0] xbar_io_masters_0_b_bits_id;
  wire xbar_io_masters_0_b_bits_user;
  wire xbar_io_masters_0_ar_ready;
  wire xbar_io_masters_0_r_valid;
  wire[1:0] xbar_io_masters_0_r_bits_resp;
  wire[63:0] xbar_io_masters_0_r_bits_data;
  wire xbar_io_masters_0_r_bits_last;
  wire[3:0] xbar_io_masters_0_r_bits_id;
  wire xbar_io_masters_0_r_bits_user;
  wire xbar_io_slaves_2_aw_valid;
  wire[31:0] xbar_io_slaves_2_aw_bits_addr;
  wire[7:0] xbar_io_slaves_2_aw_bits_len;
  wire[2:0] xbar_io_slaves_2_aw_bits_size;
  wire[1:0] xbar_io_slaves_2_aw_bits_burst;
  wire xbar_io_slaves_2_aw_bits_lock;
  wire[3:0] xbar_io_slaves_2_aw_bits_cache;
  wire[2:0] xbar_io_slaves_2_aw_bits_prot;
  wire[3:0] xbar_io_slaves_2_aw_bits_qos;
  wire[3:0] xbar_io_slaves_2_aw_bits_region;
  wire[3:0] xbar_io_slaves_2_aw_bits_id;
  wire xbar_io_slaves_2_aw_bits_user;
  wire xbar_io_slaves_2_w_valid;
  wire[63:0] xbar_io_slaves_2_w_bits_data;
  wire xbar_io_slaves_2_w_bits_last;
  wire[7:0] xbar_io_slaves_2_w_bits_strb;
  wire xbar_io_slaves_2_w_bits_user;
  wire xbar_io_slaves_2_b_ready;
  wire xbar_io_slaves_2_ar_valid;
  wire[31:0] xbar_io_slaves_2_ar_bits_addr;
  wire[7:0] xbar_io_slaves_2_ar_bits_len;
  wire[2:0] xbar_io_slaves_2_ar_bits_size;
  wire[1:0] xbar_io_slaves_2_ar_bits_burst;
  wire xbar_io_slaves_2_ar_bits_lock;
  wire[3:0] xbar_io_slaves_2_ar_bits_cache;
  wire[2:0] xbar_io_slaves_2_ar_bits_prot;
  wire[3:0] xbar_io_slaves_2_ar_bits_qos;
  wire[3:0] xbar_io_slaves_2_ar_bits_region;
  wire[3:0] xbar_io_slaves_2_ar_bits_id;
  wire xbar_io_slaves_2_ar_bits_user;
  wire xbar_io_slaves_2_r_ready;
  wire xbar_io_slaves_1_aw_valid;
  wire[31:0] xbar_io_slaves_1_aw_bits_addr;
  wire[7:0] xbar_io_slaves_1_aw_bits_len;
  wire[2:0] xbar_io_slaves_1_aw_bits_size;
  wire[1:0] xbar_io_slaves_1_aw_bits_burst;
  wire xbar_io_slaves_1_aw_bits_lock;
  wire[3:0] xbar_io_slaves_1_aw_bits_cache;
  wire[2:0] xbar_io_slaves_1_aw_bits_prot;
  wire[3:0] xbar_io_slaves_1_aw_bits_qos;
  wire[3:0] xbar_io_slaves_1_aw_bits_region;
  wire[3:0] xbar_io_slaves_1_aw_bits_id;
  wire xbar_io_slaves_1_aw_bits_user;
  wire xbar_io_slaves_1_w_valid;
  wire[63:0] xbar_io_slaves_1_w_bits_data;
  wire xbar_io_slaves_1_w_bits_last;
  wire[7:0] xbar_io_slaves_1_w_bits_strb;
  wire xbar_io_slaves_1_w_bits_user;
  wire xbar_io_slaves_1_b_ready;
  wire xbar_io_slaves_1_ar_valid;
  wire[31:0] xbar_io_slaves_1_ar_bits_addr;
  wire[7:0] xbar_io_slaves_1_ar_bits_len;
  wire[2:0] xbar_io_slaves_1_ar_bits_size;
  wire[1:0] xbar_io_slaves_1_ar_bits_burst;
  wire xbar_io_slaves_1_ar_bits_lock;
  wire[3:0] xbar_io_slaves_1_ar_bits_cache;
  wire[2:0] xbar_io_slaves_1_ar_bits_prot;
  wire[3:0] xbar_io_slaves_1_ar_bits_qos;
  wire[3:0] xbar_io_slaves_1_ar_bits_region;
  wire[3:0] xbar_io_slaves_1_ar_bits_id;
  wire xbar_io_slaves_1_ar_bits_user;
  wire xbar_io_slaves_1_r_ready;
  wire xbar_io_slaves_0_aw_valid;
  wire[31:0] xbar_io_slaves_0_aw_bits_addr;
  wire[7:0] xbar_io_slaves_0_aw_bits_len;
  wire[2:0] xbar_io_slaves_0_aw_bits_size;
  wire[1:0] xbar_io_slaves_0_aw_bits_burst;
  wire xbar_io_slaves_0_aw_bits_lock;
  wire[3:0] xbar_io_slaves_0_aw_bits_cache;
  wire[2:0] xbar_io_slaves_0_aw_bits_prot;
  wire[3:0] xbar_io_slaves_0_aw_bits_qos;
  wire[3:0] xbar_io_slaves_0_aw_bits_region;
  wire[3:0] xbar_io_slaves_0_aw_bits_id;
  wire xbar_io_slaves_0_aw_bits_user;
  wire xbar_io_slaves_0_w_valid;
  wire[63:0] xbar_io_slaves_0_w_bits_data;
  wire xbar_io_slaves_0_w_bits_last;
  wire[7:0] xbar_io_slaves_0_w_bits_strb;
  wire xbar_io_slaves_0_w_bits_user;
  wire xbar_io_slaves_0_b_ready;
  wire xbar_io_slaves_0_ar_valid;
  wire[31:0] xbar_io_slaves_0_ar_bits_addr;
  wire[7:0] xbar_io_slaves_0_ar_bits_len;
  wire[2:0] xbar_io_slaves_0_ar_bits_size;
  wire[1:0] xbar_io_slaves_0_ar_bits_burst;
  wire xbar_io_slaves_0_ar_bits_lock;
  wire[3:0] xbar_io_slaves_0_ar_bits_cache;
  wire[2:0] xbar_io_slaves_0_ar_bits_prot;
  wire[3:0] xbar_io_slaves_0_ar_bits_qos;
  wire[3:0] xbar_io_slaves_0_ar_bits_region;
  wire[3:0] xbar_io_slaves_0_ar_bits_id;
  wire xbar_io_slaves_0_ar_bits_user;
  wire xbar_io_slaves_0_r_ready;
  wire NastiRecursiveInterconnect_io_masters_0_aw_ready;
  wire NastiRecursiveInterconnect_io_masters_0_w_ready;
  wire NastiRecursiveInterconnect_io_masters_0_b_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_b_bits_resp;
  wire[3:0] NastiRecursiveInterconnect_io_masters_0_b_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_b_bits_user;
  wire NastiRecursiveInterconnect_io_masters_0_ar_ready;
  wire NastiRecursiveInterconnect_io_masters_0_r_valid;
  wire[1:0] NastiRecursiveInterconnect_io_masters_0_r_bits_resp;
  wire[63:0] NastiRecursiveInterconnect_io_masters_0_r_bits_data;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_last;
  wire[3:0] NastiRecursiveInterconnect_io_masters_0_r_bits_id;
  wire NastiRecursiveInterconnect_io_masters_0_r_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_2_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_2_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_2_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_2_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_2_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_2_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_2_r_ready;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_1_r_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_w_valid;
  wire[63:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  wire NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_b_ready;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  wire[31:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  wire[7:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  wire[1:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  wire[2:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  wire[3:0] NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  wire NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  wire NastiRecursiveInterconnect_io_slaves_0_r_ready;


  assign io_slaves_0_r_ready = xbar_io_slaves_0_r_ready;
  assign io_slaves_0_ar_bits_user = xbar_io_slaves_0_ar_bits_user;
  assign io_slaves_0_ar_bits_id = xbar_io_slaves_0_ar_bits_id;
  assign io_slaves_0_ar_bits_region = xbar_io_slaves_0_ar_bits_region;
  assign io_slaves_0_ar_bits_qos = xbar_io_slaves_0_ar_bits_qos;
  assign io_slaves_0_ar_bits_prot = xbar_io_slaves_0_ar_bits_prot;
  assign io_slaves_0_ar_bits_cache = xbar_io_slaves_0_ar_bits_cache;
  assign io_slaves_0_ar_bits_lock = xbar_io_slaves_0_ar_bits_lock;
  assign io_slaves_0_ar_bits_burst = xbar_io_slaves_0_ar_bits_burst;
  assign io_slaves_0_ar_bits_size = xbar_io_slaves_0_ar_bits_size;
  assign io_slaves_0_ar_bits_len = xbar_io_slaves_0_ar_bits_len;
  assign io_slaves_0_ar_bits_addr = xbar_io_slaves_0_ar_bits_addr;
  assign io_slaves_0_ar_valid = xbar_io_slaves_0_ar_valid;
  assign io_slaves_0_b_ready = xbar_io_slaves_0_b_ready;
  assign io_slaves_0_w_bits_user = xbar_io_slaves_0_w_bits_user;
  assign io_slaves_0_w_bits_strb = xbar_io_slaves_0_w_bits_strb;
  assign io_slaves_0_w_bits_last = xbar_io_slaves_0_w_bits_last;
  assign io_slaves_0_w_bits_data = xbar_io_slaves_0_w_bits_data;
  assign io_slaves_0_w_valid = xbar_io_slaves_0_w_valid;
  assign io_slaves_0_aw_bits_user = xbar_io_slaves_0_aw_bits_user;
  assign io_slaves_0_aw_bits_id = xbar_io_slaves_0_aw_bits_id;
  assign io_slaves_0_aw_bits_region = xbar_io_slaves_0_aw_bits_region;
  assign io_slaves_0_aw_bits_qos = xbar_io_slaves_0_aw_bits_qos;
  assign io_slaves_0_aw_bits_prot = xbar_io_slaves_0_aw_bits_prot;
  assign io_slaves_0_aw_bits_cache = xbar_io_slaves_0_aw_bits_cache;
  assign io_slaves_0_aw_bits_lock = xbar_io_slaves_0_aw_bits_lock;
  assign io_slaves_0_aw_bits_burst = xbar_io_slaves_0_aw_bits_burst;
  assign io_slaves_0_aw_bits_size = xbar_io_slaves_0_aw_bits_size;
  assign io_slaves_0_aw_bits_len = xbar_io_slaves_0_aw_bits_len;
  assign io_slaves_0_aw_bits_addr = xbar_io_slaves_0_aw_bits_addr;
  assign io_slaves_0_aw_valid = xbar_io_slaves_0_aw_valid;
  assign io_slaves_1_r_ready = NastiRecursiveInterconnect_io_slaves_0_r_ready;
  assign io_slaves_1_ar_bits_user = NastiRecursiveInterconnect_io_slaves_0_ar_bits_user;
  assign io_slaves_1_ar_bits_id = NastiRecursiveInterconnect_io_slaves_0_ar_bits_id;
  assign io_slaves_1_ar_bits_region = NastiRecursiveInterconnect_io_slaves_0_ar_bits_region;
  assign io_slaves_1_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos;
  assign io_slaves_1_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot;
  assign io_slaves_1_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache;
  assign io_slaves_1_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock;
  assign io_slaves_1_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst;
  assign io_slaves_1_ar_bits_size = NastiRecursiveInterconnect_io_slaves_0_ar_bits_size;
  assign io_slaves_1_ar_bits_len = NastiRecursiveInterconnect_io_slaves_0_ar_bits_len;
  assign io_slaves_1_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr;
  assign io_slaves_1_ar_valid = NastiRecursiveInterconnect_io_slaves_0_ar_valid;
  assign io_slaves_1_b_ready = NastiRecursiveInterconnect_io_slaves_0_b_ready;
  assign io_slaves_1_w_bits_user = NastiRecursiveInterconnect_io_slaves_0_w_bits_user;
  assign io_slaves_1_w_bits_strb = NastiRecursiveInterconnect_io_slaves_0_w_bits_strb;
  assign io_slaves_1_w_bits_last = NastiRecursiveInterconnect_io_slaves_0_w_bits_last;
  assign io_slaves_1_w_bits_data = NastiRecursiveInterconnect_io_slaves_0_w_bits_data;
  assign io_slaves_1_w_valid = NastiRecursiveInterconnect_io_slaves_0_w_valid;
  assign io_slaves_1_aw_bits_user = NastiRecursiveInterconnect_io_slaves_0_aw_bits_user;
  assign io_slaves_1_aw_bits_id = NastiRecursiveInterconnect_io_slaves_0_aw_bits_id;
  assign io_slaves_1_aw_bits_region = NastiRecursiveInterconnect_io_slaves_0_aw_bits_region;
  assign io_slaves_1_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos;
  assign io_slaves_1_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot;
  assign io_slaves_1_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache;
  assign io_slaves_1_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock;
  assign io_slaves_1_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst;
  assign io_slaves_1_aw_bits_size = NastiRecursiveInterconnect_io_slaves_0_aw_bits_size;
  assign io_slaves_1_aw_bits_len = NastiRecursiveInterconnect_io_slaves_0_aw_bits_len;
  assign io_slaves_1_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr;
  assign io_slaves_1_aw_valid = NastiRecursiveInterconnect_io_slaves_0_aw_valid;
  assign io_slaves_2_r_ready = NastiRecursiveInterconnect_io_slaves_1_r_ready;
  assign io_slaves_2_ar_bits_user = NastiRecursiveInterconnect_io_slaves_1_ar_bits_user;
  assign io_slaves_2_ar_bits_id = NastiRecursiveInterconnect_io_slaves_1_ar_bits_id;
  assign io_slaves_2_ar_bits_region = NastiRecursiveInterconnect_io_slaves_1_ar_bits_region;
  assign io_slaves_2_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos;
  assign io_slaves_2_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot;
  assign io_slaves_2_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache;
  assign io_slaves_2_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock;
  assign io_slaves_2_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst;
  assign io_slaves_2_ar_bits_size = NastiRecursiveInterconnect_io_slaves_1_ar_bits_size;
  assign io_slaves_2_ar_bits_len = NastiRecursiveInterconnect_io_slaves_1_ar_bits_len;
  assign io_slaves_2_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr;
  assign io_slaves_2_ar_valid = NastiRecursiveInterconnect_io_slaves_1_ar_valid;
  assign io_slaves_2_b_ready = NastiRecursiveInterconnect_io_slaves_1_b_ready;
  assign io_slaves_2_w_bits_user = NastiRecursiveInterconnect_io_slaves_1_w_bits_user;
  assign io_slaves_2_w_bits_strb = NastiRecursiveInterconnect_io_slaves_1_w_bits_strb;
  assign io_slaves_2_w_bits_last = NastiRecursiveInterconnect_io_slaves_1_w_bits_last;
  assign io_slaves_2_w_bits_data = NastiRecursiveInterconnect_io_slaves_1_w_bits_data;
  assign io_slaves_2_w_valid = NastiRecursiveInterconnect_io_slaves_1_w_valid;
  assign io_slaves_2_aw_bits_user = NastiRecursiveInterconnect_io_slaves_1_aw_bits_user;
  assign io_slaves_2_aw_bits_id = NastiRecursiveInterconnect_io_slaves_1_aw_bits_id;
  assign io_slaves_2_aw_bits_region = NastiRecursiveInterconnect_io_slaves_1_aw_bits_region;
  assign io_slaves_2_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos;
  assign io_slaves_2_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot;
  assign io_slaves_2_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache;
  assign io_slaves_2_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock;
  assign io_slaves_2_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst;
  assign io_slaves_2_aw_bits_size = NastiRecursiveInterconnect_io_slaves_1_aw_bits_size;
  assign io_slaves_2_aw_bits_len = NastiRecursiveInterconnect_io_slaves_1_aw_bits_len;
  assign io_slaves_2_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr;
  assign io_slaves_2_aw_valid = NastiRecursiveInterconnect_io_slaves_1_aw_valid;
  assign io_slaves_3_r_ready = NastiRecursiveInterconnect_io_slaves_2_r_ready;
  assign io_slaves_3_ar_bits_user = NastiRecursiveInterconnect_io_slaves_2_ar_bits_user;
  assign io_slaves_3_ar_bits_id = NastiRecursiveInterconnect_io_slaves_2_ar_bits_id;
  assign io_slaves_3_ar_bits_region = NastiRecursiveInterconnect_io_slaves_2_ar_bits_region;
  assign io_slaves_3_ar_bits_qos = NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos;
  assign io_slaves_3_ar_bits_prot = NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot;
  assign io_slaves_3_ar_bits_cache = NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache;
  assign io_slaves_3_ar_bits_lock = NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock;
  assign io_slaves_3_ar_bits_burst = NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst;
  assign io_slaves_3_ar_bits_size = NastiRecursiveInterconnect_io_slaves_2_ar_bits_size;
  assign io_slaves_3_ar_bits_len = NastiRecursiveInterconnect_io_slaves_2_ar_bits_len;
  assign io_slaves_3_ar_bits_addr = NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr;
  assign io_slaves_3_ar_valid = NastiRecursiveInterconnect_io_slaves_2_ar_valid;
  assign io_slaves_3_b_ready = NastiRecursiveInterconnect_io_slaves_2_b_ready;
  assign io_slaves_3_w_bits_user = NastiRecursiveInterconnect_io_slaves_2_w_bits_user;
  assign io_slaves_3_w_bits_strb = NastiRecursiveInterconnect_io_slaves_2_w_bits_strb;
  assign io_slaves_3_w_bits_last = NastiRecursiveInterconnect_io_slaves_2_w_bits_last;
  assign io_slaves_3_w_bits_data = NastiRecursiveInterconnect_io_slaves_2_w_bits_data;
  assign io_slaves_3_w_valid = NastiRecursiveInterconnect_io_slaves_2_w_valid;
  assign io_slaves_3_aw_bits_user = NastiRecursiveInterconnect_io_slaves_2_aw_bits_user;
  assign io_slaves_3_aw_bits_id = NastiRecursiveInterconnect_io_slaves_2_aw_bits_id;
  assign io_slaves_3_aw_bits_region = NastiRecursiveInterconnect_io_slaves_2_aw_bits_region;
  assign io_slaves_3_aw_bits_qos = NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos;
  assign io_slaves_3_aw_bits_prot = NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot;
  assign io_slaves_3_aw_bits_cache = NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache;
  assign io_slaves_3_aw_bits_lock = NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock;
  assign io_slaves_3_aw_bits_burst = NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst;
  assign io_slaves_3_aw_bits_size = NastiRecursiveInterconnect_io_slaves_2_aw_bits_size;
  assign io_slaves_3_aw_bits_len = NastiRecursiveInterconnect_io_slaves_2_aw_bits_len;
  assign io_slaves_3_aw_bits_addr = NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr;
  assign io_slaves_3_aw_valid = NastiRecursiveInterconnect_io_slaves_2_aw_valid;
  assign io_slaves_4_r_ready = xbar_io_slaves_2_r_ready;
  assign io_slaves_4_ar_bits_user = xbar_io_slaves_2_ar_bits_user;
  assign io_slaves_4_ar_bits_id = xbar_io_slaves_2_ar_bits_id;
  assign io_slaves_4_ar_bits_region = xbar_io_slaves_2_ar_bits_region;
  assign io_slaves_4_ar_bits_qos = xbar_io_slaves_2_ar_bits_qos;
  assign io_slaves_4_ar_bits_prot = xbar_io_slaves_2_ar_bits_prot;
  assign io_slaves_4_ar_bits_cache = xbar_io_slaves_2_ar_bits_cache;
  assign io_slaves_4_ar_bits_lock = xbar_io_slaves_2_ar_bits_lock;
  assign io_slaves_4_ar_bits_burst = xbar_io_slaves_2_ar_bits_burst;
  assign io_slaves_4_ar_bits_size = xbar_io_slaves_2_ar_bits_size;
  assign io_slaves_4_ar_bits_len = xbar_io_slaves_2_ar_bits_len;
  assign io_slaves_4_ar_bits_addr = xbar_io_slaves_2_ar_bits_addr;
  assign io_slaves_4_ar_valid = xbar_io_slaves_2_ar_valid;
  assign io_slaves_4_b_ready = xbar_io_slaves_2_b_ready;
  assign io_slaves_4_w_bits_user = xbar_io_slaves_2_w_bits_user;
  assign io_slaves_4_w_bits_strb = xbar_io_slaves_2_w_bits_strb;
  assign io_slaves_4_w_bits_last = xbar_io_slaves_2_w_bits_last;
  assign io_slaves_4_w_bits_data = xbar_io_slaves_2_w_bits_data;
  assign io_slaves_4_w_valid = xbar_io_slaves_2_w_valid;
  assign io_slaves_4_aw_bits_user = xbar_io_slaves_2_aw_bits_user;
  assign io_slaves_4_aw_bits_id = xbar_io_slaves_2_aw_bits_id;
  assign io_slaves_4_aw_bits_region = xbar_io_slaves_2_aw_bits_region;
  assign io_slaves_4_aw_bits_qos = xbar_io_slaves_2_aw_bits_qos;
  assign io_slaves_4_aw_bits_prot = xbar_io_slaves_2_aw_bits_prot;
  assign io_slaves_4_aw_bits_cache = xbar_io_slaves_2_aw_bits_cache;
  assign io_slaves_4_aw_bits_lock = xbar_io_slaves_2_aw_bits_lock;
  assign io_slaves_4_aw_bits_burst = xbar_io_slaves_2_aw_bits_burst;
  assign io_slaves_4_aw_bits_size = xbar_io_slaves_2_aw_bits_size;
  assign io_slaves_4_aw_bits_len = xbar_io_slaves_2_aw_bits_len;
  assign io_slaves_4_aw_bits_addr = xbar_io_slaves_2_aw_bits_addr;
  assign io_slaves_4_aw_valid = xbar_io_slaves_2_aw_valid;
  assign io_masters_0_r_bits_user = xbar_io_masters_0_r_bits_user;
  assign io_masters_0_r_bits_id = xbar_io_masters_0_r_bits_id;
  assign io_masters_0_r_bits_last = xbar_io_masters_0_r_bits_last;
  assign io_masters_0_r_bits_data = xbar_io_masters_0_r_bits_data;
  assign io_masters_0_r_bits_resp = xbar_io_masters_0_r_bits_resp;
  assign io_masters_0_r_valid = xbar_io_masters_0_r_valid;
  assign io_masters_0_ar_ready = xbar_io_masters_0_ar_ready;
  assign io_masters_0_b_bits_user = xbar_io_masters_0_b_bits_user;
  assign io_masters_0_b_bits_id = xbar_io_masters_0_b_bits_id;
  assign io_masters_0_b_bits_resp = xbar_io_masters_0_b_bits_resp;
  assign io_masters_0_b_valid = xbar_io_masters_0_b_valid;
  assign io_masters_0_w_ready = xbar_io_masters_0_w_ready;
  assign io_masters_0_aw_ready = xbar_io_masters_0_aw_ready;
  assign io_masters_1_r_bits_user = xbar_io_masters_1_r_bits_user;
  assign io_masters_1_r_bits_id = xbar_io_masters_1_r_bits_id;
  assign io_masters_1_r_bits_last = xbar_io_masters_1_r_bits_last;
  assign io_masters_1_r_bits_data = xbar_io_masters_1_r_bits_data;
  assign io_masters_1_r_bits_resp = xbar_io_masters_1_r_bits_resp;
  assign io_masters_1_r_valid = xbar_io_masters_1_r_valid;
  assign io_masters_1_ar_ready = xbar_io_masters_1_ar_ready;
  assign io_masters_1_b_bits_user = xbar_io_masters_1_b_bits_user;
  assign io_masters_1_b_bits_id = xbar_io_masters_1_b_bits_id;
  assign io_masters_1_b_bits_resp = xbar_io_masters_1_b_bits_resp;
  assign io_masters_1_b_valid = xbar_io_masters_1_b_valid;
  assign io_masters_1_w_ready = xbar_io_masters_1_w_ready;
  assign io_masters_1_aw_ready = xbar_io_masters_1_aw_ready;
  NastiCrossbar_0 xbar(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( xbar_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( io_masters_1_aw_valid ),
       .io_masters_1_aw_bits_addr( io_masters_1_aw_bits_addr ),
       .io_masters_1_aw_bits_len( io_masters_1_aw_bits_len ),
       .io_masters_1_aw_bits_size( io_masters_1_aw_bits_size ),
       .io_masters_1_aw_bits_burst( io_masters_1_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( io_masters_1_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( io_masters_1_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( io_masters_1_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( io_masters_1_aw_bits_qos ),
       .io_masters_1_aw_bits_region( io_masters_1_aw_bits_region ),
       .io_masters_1_aw_bits_id( io_masters_1_aw_bits_id ),
       .io_masters_1_aw_bits_user( io_masters_1_aw_bits_user ),
       .io_masters_1_w_ready( xbar_io_masters_1_w_ready ),
       .io_masters_1_w_valid( io_masters_1_w_valid ),
       .io_masters_1_w_bits_data( io_masters_1_w_bits_data ),
       .io_masters_1_w_bits_last( io_masters_1_w_bits_last ),
       .io_masters_1_w_bits_strb( io_masters_1_w_bits_strb ),
       .io_masters_1_w_bits_user( io_masters_1_w_bits_user ),
       .io_masters_1_b_ready( io_masters_1_b_ready ),
       .io_masters_1_b_valid( xbar_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( xbar_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( xbar_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( xbar_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( xbar_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( io_masters_1_ar_valid ),
       .io_masters_1_ar_bits_addr( io_masters_1_ar_bits_addr ),
       .io_masters_1_ar_bits_len( io_masters_1_ar_bits_len ),
       .io_masters_1_ar_bits_size( io_masters_1_ar_bits_size ),
       .io_masters_1_ar_bits_burst( io_masters_1_ar_bits_burst ),
       .io_masters_1_ar_bits_lock( io_masters_1_ar_bits_lock ),
       .io_masters_1_ar_bits_cache( io_masters_1_ar_bits_cache ),
       .io_masters_1_ar_bits_prot( io_masters_1_ar_bits_prot ),
       .io_masters_1_ar_bits_qos( io_masters_1_ar_bits_qos ),
       .io_masters_1_ar_bits_region( io_masters_1_ar_bits_region ),
       .io_masters_1_ar_bits_id( io_masters_1_ar_bits_id ),
       .io_masters_1_ar_bits_user( io_masters_1_ar_bits_user ),
       .io_masters_1_r_ready( io_masters_1_r_ready ),
       .io_masters_1_r_valid( xbar_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( xbar_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( xbar_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( xbar_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( xbar_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( xbar_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( xbar_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( io_masters_0_aw_valid ),
       .io_masters_0_aw_bits_addr( io_masters_0_aw_bits_addr ),
       .io_masters_0_aw_bits_len( io_masters_0_aw_bits_len ),
       .io_masters_0_aw_bits_size( io_masters_0_aw_bits_size ),
       .io_masters_0_aw_bits_burst( io_masters_0_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( io_masters_0_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( io_masters_0_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( io_masters_0_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( io_masters_0_aw_bits_qos ),
       .io_masters_0_aw_bits_region( io_masters_0_aw_bits_region ),
       .io_masters_0_aw_bits_id( io_masters_0_aw_bits_id ),
       .io_masters_0_aw_bits_user( io_masters_0_aw_bits_user ),
       .io_masters_0_w_ready( xbar_io_masters_0_w_ready ),
       .io_masters_0_w_valid( io_masters_0_w_valid ),
       .io_masters_0_w_bits_data( io_masters_0_w_bits_data ),
       .io_masters_0_w_bits_last( io_masters_0_w_bits_last ),
       .io_masters_0_w_bits_strb( io_masters_0_w_bits_strb ),
       .io_masters_0_w_bits_user( io_masters_0_w_bits_user ),
       .io_masters_0_b_ready( io_masters_0_b_ready ),
       .io_masters_0_b_valid( xbar_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( xbar_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( xbar_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( xbar_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( xbar_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( io_masters_0_ar_valid ),
       .io_masters_0_ar_bits_addr( io_masters_0_ar_bits_addr ),
       .io_masters_0_ar_bits_len( io_masters_0_ar_bits_len ),
       .io_masters_0_ar_bits_size( io_masters_0_ar_bits_size ),
       .io_masters_0_ar_bits_burst( io_masters_0_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( io_masters_0_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( io_masters_0_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( io_masters_0_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( io_masters_0_ar_bits_qos ),
       .io_masters_0_ar_bits_region( io_masters_0_ar_bits_region ),
       .io_masters_0_ar_bits_id( io_masters_0_ar_bits_id ),
       .io_masters_0_ar_bits_user( io_masters_0_ar_bits_user ),
       .io_masters_0_r_ready( io_masters_0_r_ready ),
       .io_masters_0_r_valid( xbar_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( xbar_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( xbar_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( xbar_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( xbar_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( xbar_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_4_aw_ready ),
       .io_slaves_2_aw_valid( xbar_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( xbar_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( xbar_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( xbar_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( xbar_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( xbar_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( xbar_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( xbar_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( xbar_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( xbar_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( xbar_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( xbar_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_4_w_ready ),
       .io_slaves_2_w_valid( xbar_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( xbar_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( xbar_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( xbar_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( xbar_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( xbar_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_4_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_4_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_4_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_4_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_4_ar_ready ),
       .io_slaves_2_ar_valid( xbar_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( xbar_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( xbar_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( xbar_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( xbar_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( xbar_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( xbar_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( xbar_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( xbar_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( xbar_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( xbar_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( xbar_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( xbar_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_4_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_4_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_4_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_4_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_4_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_4_r_bits_user ),
       .io_slaves_1_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_slaves_1_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_slaves_1_w_valid( xbar_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( xbar_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_slaves_1_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_slaves_1_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_slaves_1_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_slaves_1_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_slaves_1_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( xbar_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_slaves_1_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_slaves_1_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_slaves_1_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_slaves_1_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_slaves_1_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_0_aw_ready ),
       .io_slaves_0_aw_valid( xbar_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( xbar_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( xbar_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( xbar_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( xbar_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( xbar_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( xbar_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( xbar_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( xbar_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( xbar_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( xbar_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( xbar_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_0_w_ready ),
       .io_slaves_0_w_valid( xbar_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( xbar_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( xbar_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( xbar_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( xbar_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( xbar_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_0_ar_ready ),
       .io_slaves_0_ar_valid( xbar_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( xbar_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( xbar_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( xbar_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( xbar_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( xbar_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( xbar_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( xbar_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( xbar_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( xbar_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( xbar_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( xbar_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( xbar_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_0_r_bits_user )
  );
  NastiRecursiveInterconnect NastiRecursiveInterconnect(.clk(clk), .reset(reset),
       .io_masters_0_aw_ready( NastiRecursiveInterconnect_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( xbar_io_slaves_1_aw_valid ),
       .io_masters_0_aw_bits_addr( xbar_io_slaves_1_aw_bits_addr ),
       .io_masters_0_aw_bits_len( xbar_io_slaves_1_aw_bits_len ),
       .io_masters_0_aw_bits_size( xbar_io_slaves_1_aw_bits_size ),
       .io_masters_0_aw_bits_burst( xbar_io_slaves_1_aw_bits_burst ),
       .io_masters_0_aw_bits_lock( xbar_io_slaves_1_aw_bits_lock ),
       .io_masters_0_aw_bits_cache( xbar_io_slaves_1_aw_bits_cache ),
       .io_masters_0_aw_bits_prot( xbar_io_slaves_1_aw_bits_prot ),
       .io_masters_0_aw_bits_qos( xbar_io_slaves_1_aw_bits_qos ),
       .io_masters_0_aw_bits_region( xbar_io_slaves_1_aw_bits_region ),
       .io_masters_0_aw_bits_id( xbar_io_slaves_1_aw_bits_id ),
       .io_masters_0_aw_bits_user( xbar_io_slaves_1_aw_bits_user ),
       .io_masters_0_w_ready( NastiRecursiveInterconnect_io_masters_0_w_ready ),
       .io_masters_0_w_valid( xbar_io_slaves_1_w_valid ),
       .io_masters_0_w_bits_data( xbar_io_slaves_1_w_bits_data ),
       .io_masters_0_w_bits_last( xbar_io_slaves_1_w_bits_last ),
       .io_masters_0_w_bits_strb( xbar_io_slaves_1_w_bits_strb ),
       .io_masters_0_w_bits_user( xbar_io_slaves_1_w_bits_user ),
       .io_masters_0_b_ready( xbar_io_slaves_1_b_ready ),
       .io_masters_0_b_valid( NastiRecursiveInterconnect_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( NastiRecursiveInterconnect_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( NastiRecursiveInterconnect_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( NastiRecursiveInterconnect_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( NastiRecursiveInterconnect_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( xbar_io_slaves_1_ar_valid ),
       .io_masters_0_ar_bits_addr( xbar_io_slaves_1_ar_bits_addr ),
       .io_masters_0_ar_bits_len( xbar_io_slaves_1_ar_bits_len ),
       .io_masters_0_ar_bits_size( xbar_io_slaves_1_ar_bits_size ),
       .io_masters_0_ar_bits_burst( xbar_io_slaves_1_ar_bits_burst ),
       .io_masters_0_ar_bits_lock( xbar_io_slaves_1_ar_bits_lock ),
       .io_masters_0_ar_bits_cache( xbar_io_slaves_1_ar_bits_cache ),
       .io_masters_0_ar_bits_prot( xbar_io_slaves_1_ar_bits_prot ),
       .io_masters_0_ar_bits_qos( xbar_io_slaves_1_ar_bits_qos ),
       .io_masters_0_ar_bits_region( xbar_io_slaves_1_ar_bits_region ),
       .io_masters_0_ar_bits_id( xbar_io_slaves_1_ar_bits_id ),
       .io_masters_0_ar_bits_user( xbar_io_slaves_1_ar_bits_user ),
       .io_masters_0_r_ready( xbar_io_slaves_1_r_ready ),
       .io_masters_0_r_valid( NastiRecursiveInterconnect_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( NastiRecursiveInterconnect_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( NastiRecursiveInterconnect_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( NastiRecursiveInterconnect_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( NastiRecursiveInterconnect_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( NastiRecursiveInterconnect_io_masters_0_r_bits_user ),
       .io_slaves_2_aw_ready( io_slaves_3_aw_ready ),
       .io_slaves_2_aw_valid( NastiRecursiveInterconnect_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( NastiRecursiveInterconnect_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( NastiRecursiveInterconnect_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( NastiRecursiveInterconnect_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( NastiRecursiveInterconnect_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( NastiRecursiveInterconnect_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( io_slaves_3_w_ready ),
       .io_slaves_2_w_valid( NastiRecursiveInterconnect_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( NastiRecursiveInterconnect_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( NastiRecursiveInterconnect_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( NastiRecursiveInterconnect_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( NastiRecursiveInterconnect_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( NastiRecursiveInterconnect_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( io_slaves_3_b_valid ),
       .io_slaves_2_b_bits_resp( io_slaves_3_b_bits_resp ),
       .io_slaves_2_b_bits_id( io_slaves_3_b_bits_id ),
       .io_slaves_2_b_bits_user( io_slaves_3_b_bits_user ),
       .io_slaves_2_ar_ready( io_slaves_3_ar_ready ),
       .io_slaves_2_ar_valid( NastiRecursiveInterconnect_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( NastiRecursiveInterconnect_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( NastiRecursiveInterconnect_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( NastiRecursiveInterconnect_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( NastiRecursiveInterconnect_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( NastiRecursiveInterconnect_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( NastiRecursiveInterconnect_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( io_slaves_3_r_valid ),
       .io_slaves_2_r_bits_resp( io_slaves_3_r_bits_resp ),
       .io_slaves_2_r_bits_data( io_slaves_3_r_bits_data ),
       .io_slaves_2_r_bits_last( io_slaves_3_r_bits_last ),
       .io_slaves_2_r_bits_id( io_slaves_3_r_bits_id ),
       .io_slaves_2_r_bits_user( io_slaves_3_r_bits_user ),
       .io_slaves_1_aw_ready( io_slaves_2_aw_ready ),
       .io_slaves_1_aw_valid( NastiRecursiveInterconnect_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( NastiRecursiveInterconnect_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( NastiRecursiveInterconnect_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( NastiRecursiveInterconnect_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( NastiRecursiveInterconnect_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( NastiRecursiveInterconnect_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_slaves_2_w_ready ),
       .io_slaves_1_w_valid( NastiRecursiveInterconnect_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( NastiRecursiveInterconnect_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( NastiRecursiveInterconnect_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( NastiRecursiveInterconnect_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( NastiRecursiveInterconnect_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( NastiRecursiveInterconnect_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_slaves_2_b_valid ),
       .io_slaves_1_b_bits_resp( io_slaves_2_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_slaves_2_b_bits_id ),
       .io_slaves_1_b_bits_user( io_slaves_2_b_bits_user ),
       .io_slaves_1_ar_ready( io_slaves_2_ar_ready ),
       .io_slaves_1_ar_valid( NastiRecursiveInterconnect_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( NastiRecursiveInterconnect_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( NastiRecursiveInterconnect_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( NastiRecursiveInterconnect_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( NastiRecursiveInterconnect_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( NastiRecursiveInterconnect_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( NastiRecursiveInterconnect_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_slaves_2_r_valid ),
       .io_slaves_1_r_bits_resp( io_slaves_2_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_slaves_2_r_bits_data ),
       .io_slaves_1_r_bits_last( io_slaves_2_r_bits_last ),
       .io_slaves_1_r_bits_id( io_slaves_2_r_bits_id ),
       .io_slaves_1_r_bits_user( io_slaves_2_r_bits_user ),
       .io_slaves_0_aw_ready( io_slaves_1_aw_ready ),
       .io_slaves_0_aw_valid( NastiRecursiveInterconnect_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( NastiRecursiveInterconnect_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( NastiRecursiveInterconnect_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( NastiRecursiveInterconnect_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( NastiRecursiveInterconnect_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( NastiRecursiveInterconnect_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( NastiRecursiveInterconnect_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( NastiRecursiveInterconnect_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( NastiRecursiveInterconnect_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( NastiRecursiveInterconnect_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( NastiRecursiveInterconnect_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( NastiRecursiveInterconnect_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_slaves_1_w_ready ),
       .io_slaves_0_w_valid( NastiRecursiveInterconnect_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( NastiRecursiveInterconnect_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( NastiRecursiveInterconnect_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( NastiRecursiveInterconnect_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( NastiRecursiveInterconnect_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( NastiRecursiveInterconnect_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_slaves_1_b_valid ),
       .io_slaves_0_b_bits_resp( io_slaves_1_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_slaves_1_b_bits_id ),
       .io_slaves_0_b_bits_user( io_slaves_1_b_bits_user ),
       .io_slaves_0_ar_ready( io_slaves_1_ar_ready ),
       .io_slaves_0_ar_valid( NastiRecursiveInterconnect_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( NastiRecursiveInterconnect_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( NastiRecursiveInterconnect_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( NastiRecursiveInterconnect_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( NastiRecursiveInterconnect_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( NastiRecursiveInterconnect_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( NastiRecursiveInterconnect_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( NastiRecursiveInterconnect_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( NastiRecursiveInterconnect_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( NastiRecursiveInterconnect_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( NastiRecursiveInterconnect_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( NastiRecursiveInterconnect_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( NastiRecursiveInterconnect_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_slaves_1_r_valid ),
       .io_slaves_0_r_bits_resp( io_slaves_1_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_slaves_1_r_bits_data ),
       .io_slaves_0_r_bits_last( io_slaves_1_r_bits_last ),
       .io_slaves_0_r_bits_id( io_slaves_1_r_bits_id ),
       .io_slaves_0_r_bits_user( io_slaves_1_r_bits_user )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [2:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [2:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[2:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  wire T1;
  wire T2;
  wire T3;
  reg  last_grant;
  wire T52;
  wire T4;
  wire T5;
  reg  lockIdx;
  wire T53;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  reg  locked;
  wire T54;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire[1:0] T19;
  reg [1:0] R20;
  wire[1:0] T55;
  wire[1:0] T21;
  wire[127:0] T22;
  wire T23;
  wire[16:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[1:0] T27;
  wire[2:0] T28;
  wire[25:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R20 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = T2 ? 1'h1 : T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign T2 = io_in_1_valid & T3;
  assign T3 = last_grant < 1'h1;
  assign T52 = reset ? 1'h0 : T4;
  assign T4 = T5 ? chosen : last_grant;
  assign T5 = io_out_ready & io_out_valid;
  assign T53 = reset ? 1'h1 : T6;
  assign T6 = T9 ? T7 : lockIdx;
  assign T7 = T8 == 1'h0;
  assign T8 = io_in_0_ready & io_in_0_valid;
  assign T9 = T11 & T10;
  assign T10 = locked ^ 1'h1;
  assign T11 = T14 & T12;
  assign T12 = io_out_bits_is_builtin_type & T13;
  assign T13 = 3'h3 == io_out_bits_a_type;
  assign T14 = io_out_ready & io_out_valid;
  assign T54 = reset ? 1'h0 : T15;
  assign T15 = T17 ? 1'h0 : T16;
  assign T16 = T9 ? 1'h1 : locked;
  assign T17 = T14 & T18;
  assign T18 = T19 == 2'h0;
  assign T19 = R20 + 2'h1;
  assign T55 = reset ? 2'h0 : T21;
  assign T21 = T11 ? T19 : R20;
  assign io_out_bits_data = T22;
  assign T22 = T23 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T23 = chosen;
  assign io_out_bits_union = T24;
  assign T24 = T23 ? io_in_1_bits_union : io_in_0_bits_union;
  assign io_out_bits_a_type = T25;
  assign T25 = T23 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_is_builtin_type = T26;
  assign T26 = T23 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_addr_beat = T27;
  assign T27 = T23 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_bits_client_xact_id = T28;
  assign T28 = T23 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T29;
  assign T29 = T23 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_valid = T30;
  assign T30 = T23 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T41 : T33;
  assign T33 = T40 | T34;
  assign T34 = T35 ^ 1'h1;
  assign T35 = T38 | T36;
  assign T36 = io_in_1_valid & T37;
  assign T37 = last_grant < 1'h1;
  assign T38 = io_in_0_valid & T39;
  assign T39 = last_grant < 1'h0;
  assign T40 = last_grant < 1'h0;
  assign T41 = lockIdx == 1'h0;
  assign io_in_1_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = locked ? T51 : T44;
  assign T44 = T48 | T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = T47 | io_in_0_valid;
  assign T47 = T38 | T36;
  assign T48 = T50 & T49;
  assign T49 = last_grant < 1'h1;
  assign T50 = T38 ^ 1'h1;
  assign T51 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T5) begin
      last_grant <= chosen;
    end
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T9) begin
      lockIdx <= T7;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T17) begin
      locked <= 1'h0;
    end else if(T9) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R20 <= 2'h0;
    end else if(T11) begin
      R20 <= T19;
    end
  end
endmodule

module ReorderQueue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_data,
    input [2:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [2:0] io_deq_tag,
    output io_deq_data,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_5;
  wire T1;
  reg  roq_free_5;
  wire T122;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[7:0] T6;
  wire[2:0] T7;
  wire[2:0] roq_enq_addr;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  reg  roq_free_4;
  wire T123;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[2:0] T19;
  wire[2:0] roq_deq_addr;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire roq_matches_4;
  wire T24;
  wire T25;
  reg [2:0] roq_tags_4;
  wire[2:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[2:0] T30;
  wire roq_matches_3;
  wire T31;
  wire T32;
  reg [2:0] roq_tags_3;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire roq_matches_2;
  wire T36;
  wire T37;
  reg [2:0] roq_tags_2;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire roq_matches_1;
  wire T41;
  wire T42;
  reg [2:0] roq_tags_1;
  wire[2:0] T43;
  wire T44;
  wire T45;
  wire roq_matches_0;
  wire T46;
  wire T47;
  reg [2:0] roq_tags_0;
  wire[2:0] T48;
  wire T49;
  wire T50;
  reg  roq_free_3;
  wire T124;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  reg  roq_free_2;
  wire T125;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  roq_free_1;
  wire T126;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  reg  roq_free_0;
  wire T127;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [2:0] roq_tags_5;
  wire[2:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  reg  roq_data_0;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[2:0] T93;
  reg  roq_data_1;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[2:0] T98;
  wire T99;
  reg  roq_data_2;
  wire T100;
  wire T101;
  wire T102;
  reg  roq_data_3;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  reg  roq_data_4;
  wire T109;
  wire T110;
  wire T111;
  reg  roq_data_5;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_data_0 = {1{$random}};
    roq_data_1 = {1{$random}};
    roq_data_2 = {1{$random}};
    roq_data_3 = {1{$random}};
    roq_data_4 = {1{$random}};
    roq_data_5 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T82 | roq_matches_5;
  assign roq_matches_5 = T78 & T1;
  assign T1 = roq_free_5 ^ 1'h1;
  assign T122 = reset ? 1'h1 : T2;
  assign T2 = T76 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_5;
  assign T4 = T75 & T5;
  assign T5 = T6[3'h5:3'h5];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 3'h0 : T8;
  assign T8 = roq_free_1 ? 3'h1 : T9;
  assign T9 = roq_free_2 ? 3'h2 : T10;
  assign T10 = roq_free_3 ? 3'h3 : T11;
  assign T11 = roq_free_4 ? 3'h4 : 3'h5;
  assign T123 = reset ? 1'h1 : T12;
  assign T12 = T16 ? 1'h1 : T13;
  assign T13 = T14 ? 1'h0 : roq_free_4;
  assign T14 = T75 & T15;
  assign T15 = T6[3'h4:3'h4];
  assign T16 = io_deq_valid & T17;
  assign T17 = T18[3'h4:3'h4];
  assign T18 = 1'h1 << T19;
  assign T19 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 3'h0 : T20;
  assign T20 = roq_matches_1 ? 3'h1 : T21;
  assign T21 = roq_matches_2 ? 3'h2 : T22;
  assign T22 = roq_matches_3 ? 3'h3 : T23;
  assign T23 = roq_matches_4 ? 3'h4 : 3'h5;
  assign roq_matches_4 = T25 & T24;
  assign T24 = roq_free_4 ^ 1'h1;
  assign T25 = roq_tags_4 == io_deq_tag;
  assign T26 = T27 ? io_enq_bits_tag : roq_tags_4;
  assign T27 = T75 & T28;
  assign T28 = T29[3'h4:3'h4];
  assign T29 = 1'h1 << T30;
  assign T30 = roq_enq_addr;
  assign roq_matches_3 = T32 & T31;
  assign T31 = roq_free_3 ^ 1'h1;
  assign T32 = roq_tags_3 == io_deq_tag;
  assign T33 = T34 ? io_enq_bits_tag : roq_tags_3;
  assign T34 = T75 & T35;
  assign T35 = T29[2'h3:2'h3];
  assign roq_matches_2 = T37 & T36;
  assign T36 = roq_free_2 ^ 1'h1;
  assign T37 = roq_tags_2 == io_deq_tag;
  assign T38 = T39 ? io_enq_bits_tag : roq_tags_2;
  assign T39 = T75 & T40;
  assign T40 = T29[2'h2:2'h2];
  assign roq_matches_1 = T42 & T41;
  assign T41 = roq_free_1 ^ 1'h1;
  assign T42 = roq_tags_1 == io_deq_tag;
  assign T43 = T44 ? io_enq_bits_tag : roq_tags_1;
  assign T44 = T75 & T45;
  assign T45 = T29[1'h1:1'h1];
  assign roq_matches_0 = T47 & T46;
  assign T46 = roq_free_0 ^ 1'h1;
  assign T47 = roq_tags_0 == io_deq_tag;
  assign T48 = T49 ? io_enq_bits_tag : roq_tags_0;
  assign T49 = T75 & T50;
  assign T50 = T29[1'h0:1'h0];
  assign T124 = reset ? 1'h1 : T51;
  assign T51 = T55 ? 1'h1 : T52;
  assign T52 = T53 ? 1'h0 : roq_free_3;
  assign T53 = T75 & T54;
  assign T54 = T6[2'h3:2'h3];
  assign T55 = io_deq_valid & T56;
  assign T56 = T18[2'h3:2'h3];
  assign T125 = reset ? 1'h1 : T57;
  assign T57 = T61 ? 1'h1 : T58;
  assign T58 = T59 ? 1'h0 : roq_free_2;
  assign T59 = T75 & T60;
  assign T60 = T6[2'h2:2'h2];
  assign T61 = io_deq_valid & T62;
  assign T62 = T18[2'h2:2'h2];
  assign T126 = reset ? 1'h1 : T63;
  assign T63 = T67 ? 1'h1 : T64;
  assign T64 = T65 ? 1'h0 : roq_free_1;
  assign T65 = T75 & T66;
  assign T66 = T6[1'h1:1'h1];
  assign T67 = io_deq_valid & T68;
  assign T68 = T18[1'h1:1'h1];
  assign T127 = reset ? 1'h1 : T69;
  assign T69 = T73 ? 1'h1 : T70;
  assign T70 = T71 ? 1'h0 : roq_free_0;
  assign T71 = T75 & T72;
  assign T72 = T6[1'h0:1'h0];
  assign T73 = io_deq_valid & T74;
  assign T74 = T18[1'h0:1'h0];
  assign T75 = io_enq_valid & io_enq_ready;
  assign T76 = io_deq_valid & T77;
  assign T77 = T18[3'h5:3'h5];
  assign T78 = roq_tags_5 == io_deq_tag;
  assign T79 = T80 ? io_enq_bits_tag : roq_tags_5;
  assign T80 = T75 & T81;
  assign T81 = T29[3'h5:3'h5];
  assign T82 = T83 | roq_matches_4;
  assign T83 = T84 | roq_matches_3;
  assign T84 = T85 | roq_matches_2;
  assign T85 = roq_matches_0 | roq_matches_1;
  assign io_deq_data = T86;
  assign T86 = T116 ? T108 : T87;
  assign T87 = T107 ? T99 : T88;
  assign T88 = T97 ? roq_data_1 : roq_data_0;
  assign T89 = T90 ? io_enq_bits_data : roq_data_0;
  assign T90 = T75 & T91;
  assign T91 = T92[1'h0:1'h0];
  assign T92 = 1'h1 << T93;
  assign T93 = roq_enq_addr;
  assign T94 = T95 ? io_enq_bits_data : roq_data_1;
  assign T95 = T75 & T96;
  assign T96 = T92[1'h1:1'h1];
  assign T97 = T98[1'h0:1'h0];
  assign T98 = roq_deq_addr;
  assign T99 = T106 ? roq_data_3 : roq_data_2;
  assign T100 = T101 ? io_enq_bits_data : roq_data_2;
  assign T101 = T75 & T102;
  assign T102 = T92[2'h2:2'h2];
  assign T103 = T104 ? io_enq_bits_data : roq_data_3;
  assign T104 = T75 & T105;
  assign T105 = T92[2'h3:2'h3];
  assign T106 = T98[1'h0:1'h0];
  assign T107 = T98[1'h1:1'h1];
  assign T108 = T115 ? roq_data_5 : roq_data_4;
  assign T109 = T110 ? io_enq_bits_data : roq_data_4;
  assign T110 = T75 & T111;
  assign T111 = T92[3'h4:3'h4];
  assign T112 = T113 ? io_enq_bits_data : roq_data_5;
  assign T113 = T75 & T114;
  assign T114 = T92[3'h5:3'h5];
  assign T115 = T98[1'h0:1'h0];
  assign T116 = T98[2'h2:2'h2];
  assign io_enq_ready = T117;
  assign T117 = T118 | roq_free_5;
  assign T118 = T119 | roq_free_4;
  assign T119 = T120 | roq_free_3;
  assign T120 = T121 | roq_free_2;
  assign T121 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T76) begin
      roq_free_5 <= 1'h1;
    end else if(T4) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T16) begin
      roq_free_4 <= 1'h1;
    end else if(T14) begin
      roq_free_4 <= 1'h0;
    end
    if(T27) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T34) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T39) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T44) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T49) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T55) begin
      roq_free_3 <= 1'h1;
    end else if(T53) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T61) begin
      roq_free_2 <= 1'h1;
    end else if(T59) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T67) begin
      roq_free_1 <= 1'h1;
    end else if(T65) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T73) begin
      roq_free_0 <= 1'h1;
    end else if(T71) begin
      roq_free_0 <= 1'h0;
    end
    if(T80) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T90) begin
      roq_data_0 <= io_enq_bits_data;
    end
    if(T95) begin
      roq_data_1 <= io_enq_bits_data;
    end
    if(T101) begin
      roq_data_2 <= io_enq_bits_data;
    end
    if(T104) begin
      roq_data_3 <= io_enq_bits_data;
    end
    if(T110) begin
      roq_data_4 <= io_enq_bits_data;
    end
    if(T113) begin
      roq_data_5 <= io_enq_bits_data;
    end
  end
endmodule

module ClientTileLinkIOUnwrapper(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [2:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[2:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_in_probe_ready,
    output io_in_probe_valid,
    //output[25:0] io_in_probe_bits_addr_block
    //output[1:0] io_in_probe_bits_p_type
    output io_in_release_ready,
    input  io_in_release_valid,
    input [1:0] io_in_release_bits_addr_beat,
    input [25:0] io_in_release_bits_addr_block,
    input [2:0] io_in_release_bits_client_xact_id,
    input  io_in_release_bits_voluntary,
    input [2:0] io_in_release_bits_r_type,
    input [127:0] io_in_release_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire rel_roq_enq;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire acq_roq_enq;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire[127:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire T36;
  wire[1:0] T37;
  wire[2:0] T38;
  wire[25:0] T39;
  wire T40;
  wire acq_roq_ready;
  wire T41;
  wire[127:0] T42;
  wire[16:0] T43;
  wire[16:0] T44;
  wire[15:0] T45;
  wire[2:0] T46;
  wire T47;
  wire[1:0] T48;
  wire[2:0] T49;
  wire[25:0] T50;
  wire T51;
  wire rel_roq_ready;
  wire T52;
  wire T53;
  wire[127:0] T54;
  wire[127:0] rel_grant_data;
  wire[127:0] acq_grant_data;
  wire[3:0] T55;
  wire[3:0] rel_grant_g_type;
  wire[3:0] T56;
  wire[3:0] acq_grant_g_type;
  wire[3:0] T57;
  wire T58;
  wire rel_grant_is_builtin_type;
  wire acq_grant_is_builtin_type;
  wire T59;
  wire rel_grant_manager_xact_id;
  wire acq_grant_manager_xact_id;
  wire[2:0] T60;
  wire[2:0] rel_grant_client_xact_id;
  wire[2:0] acq_grant_client_xact_id;
  wire[1:0] T61;
  wire[1:0] rel_grant_addr_beat;
  wire[1:0] acq_grant_addr_beat;
  wire T62;
  wire acqArb_io_in_1_ready;
  wire acqArb_io_in_0_ready;
  wire acqArb_io_out_valid;
  wire[25:0] acqArb_io_out_bits_addr_block;
  wire[2:0] acqArb_io_out_bits_client_xact_id;
  wire[1:0] acqArb_io_out_bits_addr_beat;
  wire acqArb_io_out_bits_is_builtin_type;
  wire[2:0] acqArb_io_out_bits_a_type;
  wire[16:0] acqArb_io_out_bits_union;
  wire[127:0] acqArb_io_out_bits_data;
  wire acqRoq_io_enq_ready;
  wire acqRoq_io_deq_data;
  wire acqRoq_io_deq_matches;
  wire relRoq_io_enq_ready;
  wire relRoq_io_deq_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_in_probe_bits_p_type = {1{$random}};
//  assign io_in_probe_bits_addr_block = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = T7 & T1;
  assign T1 = T3 | T2;
  assign T2 = io_out_grant_bits_addr_beat == 2'h3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = io_out_grant_bits_is_builtin_type ? T6 : T5;
  assign T5 = 4'h0 == io_out_grant_bits_g_type;
  assign T6 = 4'h5 == io_out_grant_bits_g_type;
  assign T7 = io_out_grant_ready & io_out_grant_valid;
  assign T8 = T16 & rel_roq_enq;
  assign rel_roq_enq = T10 | T9;
  assign T9 = io_in_release_bits_addr_beat == 2'h0;
  assign T10 = T11 ^ 1'h1;
  assign T11 = T13 | T12;
  assign T12 = 3'h2 == io_in_release_bits_r_type;
  assign T13 = T15 | T14;
  assign T14 = 3'h1 == io_in_release_bits_r_type;
  assign T15 = 3'h0 == io_in_release_bits_r_type;
  assign T16 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T17 = T24 & T18;
  assign T18 = T20 | T19;
  assign T19 = io_out_grant_bits_addr_beat == 2'h3;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_out_grant_bits_is_builtin_type ? T23 : T22;
  assign T22 = 4'h0 == io_out_grant_bits_g_type;
  assign T23 = 4'h5 == io_out_grant_bits_g_type;
  assign T24 = io_out_grant_ready & io_out_grant_valid;
  assign T25 = T30 & acq_roq_enq;
  assign acq_roq_enq = T27 | T26;
  assign T26 = io_in_acquire_bits_addr_beat == 2'h0;
  assign T27 = T28 ^ 1'h1;
  assign T28 = io_in_acquire_bits_is_builtin_type & T29;
  assign T29 = 3'h3 == io_in_acquire_bits_a_type;
  assign T30 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T31 = io_in_acquire_bits_data;
  assign T32 = T33;
  assign T33 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : 17'h1c1;
  assign T34 = T35;
  assign T35 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T36 = 1'h1;
  assign T37 = io_in_acquire_bits_addr_beat;
  assign T38 = io_in_acquire_bits_client_xact_id;
  assign T39 = io_in_acquire_bits_addr_block;
  assign T40 = io_in_acquire_valid & acq_roq_ready;
  assign acq_roq_ready = T41 | acqRoq_io_enq_ready;
  assign T41 = acq_roq_enq ^ 1'h1;
  assign T42 = io_in_release_bits_data;
  assign T43 = T44;
  assign T44 = {T45, 1'h1};
  assign T45 = 16'hffff;
  assign T46 = 3'h3;
  assign T47 = 1'h1;
  assign T48 = io_in_release_bits_addr_beat;
  assign T49 = io_in_release_bits_client_xact_id;
  assign T50 = io_in_release_bits_addr_block;
  assign T51 = io_in_release_valid & rel_roq_ready;
  assign rel_roq_ready = T52 | relRoq_io_enq_ready;
  assign T52 = rel_roq_enq ^ 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_in_release_ready = T53;
  assign T53 = rel_roq_ready & acqArb_io_in_1_ready;
  assign io_in_probe_valid = 1'h0;
  assign io_in_grant_bits_data = T54;
  assign T54 = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
  assign rel_grant_data = io_out_grant_bits_data;
  assign acq_grant_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = T55;
  assign T55 = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign rel_grant_g_type = T56;
  assign T56 = relRoq_io_deq_data ? 4'h0 : io_out_grant_bits_g_type;
  assign acq_grant_g_type = T57;
  assign T57 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign io_in_grant_bits_is_builtin_type = T58;
  assign T58 = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign rel_grant_is_builtin_type = 1'h1;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign io_in_grant_bits_manager_xact_id = T59;
  assign T59 = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = T60;
  assign T60 = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = T61;
  assign T61 = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = T62;
  assign T62 = acq_roq_ready & acqArb_io_in_0_ready;
  LockingRRArbiter_4 acqArb(.clk(clk), .reset(reset),
       .io_in_1_ready( acqArb_io_in_1_ready ),
       .io_in_1_valid( T51 ),
       .io_in_1_bits_addr_block( T50 ),
       .io_in_1_bits_client_xact_id( T49 ),
       .io_in_1_bits_addr_beat( T48 ),
       .io_in_1_bits_is_builtin_type( T47 ),
       .io_in_1_bits_a_type( T46 ),
       .io_in_1_bits_union( T43 ),
       .io_in_1_bits_data( T42 ),
       .io_in_0_ready( acqArb_io_in_0_ready ),
       .io_in_0_valid( T40 ),
       .io_in_0_bits_addr_block( T39 ),
       .io_in_0_bits_client_xact_id( T38 ),
       .io_in_0_bits_addr_beat( T37 ),
       .io_in_0_bits_is_builtin_type( T36 ),
       .io_in_0_bits_a_type( T34 ),
       .io_in_0_bits_union( T32 ),
       .io_in_0_bits_data( T31 ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( acqArb_io_out_valid ),
       .io_out_bits_addr_block( acqArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( acqArb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( acqArb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( acqArb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( acqArb_io_out_bits_a_type ),
       .io_out_bits_union( acqArb_io_out_bits_union ),
       .io_out_bits_data( acqArb_io_out_bits_data )
       //.io_chosen(  )
  );
  ReorderQueue_0 acqRoq(.clk(clk), .reset(reset),
       .io_enq_ready( acqRoq_io_enq_ready ),
       .io_enq_valid( T25 ),
       .io_enq_bits_data( io_in_acquire_bits_is_builtin_type ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T17 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( acqRoq_io_deq_data ),
       .io_deq_matches( acqRoq_io_deq_matches )
  );
  ReorderQueue_0 relRoq(.clk(clk), .reset(reset),
       .io_enq_ready( relRoq_io_enq_ready ),
       .io_enq_valid( T8 ),
       .io_enq_bits_data( io_in_release_bits_voluntary ),
       .io_enq_bits_tag( io_in_release_bits_client_xact_id ),
       .io_deq_valid( T0 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( relRoq_io_deq_data )
       //.io_deq_matches(  )
  );
endmodule

module TileLinkIONarrower(input clk, input reset,
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [2:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[2:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[2:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[11:0] io_out_acquire_bits_union,
    output[63:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [2:0] io_out_grant_bits_addr_beat,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [63:0] io_out_grant_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg[0:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  wire[7:0] T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[15:0] T37;
  wire[15:0] T38;
  wire[7:0] T39;
  wire[7:0] T303;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire[3:0] T43;
  wire[7:0] T44;
  wire[7:0] T304;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[7:0] T49;
  wire[15:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[15:0] T58;
  wire[15:0] T59;
  wire[7:0] T60;
  wire[7:0] T305;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire[3:0] T64;
  wire[7:0] T65;
  wire[7:0] T306;
  wire T66;
  wire T67;
  wire T68;
  wire[1:0] T307;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[31:0] T78;
  wire[5:0] T79;
  wire[3:0] T80;
  wire T81;
  wire T82;
  reg  R83;
  wire T308;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  reg  R91;
  wire T309;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  reg  R103;
  wire T310;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg  R108;
  wire T311;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire[63:0] T312;
  wire[127:0] T115;
  wire[127:0] T116;
  wire[127:0] T117;
  wire[127:0] T118;
  wire[127:0] T313;
  wire[63:0] T119;
  wire[127:0] T314;
  wire[63:0] T120;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire[127:0] T315;
  wire[63:0] T128;
  wire T129;
  wire[127:0] T316;
  wire[63:0] T130;
  wire[63:0] T131;
  reg [127:0] R132;
  wire[127:0] T133;
  wire[127:0] T134;
  wire[127:0] T317;
  wire[63:0] T135;
  wire[11:0] T318;
  wire[16:0] T136;
  wire[16:0] T137;
  wire[16:0] T138;
  wire[16:0] T139;
  wire[16:0] T319;
  wire[11:0] T140;
  wire[11:0] T141;
  wire[5:0] T142;
  wire T143;
  wire[5:0] T144;
  wire[2:0] T145;
  wire[2:0] T146;
  wire[31:0] T147;
  wire[5:0] T148;
  wire[3:0] T149;
  wire[16:0] T320;
  wire[11:0] T150;
  wire[11:0] T321;
  wire[8:0] T151;
  wire[7:0] T152;
  wire[7:0] T153;
  wire T154;
  wire[7:0] T155;
  wire T156;
  wire[16:0] T322;
  wire[11:0] T157;
  wire[11:0] T323;
  wire[8:0] T158;
  wire[5:0] T159;
  wire T160;
  wire[16:0] T324;
  wire[11:0] T161;
  wire[11:0] T325;
  wire[8:0] T162;
  wire[7:0] T163;
  reg [15:0] R164;
  wire[15:0] T165;
  wire[15:0] T166;
  wire[15:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[15:0] T175;
  wire[15:0] T176;
  wire[7:0] T177;
  wire[7:0] T326;
  wire T178;
  wire[1:0] T179;
  wire T180;
  wire[3:0] T181;
  wire[7:0] T182;
  wire[7:0] T327;
  wire T183;
  wire T184;
  wire T185;
  wire[15:0] T328;
  wire[7:0] T186;
  wire[2:0] T187;
  wire[2:0] T188;
  wire[2:0] T189;
  wire[2:0] T190;
  wire[2:0] T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[2:0] T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[2:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[2:0] T206;
  wire[2:0] T329;
  wire[2:0] T207;
  wire[2:0] T208;
  wire[31:0] T209;
  wire[5:0] T210;
  wire[3:0] T211;
  wire[2:0] T212;
  wire[2:0] T213;
  wire T330;
  wire T331;
  wire[2:0] T215;
  wire[2:0] T216;
  wire[2:0] T217;
  reg [1:0] R218;
  wire[1:0] T219;
  wire[2:0] T220;
  wire[2:0] T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire[2:0] T224;
  wire[2:0] T225;
  wire[2:0] T226;
  wire[2:0] T227;
  reg [2:0] R228;
  wire[2:0] T229;
  wire[25:0] T230;
  wire[25:0] T231;
  wire[25:0] T232;
  wire[25:0] T233;
  wire[25:0] T234;
  wire[25:0] T235;
  wire[25:0] T236;
  wire[25:0] T237;
  reg [25:0] R238;
  wire[25:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[127:0] T247;
  wire[127:0] T248;
  wire[127:0] T332;
  wire[127:0] T249;
  wire[127:0] T333;
  wire[190:0] T250;
  wire[6:0] T251;
  wire[127:0] T252;
  wire[127:0] T253;
  wire[127:0] T254;
  reg [63:0] R255;
  wire[63:0] T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  wire T260;
  reg [63:0] R261;
  wire[63:0] T262;
  wire T263;
  wire T264;
  wire[3:0] T265;
  wire[3:0] T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  reg  R277;
  wire T278;
  wire[2:0] T279;
  wire[2:0] T280;
  wire[2:0] T281;
  wire[2:0] T282;
  reg [2:0] R283;
  wire[2:0] T284;
  wire[1:0] T334;
  wire[2:0] T285;
  wire[2:0] T286;
  wire[2:0] T335;
  wire[1:0] T287;
  wire[1:0] T288;
  wire[2:0] T336;
  wire[1:0] T289;
  reg [1:0] R290;
  wire[1:0] T337;
  wire[1:0] T291;
  wire[1:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire ReorderQueue_io_enq_ready;
  wire ReorderQueue_io_deq_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T19 = 1'b0;
    R83 = {1{$random}};
    R91 = {1{$random}};
    R103 = {1{$random}};
    R108 = {1{$random}};
    R132 = {4{$random}};
    R164 = {1{$random}};
    R218 = {1{$random}};
    R228 = {1{$random}};
    R238 = {1{$random}};
    R255 = {2{$random}};
    R261 = {2{$random}};
    R277 = {1{$random}};
    R283 = {1{$random}};
    R290 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T15 | T3;
  assign T3 = T14 ? 1'h1 : T4;
  assign T4 = T13 ? 1'h1 : T5;
  assign T5 = T12 ? 1'h1 : T6;
  assign T6 = T11 ? 1'h1 : T7;
  assign T7 = T10 ? 1'h1 : T8;
  assign T8 = T9 == 3'h3;
  assign T9 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T10 = T9 == 3'h2;
  assign T11 = T9 == 3'h5;
  assign T12 = T9 == 3'h1;
  assign T13 = T9 == 3'h4;
  assign T14 = T9 == 3'h0;
  assign T15 = T18 | T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = io_in_acquire_bits_a_type == 3'h0;
  assign T18 = io_in_acquire_valid ^ 1'h1;
  assign T20 = T21 | reset;
  assign T21 = T70 | T22;
  assign T22 = T23 <= 2'h1;
  assign T23 = T307 + T24;
  assign T24 = {1'h0, T25};
  assign T25 = T26[1'h1:1'h1];
  assign T26 = {T48, T27};
  assign T27 = T28 != 8'h0;
  assign T28 = T29[3'h7:1'h0];
  assign T29 = T46 ? T37 : T30;
  assign T30 = T32 ? T31 : 16'h0;
  assign T31 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T32 = T35 | T33;
  assign T33 = io_in_acquire_bits_is_builtin_type & T34;
  assign T34 = io_in_acquire_bits_a_type == 3'h2;
  assign T35 = io_in_acquire_bits_is_builtin_type & T36;
  assign T36 = io_in_acquire_bits_a_type == 3'h3;
  assign T37 = T38;
  assign T38 = {T44, T39};
  assign T39 = 8'h0 - T303;
  assign T303 = {7'h0, T40};
  assign T40 = T41[1'h0:1'h0];
  assign T41 = 1'h1 << T42;
  assign T42 = T43[2'h3:2'h3];
  assign T43 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T44 = 8'h0 - T304;
  assign T304 = {7'h0, T45};
  assign T45 = T41[1'h1:1'h1];
  assign T46 = io_in_acquire_bits_is_builtin_type & T47;
  assign T47 = io_in_acquire_bits_a_type == 3'h4;
  assign T48 = T49 != 8'h0;
  assign T49 = T50[4'hf:4'h8];
  assign T50 = T67 ? T58 : T51;
  assign T51 = T53 ? T52 : 16'h0;
  assign T52 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T53 = T56 | T54;
  assign T54 = io_in_acquire_bits_is_builtin_type & T55;
  assign T55 = io_in_acquire_bits_a_type == 3'h2;
  assign T56 = io_in_acquire_bits_is_builtin_type & T57;
  assign T57 = io_in_acquire_bits_a_type == 3'h3;
  assign T58 = T59;
  assign T59 = {T65, T60};
  assign T60 = 8'h0 - T305;
  assign T305 = {7'h0, T61};
  assign T61 = T62[1'h0:1'h0];
  assign T62 = 1'h1 << T63;
  assign T63 = T64[2'h3:2'h3];
  assign T64 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T65 = 8'h0 - T306;
  assign T306 = {7'h0, T66};
  assign T66 = T62[1'h1:1'h1];
  assign T67 = io_in_acquire_bits_is_builtin_type & T68;
  assign T68 = io_in_acquire_bits_a_type == 3'h4;
  assign T307 = {1'h0, T69};
  assign T69 = T26[1'h0:1'h0];
  assign T70 = T73 | T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = io_in_acquire_bits_a_type == 3'h2;
  assign T73 = io_in_acquire_valid ^ 1'h1;
  assign T74 = T76 & T75;
  assign T75 = io_out_grant_bits_g_type == 4'h4;
  assign T76 = io_out_grant_ready & io_out_grant_valid;
  assign T77 = T78[2'h3:2'h3];
  assign T78 = {io_in_acquire_bits_addr_block, T79};
  assign T79 = {io_in_acquire_bits_addr_beat, T80};
  assign T80 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T81 = T95 & T82;
  assign T82 = R83 ^ 1'h1;
  assign T308 = reset ? 1'h0 : T84;
  assign T84 = T89 ? 1'h0 : T85;
  assign T85 = T86 ? 1'h1 : R83;
  assign T86 = T88 & T87;
  assign T87 = io_in_acquire_bits_a_type == 3'h3;
  assign T88 = io_in_acquire_ready & io_in_acquire_valid;
  assign T89 = T94 & T90;
  assign T90 = R91 == 1'h1;
  assign T309 = reset ? 1'h0 : T92;
  assign T92 = T94 ? T93 : R91;
  assign T93 = R91 + 1'h1;
  assign T94 = R83 & io_out_acquire_ready;
  assign T95 = T96 & io_out_acquire_ready;
  assign T96 = T17 & io_in_acquire_valid;
  assign io_out_grant_ready = T97;
  assign T97 = T102 & T98;
  assign T98 = T99 | io_in_grant_ready;
  assign T99 = io_out_grant_bits_is_builtin_type ? T101 : T100;
  assign T100 = 4'h0 == io_out_grant_bits_g_type;
  assign T101 = 4'h5 == io_out_grant_bits_g_type;
  assign T102 = R103 ^ 1'h1;
  assign T310 = reset ? 1'h0 : T104;
  assign T104 = T114 ? 1'h0 : T105;
  assign T105 = T106 ? 1'h1 : R103;
  assign T106 = T111 & T107;
  assign T107 = R108 == 1'h1;
  assign T311 = reset ? 1'h0 : T109;
  assign T109 = T111 ? T110 : R108;
  assign T110 = R108 + 1'h1;
  assign T111 = T113 & T112;
  assign T112 = R103 ^ 1'h1;
  assign T113 = io_out_grant_valid & T99;
  assign T114 = io_in_grant_ready & R103;
  assign io_out_acquire_bits_data = T312;
  assign T312 = T115[6'h3f:1'h0];
  assign T115 = R83 ? T316 : T116;
  assign T116 = T129 ? T315 : T117;
  assign T117 = T72 ? T314 : T118;
  assign T118 = T17 ? T313 : io_in_acquire_bits_data;
  assign T313 = {64'h0, T119};
  assign T119 = 64'h0;
  assign T314 = {64'h0, T120};
  assign T120 = T121;
  assign T121 = T125 | T122;
  assign T122 = T124 ? T123 : 64'h0;
  assign T123 = io_in_acquire_bits_data[7'h7f:7'h40];
  assign T124 = T26[1'h1:1'h1];
  assign T125 = T127 ? T126 : 64'h0;
  assign T126 = io_in_acquire_bits_data[6'h3f:1'h0];
  assign T127 = T26[1'h0:1'h0];
  assign T315 = {64'h0, T128};
  assign T128 = 64'h0;
  assign T129 = io_in_acquire_bits_a_type == 3'h1;
  assign T316 = {64'h0, T130};
  assign T130 = T131;
  assign T131 = R132[6'h3f:1'h0];
  assign T133 = T94 ? T317 : T134;
  assign T134 = T86 ? io_in_acquire_bits_data : R132;
  assign T317 = {64'h0, T135};
  assign T135 = R132 >> 7'h40;
  assign io_out_acquire_bits_union = T318;
  assign T318 = T136[4'hb:1'h0];
  assign T136 = R83 ? T324 : T137;
  assign T137 = T129 ? T322 : T138;
  assign T138 = T72 ? T320 : T139;
  assign T139 = T17 ? T319 : io_in_acquire_bits_union;
  assign T319 = {5'h0, T140};
  assign T140 = T141;
  assign T141 = {T144, T142};
  assign T142 = {5'h0, T143};
  assign T143 = io_in_acquire_bits_union[1'h0:1'h0];
  assign T144 = {T146, T145};
  assign T145 = io_in_acquire_bits_union[4'h8:3'h6];
  assign T146 = T147[2'h2:1'h0];
  assign T147 = {io_in_acquire_bits_addr_block, T148};
  assign T148 = {io_in_acquire_bits_addr_beat, T149};
  assign T149 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T320 = {5'h0, T150};
  assign T150 = T321;
  assign T321 = {3'h0, T151};
  assign T151 = {T152, 1'h1};
  assign T152 = T155 | T153;
  assign T153 = T154 ? T49 : 8'h0;
  assign T154 = T26[1'h1:1'h1];
  assign T155 = T156 ? T28 : 8'h0;
  assign T156 = T26[1'h0:1'h0];
  assign T322 = {5'h0, T157};
  assign T157 = T323;
  assign T323 = {3'h0, T158};
  assign T158 = {3'h7, T159};
  assign T159 = {5'h0, T160};
  assign T160 = io_in_acquire_bits_union[1'h0:1'h0];
  assign T324 = {5'h0, T161};
  assign T161 = T325;
  assign T325 = {3'h0, T162};
  assign T162 = {T163, 1'h1};
  assign T163 = R164[3'h7:1'h0];
  assign T165 = T94 ? T328 : T166;
  assign T166 = T86 ? T167 : R164;
  assign T167 = T184 ? T175 : T168;
  assign T168 = T170 ? T169 : 16'h0;
  assign T169 = io_in_acquire_bits_union[5'h10:1'h1];
  assign T170 = T173 | T171;
  assign T171 = io_in_acquire_bits_is_builtin_type & T172;
  assign T172 = io_in_acquire_bits_a_type == 3'h2;
  assign T173 = io_in_acquire_bits_is_builtin_type & T174;
  assign T174 = io_in_acquire_bits_a_type == 3'h3;
  assign T175 = T176;
  assign T176 = {T182, T177};
  assign T177 = 8'h0 - T326;
  assign T326 = {7'h0, T178};
  assign T178 = T179[1'h0:1'h0];
  assign T179 = 1'h1 << T180;
  assign T180 = T181[2'h3:2'h3];
  assign T181 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T182 = 8'h0 - T327;
  assign T327 = {7'h0, T183};
  assign T183 = T179[1'h1:1'h1];
  assign T184 = io_in_acquire_bits_is_builtin_type & T185;
  assign T185 = io_in_acquire_bits_a_type == 3'h4;
  assign T328 = {8'h0, T186};
  assign T186 = R164 >> 4'h8;
  assign io_out_acquire_bits_a_type = T187;
  assign T187 = R83 ? T194 : T188;
  assign T188 = T129 ? T193 : T189;
  assign T189 = T72 ? T192 : T190;
  assign T190 = T17 ? T191 : io_in_acquire_bits_a_type;
  assign T191 = 3'h0;
  assign T192 = 3'h2;
  assign T193 = 3'h1;
  assign T194 = 3'h3;
  assign io_out_acquire_bits_is_builtin_type = T195;
  assign T195 = R83 ? T202 : T196;
  assign T196 = T129 ? T201 : T197;
  assign T197 = T72 ? T200 : T198;
  assign T198 = T17 ? T199 : io_in_acquire_bits_is_builtin_type;
  assign T199 = 1'h1;
  assign T200 = 1'h1;
  assign T201 = 1'h1;
  assign T202 = 1'h1;
  assign io_out_acquire_bits_addr_beat = T203;
  assign T203 = R83 ? T216 : T204;
  assign T204 = T129 ? T215 : T205;
  assign T205 = T72 ? T212 : T206;
  assign T206 = T17 ? T207 : T329;
  assign T329 = {1'h0, io_in_acquire_bits_addr_beat};
  assign T207 = T208;
  assign T208 = T209[3'h5:2'h3];
  assign T209 = {io_in_acquire_bits_addr_block, T210};
  assign T210 = {io_in_acquire_bits_addr_beat, T211};
  assign T211 = io_in_acquire_bits_union[4'hc:4'h9];
  assign T212 = T213;
  assign T213 = {io_in_acquire_bits_addr_beat, T330};
  assign T330 = T331 == 1'h0;
  assign T331 = T26[1'h0:1'h0];
  assign T215 = 3'h0;
  assign T216 = T217;
  assign T217 = {R218, R91};
  assign T219 = T86 ? io_in_acquire_bits_addr_beat : R218;
  assign io_out_acquire_bits_client_xact_id = T220;
  assign T220 = R83 ? T227 : T221;
  assign T221 = T129 ? T226 : T222;
  assign T222 = T72 ? T225 : T223;
  assign T223 = T17 ? T224 : io_in_acquire_bits_client_xact_id;
  assign T224 = io_in_acquire_bits_client_xact_id;
  assign T225 = io_in_acquire_bits_client_xact_id;
  assign T226 = io_in_acquire_bits_client_xact_id;
  assign T227 = R228;
  assign T229 = T86 ? io_in_acquire_bits_client_xact_id : R228;
  assign io_out_acquire_bits_addr_block = T230;
  assign T230 = R83 ? T237 : T231;
  assign T231 = T129 ? T236 : T232;
  assign T232 = T72 ? T235 : T233;
  assign T233 = T17 ? T234 : io_in_acquire_bits_addr_block;
  assign T234 = io_in_acquire_bits_addr_block;
  assign T235 = io_in_acquire_bits_addr_block;
  assign T236 = io_in_acquire_bits_addr_block;
  assign T237 = R238;
  assign T239 = T86 ? io_in_acquire_bits_addr_block : R238;
  assign io_out_acquire_valid = T240;
  assign T240 = T242 | T241;
  assign T241 = T96 & ReorderQueue_io_enq_ready;
  assign T242 = R83 | T243;
  assign T243 = T245 & T244;
  assign T244 = T17 ^ 1'h1;
  assign T245 = io_in_acquire_valid & T246;
  assign T246 = T87 ^ 1'h1;
  assign io_in_grant_bits_data = T247;
  assign T247 = R103 ? T252 : T248;
  assign T248 = T75 ? T249 : T332;
  assign T332 = {64'h0, io_out_grant_bits_data};
  assign T249 = T333;
  assign T333 = T250[7'h7f:1'h0];
  assign T250 = io_out_grant_bits_data << T251;
  assign T251 = {ReorderQueue_io_deq_data, 6'h0};
  assign T252 = T253;
  assign T253 = T254;
  assign T254 = {R261, R255};
  assign T256 = T257 ? io_out_grant_bits_data : R255;
  assign T257 = T111 & T258;
  assign T258 = T259[1'h0:1'h0];
  assign T259 = 1'h1 << T260;
  assign T260 = R108;
  assign T262 = T263 ? io_out_grant_bits_data : R261;
  assign T263 = T111 & T264;
  assign T264 = T259[1'h1:1'h1];
  assign io_in_grant_bits_g_type = T265;
  assign T265 = R103 ? T268 : T266;
  assign T266 = T75 ? T267 : io_out_grant_bits_g_type;
  assign T267 = 4'h4;
  assign T268 = 4'h5;
  assign io_in_grant_bits_is_builtin_type = T269;
  assign T269 = R103 ? T272 : T270;
  assign T270 = T75 ? T271 : io_out_grant_bits_is_builtin_type;
  assign T271 = 1'h1;
  assign T272 = 1'h1;
  assign io_in_grant_bits_manager_xact_id = T273;
  assign T273 = R103 ? T276 : T274;
  assign T274 = T75 ? T275 : io_out_grant_bits_manager_xact_id;
  assign T275 = io_out_grant_bits_manager_xact_id;
  assign T276 = R277;
  assign T278 = T106 ? io_out_grant_bits_manager_xact_id : R277;
  assign io_in_grant_bits_client_xact_id = T279;
  assign T279 = R103 ? T282 : T280;
  assign T280 = T75 ? T281 : io_out_grant_bits_client_xact_id;
  assign T281 = io_out_grant_bits_client_xact_id;
  assign T282 = R283;
  assign T284 = T106 ? io_out_grant_bits_client_xact_id : R283;
  assign io_in_grant_bits_addr_beat = T334;
  assign T334 = T285[1'h1:1'h0];
  assign T285 = R103 ? T336 : T286;
  assign T286 = T75 ? T335 : io_out_grant_bits_addr_beat;
  assign T335 = {1'h0, T287};
  assign T287 = T288;
  assign T288 = io_out_grant_bits_addr_beat >> 1'h1;
  assign T336 = {1'h0, T289};
  assign T289 = R290;
  assign T337 = reset ? 2'h0 : T291;
  assign T291 = T114 ? T292 : R290;
  assign T292 = R290 + 2'h1;
  assign io_in_grant_valid = T293;
  assign T293 = R103 | T294;
  assign T294 = io_out_grant_valid & T295;
  assign T295 = T99 ^ 1'h1;
  assign io_in_acquire_ready = T296;
  assign T296 = T302 & T297;
  assign T297 = T299 | T298;
  assign T298 = ReorderQueue_io_enq_ready & io_out_acquire_ready;
  assign T299 = T87 | T300;
  assign T300 = T301 & io_out_acquire_ready;
  assign T301 = T17 ^ 1'h1;
  assign T302 = R83 ^ 1'h1;
  ReorderQueue_0 ReorderQueue(.clk(clk), .reset(reset),
       .io_enq_ready( ReorderQueue_io_enq_ready ),
       .io_enq_valid( T81 ),
       .io_enq_bits_data( T77 ),
       .io_enq_bits_tag( io_in_acquire_bits_client_xact_id ),
       .io_deq_valid( T74 ),
       .io_deq_tag( io_out_grant_bits_client_xact_id ),
       .io_deq_data( ReorderQueue_io_deq_data )
       //.io_deq_matches(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T19 <= 1'b1;
  if(!T20 && T19 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Put wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't perform Get wider than outer width");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R83 <= 1'h0;
    end else if(T89) begin
      R83 <= 1'h0;
    end else if(T86) begin
      R83 <= 1'h1;
    end
    if(reset) begin
      R91 <= 1'h0;
    end else if(T94) begin
      R91 <= T93;
    end
    if(reset) begin
      R103 <= 1'h0;
    end else if(T114) begin
      R103 <= 1'h0;
    end else if(T106) begin
      R103 <= 1'h1;
    end
    if(reset) begin
      R108 <= 1'h0;
    end else if(T111) begin
      R108 <= T110;
    end
    if(T94) begin
      R132 <= T317;
    end else if(T86) begin
      R132 <= io_in_acquire_bits_data;
    end
    if(T94) begin
      R164 <= T328;
    end else if(T86) begin
      R164 <= T167;
    end
    if(T86) begin
      R218 <= io_in_acquire_bits_addr_beat;
    end
    if(T86) begin
      R228 <= io_in_acquire_bits_client_xact_id;
    end
    if(T86) begin
      R238 <= io_in_acquire_bits_addr_block;
    end
    if(T257) begin
      R255 <= io_out_grant_bits_data;
    end
    if(T263) begin
      R261 <= io_out_grant_bits_data;
    end
    if(T106) begin
      R277 <= io_out_grant_bits_manager_xact_id;
    end
    if(T106) begin
      R283 <= io_out_grant_bits_client_xact_id;
    end
    if(reset) begin
      R290 <= 2'h0;
    end else if(T114) begin
      R290 <= T292;
    end
  end
endmodule

module ReorderQueue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [2:0] io_enq_bits_data_addr_beat,
    input [2:0] io_enq_bits_data_byteOff,
    input  io_enq_bits_data_subblock,
    input [3:0] io_enq_bits_tag,
    input  io_deq_valid,
    input [3:0] io_deq_tag,
    output[2:0] io_deq_data_addr_beat,
    output[2:0] io_deq_data_byteOff,
    output io_deq_data_subblock,
    output io_deq_matches
);

  wire T0;
  wire roq_matches_5;
  wire T1;
  reg  roq_free_5;
  wire T166;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire[7:0] T6;
  wire[2:0] T7;
  wire[2:0] roq_enq_addr;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  reg  roq_free_4;
  wire T167;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[7:0] T18;
  wire[2:0] T19;
  wire[2:0] roq_deq_addr;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire roq_matches_4;
  wire T24;
  wire T25;
  reg [3:0] roq_tags_4;
  wire[3:0] T26;
  wire T27;
  wire T28;
  wire[7:0] T29;
  wire[2:0] T30;
  wire roq_matches_3;
  wire T31;
  wire T32;
  reg [3:0] roq_tags_3;
  wire[3:0] T33;
  wire T34;
  wire T35;
  wire roq_matches_2;
  wire T36;
  wire T37;
  reg [3:0] roq_tags_2;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire roq_matches_1;
  wire T41;
  wire T42;
  reg [3:0] roq_tags_1;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire roq_matches_0;
  wire T46;
  wire T47;
  reg [3:0] roq_tags_0;
  wire[3:0] T48;
  wire T49;
  wire T50;
  reg  roq_free_3;
  wire T168;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  reg  roq_free_2;
  wire T169;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  roq_free_1;
  wire T170;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  reg  roq_free_0;
  wire T171;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [3:0] roq_tags_5;
  wire[3:0] T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  reg  roq_data_0_subblock;
  wire T89;
  wire T90;
  wire T91;
  wire[7:0] T92;
  wire[2:0] T93;
  reg  roq_data_1_subblock;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire[2:0] T98;
  wire T99;
  reg  roq_data_2_subblock;
  wire T100;
  wire T101;
  wire T102;
  reg  roq_data_3_subblock;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  reg  roq_data_4_subblock;
  wire T109;
  wire T110;
  wire T111;
  reg  roq_data_5_subblock;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire[2:0] T119;
  reg [2:0] roq_data_0_byteOff;
  wire[2:0] T120;
  wire T121;
  reg [2:0] roq_data_1_byteOff;
  wire[2:0] T122;
  wire T123;
  wire T124;
  wire[2:0] T125;
  reg [2:0] roq_data_2_byteOff;
  wire[2:0] T126;
  wire T127;
  reg [2:0] roq_data_3_byteOff;
  wire[2:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  reg [2:0] roq_data_4_byteOff;
  wire[2:0] T133;
  wire T134;
  reg [2:0] roq_data_5_byteOff;
  wire[2:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire[2:0] T139;
  wire[2:0] T140;
  wire[2:0] T141;
  reg [2:0] roq_data_0_addr_beat;
  wire[2:0] T142;
  wire T143;
  reg [2:0] roq_data_1_addr_beat;
  wire[2:0] T144;
  wire T145;
  wire T146;
  wire[2:0] T147;
  reg [2:0] roq_data_2_addr_beat;
  wire[2:0] T148;
  wire T149;
  reg [2:0] roq_data_3_addr_beat;
  wire[2:0] T150;
  wire T151;
  wire T152;
  wire T153;
  wire[2:0] T154;
  reg [2:0] roq_data_4_addr_beat;
  wire[2:0] T155;
  wire T156;
  reg [2:0] roq_data_5_addr_beat;
  wire[2:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    roq_free_5 = {1{$random}};
    roq_free_4 = {1{$random}};
    roq_tags_4 = {1{$random}};
    roq_tags_3 = {1{$random}};
    roq_tags_2 = {1{$random}};
    roq_tags_1 = {1{$random}};
    roq_tags_0 = {1{$random}};
    roq_free_3 = {1{$random}};
    roq_free_2 = {1{$random}};
    roq_free_1 = {1{$random}};
    roq_free_0 = {1{$random}};
    roq_tags_5 = {1{$random}};
    roq_data_0_subblock = {1{$random}};
    roq_data_1_subblock = {1{$random}};
    roq_data_2_subblock = {1{$random}};
    roq_data_3_subblock = {1{$random}};
    roq_data_4_subblock = {1{$random}};
    roq_data_5_subblock = {1{$random}};
    roq_data_0_byteOff = {1{$random}};
    roq_data_1_byteOff = {1{$random}};
    roq_data_2_byteOff = {1{$random}};
    roq_data_3_byteOff = {1{$random}};
    roq_data_4_byteOff = {1{$random}};
    roq_data_5_byteOff = {1{$random}};
    roq_data_0_addr_beat = {1{$random}};
    roq_data_1_addr_beat = {1{$random}};
    roq_data_2_addr_beat = {1{$random}};
    roq_data_3_addr_beat = {1{$random}};
    roq_data_4_addr_beat = {1{$random}};
    roq_data_5_addr_beat = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_deq_matches = T0;
  assign T0 = T82 | roq_matches_5;
  assign roq_matches_5 = T78 & T1;
  assign T1 = roq_free_5 ^ 1'h1;
  assign T166 = reset ? 1'h1 : T2;
  assign T2 = T76 ? 1'h1 : T3;
  assign T3 = T4 ? 1'h0 : roq_free_5;
  assign T4 = T75 & T5;
  assign T5 = T6[3'h5:3'h5];
  assign T6 = 1'h1 << T7;
  assign T7 = roq_enq_addr;
  assign roq_enq_addr = roq_free_0 ? 3'h0 : T8;
  assign T8 = roq_free_1 ? 3'h1 : T9;
  assign T9 = roq_free_2 ? 3'h2 : T10;
  assign T10 = roq_free_3 ? 3'h3 : T11;
  assign T11 = roq_free_4 ? 3'h4 : 3'h5;
  assign T167 = reset ? 1'h1 : T12;
  assign T12 = T16 ? 1'h1 : T13;
  assign T13 = T14 ? 1'h0 : roq_free_4;
  assign T14 = T75 & T15;
  assign T15 = T6[3'h4:3'h4];
  assign T16 = io_deq_valid & T17;
  assign T17 = T18[3'h4:3'h4];
  assign T18 = 1'h1 << T19;
  assign T19 = roq_deq_addr;
  assign roq_deq_addr = roq_matches_0 ? 3'h0 : T20;
  assign T20 = roq_matches_1 ? 3'h1 : T21;
  assign T21 = roq_matches_2 ? 3'h2 : T22;
  assign T22 = roq_matches_3 ? 3'h3 : T23;
  assign T23 = roq_matches_4 ? 3'h4 : 3'h5;
  assign roq_matches_4 = T25 & T24;
  assign T24 = roq_free_4 ^ 1'h1;
  assign T25 = roq_tags_4 == io_deq_tag;
  assign T26 = T27 ? io_enq_bits_tag : roq_tags_4;
  assign T27 = T75 & T28;
  assign T28 = T29[3'h4:3'h4];
  assign T29 = 1'h1 << T30;
  assign T30 = roq_enq_addr;
  assign roq_matches_3 = T32 & T31;
  assign T31 = roq_free_3 ^ 1'h1;
  assign T32 = roq_tags_3 == io_deq_tag;
  assign T33 = T34 ? io_enq_bits_tag : roq_tags_3;
  assign T34 = T75 & T35;
  assign T35 = T29[2'h3:2'h3];
  assign roq_matches_2 = T37 & T36;
  assign T36 = roq_free_2 ^ 1'h1;
  assign T37 = roq_tags_2 == io_deq_tag;
  assign T38 = T39 ? io_enq_bits_tag : roq_tags_2;
  assign T39 = T75 & T40;
  assign T40 = T29[2'h2:2'h2];
  assign roq_matches_1 = T42 & T41;
  assign T41 = roq_free_1 ^ 1'h1;
  assign T42 = roq_tags_1 == io_deq_tag;
  assign T43 = T44 ? io_enq_bits_tag : roq_tags_1;
  assign T44 = T75 & T45;
  assign T45 = T29[1'h1:1'h1];
  assign roq_matches_0 = T47 & T46;
  assign T46 = roq_free_0 ^ 1'h1;
  assign T47 = roq_tags_0 == io_deq_tag;
  assign T48 = T49 ? io_enq_bits_tag : roq_tags_0;
  assign T49 = T75 & T50;
  assign T50 = T29[1'h0:1'h0];
  assign T168 = reset ? 1'h1 : T51;
  assign T51 = T55 ? 1'h1 : T52;
  assign T52 = T53 ? 1'h0 : roq_free_3;
  assign T53 = T75 & T54;
  assign T54 = T6[2'h3:2'h3];
  assign T55 = io_deq_valid & T56;
  assign T56 = T18[2'h3:2'h3];
  assign T169 = reset ? 1'h1 : T57;
  assign T57 = T61 ? 1'h1 : T58;
  assign T58 = T59 ? 1'h0 : roq_free_2;
  assign T59 = T75 & T60;
  assign T60 = T6[2'h2:2'h2];
  assign T61 = io_deq_valid & T62;
  assign T62 = T18[2'h2:2'h2];
  assign T170 = reset ? 1'h1 : T63;
  assign T63 = T67 ? 1'h1 : T64;
  assign T64 = T65 ? 1'h0 : roq_free_1;
  assign T65 = T75 & T66;
  assign T66 = T6[1'h1:1'h1];
  assign T67 = io_deq_valid & T68;
  assign T68 = T18[1'h1:1'h1];
  assign T171 = reset ? 1'h1 : T69;
  assign T69 = T73 ? 1'h1 : T70;
  assign T70 = T71 ? 1'h0 : roq_free_0;
  assign T71 = T75 & T72;
  assign T72 = T6[1'h0:1'h0];
  assign T73 = io_deq_valid & T74;
  assign T74 = T18[1'h0:1'h0];
  assign T75 = io_enq_valid & io_enq_ready;
  assign T76 = io_deq_valid & T77;
  assign T77 = T18[3'h5:3'h5];
  assign T78 = roq_tags_5 == io_deq_tag;
  assign T79 = T80 ? io_enq_bits_tag : roq_tags_5;
  assign T80 = T75 & T81;
  assign T81 = T29[3'h5:3'h5];
  assign T82 = T83 | roq_matches_4;
  assign T83 = T84 | roq_matches_3;
  assign T84 = T85 | roq_matches_2;
  assign T85 = roq_matches_0 | roq_matches_1;
  assign io_deq_data_subblock = T86;
  assign T86 = T116 ? T108 : T87;
  assign T87 = T107 ? T99 : T88;
  assign T88 = T97 ? roq_data_1_subblock : roq_data_0_subblock;
  assign T89 = T90 ? io_enq_bits_data_subblock : roq_data_0_subblock;
  assign T90 = T75 & T91;
  assign T91 = T92[1'h0:1'h0];
  assign T92 = 1'h1 << T93;
  assign T93 = roq_enq_addr;
  assign T94 = T95 ? io_enq_bits_data_subblock : roq_data_1_subblock;
  assign T95 = T75 & T96;
  assign T96 = T92[1'h1:1'h1];
  assign T97 = T98[1'h0:1'h0];
  assign T98 = roq_deq_addr;
  assign T99 = T106 ? roq_data_3_subblock : roq_data_2_subblock;
  assign T100 = T101 ? io_enq_bits_data_subblock : roq_data_2_subblock;
  assign T101 = T75 & T102;
  assign T102 = T92[2'h2:2'h2];
  assign T103 = T104 ? io_enq_bits_data_subblock : roq_data_3_subblock;
  assign T104 = T75 & T105;
  assign T105 = T92[2'h3:2'h3];
  assign T106 = T98[1'h0:1'h0];
  assign T107 = T98[1'h1:1'h1];
  assign T108 = T115 ? roq_data_5_subblock : roq_data_4_subblock;
  assign T109 = T110 ? io_enq_bits_data_subblock : roq_data_4_subblock;
  assign T110 = T75 & T111;
  assign T111 = T92[3'h4:3'h4];
  assign T112 = T113 ? io_enq_bits_data_subblock : roq_data_5_subblock;
  assign T113 = T75 & T114;
  assign T114 = T92[3'h5:3'h5];
  assign T115 = T98[1'h0:1'h0];
  assign T116 = T98[2'h2:2'h2];
  assign io_deq_data_byteOff = T117;
  assign T117 = T138 ? T132 : T118;
  assign T118 = T131 ? T125 : T119;
  assign T119 = T124 ? roq_data_1_byteOff : roq_data_0_byteOff;
  assign T120 = T121 ? io_enq_bits_data_byteOff : roq_data_0_byteOff;
  assign T121 = T75 & T91;
  assign T122 = T123 ? io_enq_bits_data_byteOff : roq_data_1_byteOff;
  assign T123 = T75 & T96;
  assign T124 = T98[1'h0:1'h0];
  assign T125 = T130 ? roq_data_3_byteOff : roq_data_2_byteOff;
  assign T126 = T127 ? io_enq_bits_data_byteOff : roq_data_2_byteOff;
  assign T127 = T75 & T102;
  assign T128 = T129 ? io_enq_bits_data_byteOff : roq_data_3_byteOff;
  assign T129 = T75 & T105;
  assign T130 = T98[1'h0:1'h0];
  assign T131 = T98[1'h1:1'h1];
  assign T132 = T137 ? roq_data_5_byteOff : roq_data_4_byteOff;
  assign T133 = T134 ? io_enq_bits_data_byteOff : roq_data_4_byteOff;
  assign T134 = T75 & T111;
  assign T135 = T136 ? io_enq_bits_data_byteOff : roq_data_5_byteOff;
  assign T136 = T75 & T114;
  assign T137 = T98[1'h0:1'h0];
  assign T138 = T98[2'h2:2'h2];
  assign io_deq_data_addr_beat = T139;
  assign T139 = T160 ? T154 : T140;
  assign T140 = T153 ? T147 : T141;
  assign T141 = T146 ? roq_data_1_addr_beat : roq_data_0_addr_beat;
  assign T142 = T143 ? io_enq_bits_data_addr_beat : roq_data_0_addr_beat;
  assign T143 = T75 & T91;
  assign T144 = T145 ? io_enq_bits_data_addr_beat : roq_data_1_addr_beat;
  assign T145 = T75 & T96;
  assign T146 = T98[1'h0:1'h0];
  assign T147 = T152 ? roq_data_3_addr_beat : roq_data_2_addr_beat;
  assign T148 = T149 ? io_enq_bits_data_addr_beat : roq_data_2_addr_beat;
  assign T149 = T75 & T102;
  assign T150 = T151 ? io_enq_bits_data_addr_beat : roq_data_3_addr_beat;
  assign T151 = T75 & T105;
  assign T152 = T98[1'h0:1'h0];
  assign T153 = T98[1'h1:1'h1];
  assign T154 = T159 ? roq_data_5_addr_beat : roq_data_4_addr_beat;
  assign T155 = T156 ? io_enq_bits_data_addr_beat : roq_data_4_addr_beat;
  assign T156 = T75 & T111;
  assign T157 = T158 ? io_enq_bits_data_addr_beat : roq_data_5_addr_beat;
  assign T158 = T75 & T114;
  assign T159 = T98[1'h0:1'h0];
  assign T160 = T98[2'h2:2'h2];
  assign io_enq_ready = T161;
  assign T161 = T162 | roq_free_5;
  assign T162 = T163 | roq_free_4;
  assign T163 = T164 | roq_free_3;
  assign T164 = T165 | roq_free_2;
  assign T165 = roq_free_0 | roq_free_1;

  always @(posedge clk) begin
    if(reset) begin
      roq_free_5 <= 1'h1;
    end else if(T76) begin
      roq_free_5 <= 1'h1;
    end else if(T4) begin
      roq_free_5 <= 1'h0;
    end
    if(reset) begin
      roq_free_4 <= 1'h1;
    end else if(T16) begin
      roq_free_4 <= 1'h1;
    end else if(T14) begin
      roq_free_4 <= 1'h0;
    end
    if(T27) begin
      roq_tags_4 <= io_enq_bits_tag;
    end
    if(T34) begin
      roq_tags_3 <= io_enq_bits_tag;
    end
    if(T39) begin
      roq_tags_2 <= io_enq_bits_tag;
    end
    if(T44) begin
      roq_tags_1 <= io_enq_bits_tag;
    end
    if(T49) begin
      roq_tags_0 <= io_enq_bits_tag;
    end
    if(reset) begin
      roq_free_3 <= 1'h1;
    end else if(T55) begin
      roq_free_3 <= 1'h1;
    end else if(T53) begin
      roq_free_3 <= 1'h0;
    end
    if(reset) begin
      roq_free_2 <= 1'h1;
    end else if(T61) begin
      roq_free_2 <= 1'h1;
    end else if(T59) begin
      roq_free_2 <= 1'h0;
    end
    if(reset) begin
      roq_free_1 <= 1'h1;
    end else if(T67) begin
      roq_free_1 <= 1'h1;
    end else if(T65) begin
      roq_free_1 <= 1'h0;
    end
    if(reset) begin
      roq_free_0 <= 1'h1;
    end else if(T73) begin
      roq_free_0 <= 1'h1;
    end else if(T71) begin
      roq_free_0 <= 1'h0;
    end
    if(T80) begin
      roq_tags_5 <= io_enq_bits_tag;
    end
    if(T90) begin
      roq_data_0_subblock <= io_enq_bits_data_subblock;
    end
    if(T95) begin
      roq_data_1_subblock <= io_enq_bits_data_subblock;
    end
    if(T101) begin
      roq_data_2_subblock <= io_enq_bits_data_subblock;
    end
    if(T104) begin
      roq_data_3_subblock <= io_enq_bits_data_subblock;
    end
    if(T110) begin
      roq_data_4_subblock <= io_enq_bits_data_subblock;
    end
    if(T113) begin
      roq_data_5_subblock <= io_enq_bits_data_subblock;
    end
    if(T121) begin
      roq_data_0_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T123) begin
      roq_data_1_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T127) begin
      roq_data_2_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T129) begin
      roq_data_3_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T134) begin
      roq_data_4_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T136) begin
      roq_data_5_byteOff <= io_enq_bits_data_byteOff;
    end
    if(T143) begin
      roq_data_0_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T145) begin
      roq_data_1_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T149) begin
      roq_data_2_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T151) begin
      roq_data_3_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T156) begin
      roq_data_4_addr_beat <= io_enq_bits_data_addr_beat;
    end
    if(T158) begin
      roq_data_5_addr_beat <= io_enq_bits_data_addr_beat;
    end
  end
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [2:0] io_in_1_bits_addr_beat,
    input [2:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_manager_xact_id,
    input  io_in_1_bits_is_builtin_type,
    input [3:0] io_in_1_bits_g_type,
    input [63:0] io_in_1_bits_data,
    input  io_in_1_bits_client_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [2:0] io_in_0_bits_addr_beat,
    input [2:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_manager_xact_id,
    input  io_in_0_bits_is_builtin_type,
    input [3:0] io_in_0_bits_g_type,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_client_id,
    input  io_out_ready,
    output io_out_valid,
    output[2:0] io_out_bits_addr_beat,
    output[2:0] io_out_bits_client_xact_id,
    output io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[63:0] io_out_bits_data,
    output io_out_bits_client_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[3:0] T3;
  wire T4;
  wire T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_client_id = T0;
  assign T0 = T1 ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_g_type = T3;
  assign T3 = T1 ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign io_out_bits_is_builtin_type = T4;
  assign T4 = T1 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module NastiIOTileLinkIOConverter(input clk, input reset,
    output io_tl_acquire_ready,
    input  io_tl_acquire_valid,
    input [25:0] io_tl_acquire_bits_addr_block,
    input [2:0] io_tl_acquire_bits_client_xact_id,
    input [2:0] io_tl_acquire_bits_addr_beat,
    input  io_tl_acquire_bits_is_builtin_type,
    input [2:0] io_tl_acquire_bits_a_type,
    input [11:0] io_tl_acquire_bits_union,
    input [63:0] io_tl_acquire_bits_data,
    input  io_tl_grant_ready,
    output io_tl_grant_valid,
    output[2:0] io_tl_grant_bits_addr_beat,
    output[2:0] io_tl_grant_bits_client_xact_id,
    output io_tl_grant_bits_manager_xact_id,
    output io_tl_grant_bits_is_builtin_type,
    output[3:0] io_tl_grant_bits_g_type,
    output[63:0] io_tl_grant_bits_data,
    input  io_nasti_aw_ready,
    output io_nasti_aw_valid,
    output[31:0] io_nasti_aw_bits_addr,
    output[7:0] io_nasti_aw_bits_len,
    output[2:0] io_nasti_aw_bits_size,
    output[1:0] io_nasti_aw_bits_burst,
    output io_nasti_aw_bits_lock,
    output[3:0] io_nasti_aw_bits_cache,
    output[2:0] io_nasti_aw_bits_prot,
    output[3:0] io_nasti_aw_bits_qos,
    output[3:0] io_nasti_aw_bits_region,
    output[3:0] io_nasti_aw_bits_id,
    output io_nasti_aw_bits_user,
    input  io_nasti_w_ready,
    output io_nasti_w_valid,
    output[63:0] io_nasti_w_bits_data,
    output io_nasti_w_bits_last,
    output[7:0] io_nasti_w_bits_strb,
    output io_nasti_w_bits_user,
    output io_nasti_b_ready,
    input  io_nasti_b_valid,
    input [1:0] io_nasti_b_bits_resp,
    input [3:0] io_nasti_b_bits_id,
    input  io_nasti_b_bits_user,
    input  io_nasti_ar_ready,
    output io_nasti_ar_valid,
    output[31:0] io_nasti_ar_bits_addr,
    output[7:0] io_nasti_ar_bits_len,
    output[2:0] io_nasti_ar_bits_size,
    output[1:0] io_nasti_ar_bits_burst,
    output io_nasti_ar_bits_lock,
    output[3:0] io_nasti_ar_bits_cache,
    output[2:0] io_nasti_ar_bits_prot,
    output[3:0] io_nasti_ar_bits_qos,
    output[3:0] io_nasti_ar_bits_region,
    output[3:0] io_nasti_ar_bits_id,
    output io_nasti_ar_bits_user,
    output io_nasti_r_ready,
    input  io_nasti_r_valid,
    input [1:0] io_nasti_r_bits_resp,
    input [63:0] io_nasti_r_bits_data,
    input  io_nasti_r_bits_last,
    input [3:0] io_nasti_r_bits_id,
    input  io_nasti_r_bits_user
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg[0:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[63:0] T145;
  wire[126:0] r_aligned_data;
  wire[126:0] T146;
  wire[126:0] T11;
  wire[5:0] T12;
  wire[3:0] T13;
  wire[3:0] T147;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[2:0] T148;
  wire[2:0] T18;
  wire[2:0] T19;
  reg [2:0] tl_cnt_in;
  wire[2:0] T149;
  wire[2:0] T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[63:0] T27;
  wire[3:0] T28;
  wire T29;
  wire T30;
  wire[2:0] T31;
  wire[2:0] T150;
  wire[2:0] T32;
  wire T33;
  wire T34;
  wire nasti_wrap_out;
  wire T35;
  reg [2:0] nasti_cnt_out;
  wire[2:0] T151;
  wire[2:0] T36;
  wire[2:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire is_subblock;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[2:0] T47;
  wire T48;
  wire get_valid;
  wire T49;
  wire has_data;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T152;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[2:0] T59;
  wire[3:0] T60;
  wire T61;
  wire[1:0] T62;
  wire[2:0] T63;
  wire[2:0] T64;
  wire[2:0] T65;
  wire[2:0] T66;
  wire[2:0] T67;
  wire[2:0] T68;
  wire[2:0] T69;
  wire[2:0] T70;
  wire[2:0] T71;
  wire T72;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[7:0] T80;
  wire[7:0] T153;
  wire[2:0] T81;
  wire[31:0] T82;
  wire[31:0] T83;
  wire[5:0] T84;
  wire[2:0] T85;
  wire T86;
  wire T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T154;
  wire T99;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire tl_wrap_out;
  wire T109;
  reg [2:0] tl_cnt_out;
  wire[2:0] T155;
  wire[2:0] T110;
  wire[2:0] T111;
  wire T112;
  wire is_multibeat;
  wire T113;
  wire T114;
  wire[63:0] T115;
  wire T116;
  wire aw_ready;
  reg  w_inflight;
  wire T156;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire put_valid;
  wire T124;
  wire[3:0] T125;
  wire[3:0] T157;
  wire[3:0] T126;
  wire[3:0] T127;
  wire[2:0] T128;
  wire[3:0] T129;
  wire T130;
  wire[1:0] T131;
  wire[2:0] T132;
  wire[7:0] T133;
  wire[7:0] T158;
  wire[2:0] T134;
  wire[31:0] T135;
  wire[31:0] T136;
  wire[5:0] T137;
  wire[2:0] T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire roq_io_enq_ready;
  wire[2:0] roq_io_deq_data_addr_beat;
  wire[2:0] roq_io_deq_data_byteOff;
  wire roq_io_deq_data_subblock;
  wire gnt_arb_io_in_1_ready;
  wire gnt_arb_io_in_0_ready;
  wire gnt_arb_io_out_valid;
  wire[2:0] gnt_arb_io_out_bits_addr_beat;
  wire[2:0] gnt_arb_io_out_bits_client_xact_id;
  wire gnt_arb_io_out_bits_manager_xact_id;
  wire gnt_arb_io_out_bits_is_builtin_type;
  wire[3:0] gnt_arb_io_out_bits_g_type;
  wire[63:0] gnt_arb_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T5 = 1'b0;
    tl_cnt_in = {1{$random}};
    nasti_cnt_out = {1{$random}};
    tl_cnt_out = {1{$random}};
    w_inflight = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = io_nasti_b_bits_resp == 2'h0;
  assign T4 = io_nasti_b_valid ^ 1'h1;
  assign T6 = T7 | reset;
  assign T7 = T9 | T8;
  assign T8 = io_nasti_r_bits_resp == 2'h0;
  assign T9 = io_nasti_r_valid ^ 1'h1;
  assign T10 = T145;
  assign T145 = r_aligned_data[6'h3f:1'h0];
  assign r_aligned_data = roq_io_deq_data_subblock ? T11 : T146;
  assign T146 = {63'h0, io_nasti_r_bits_data};
  assign T11 = io_nasti_r_bits_data << T12;
  assign T12 = {roq_io_deq_data_byteOff, 3'h0};
  assign T13 = T147;
  assign T147 = {1'h0, T14};
  assign T14 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T15 = 1'h1;
  assign T16 = 1'h0;
  assign T17 = T148;
  assign T148 = io_nasti_r_bits_id[2'h2:1'h0];
  assign T18 = T19;
  assign T19 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T149 = reset ? 3'h0 : T20;
  assign T20 = T22 ? T21 : tl_cnt_in;
  assign T21 = tl_cnt_in + 3'h1;
  assign T22 = T26 & T23;
  assign T23 = io_tl_grant_bits_is_builtin_type ? T25 : T24;
  assign T24 = 4'h0 == io_tl_grant_bits_g_type;
  assign T25 = 4'h5 == io_tl_grant_bits_g_type;
  assign T26 = io_tl_grant_ready & io_tl_grant_valid;
  assign T27 = 64'h0;
  assign T28 = 4'h3;
  assign T29 = 1'h1;
  assign T30 = 1'h0;
  assign T31 = T150;
  assign T150 = io_nasti_b_bits_id[2'h2:1'h0];
  assign T32 = 3'h0;
  assign T33 = T41 & T34;
  assign T34 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign nasti_wrap_out = T38 & T35;
  assign T35 = nasti_cnt_out == 3'h7;
  assign T151 = reset ? 3'h0 : T36;
  assign T36 = T38 ? T37 : nasti_cnt_out;
  assign T37 = nasti_cnt_out + 3'h1;
  assign T38 = T40 & T39;
  assign T39 = roq_io_deq_data_subblock ^ 1'h1;
  assign T40 = io_nasti_r_ready & io_nasti_r_valid;
  assign T41 = io_nasti_r_ready & io_nasti_r_valid;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T42;
  assign T42 = T44 | T43;
  assign T43 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T44 = T46 | T45;
  assign T45 = 3'h0 == io_tl_acquire_bits_a_type;
  assign T46 = 3'h2 == io_tl_acquire_bits_a_type;
  assign T47 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign T48 = get_valid & io_nasti_ar_ready;
  assign get_valid = io_tl_acquire_valid & T49;
  assign T49 = has_data ^ 1'h1;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T50;
  assign T50 = T52 | T51;
  assign T51 = 3'h4 == io_tl_acquire_bits_a_type;
  assign T52 = T54 | T53;
  assign T53 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T54 = 3'h2 == io_tl_acquire_bits_a_type;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign io_nasti_ar_bits_user = T55;
  assign T55 = 1'h0;
  assign io_nasti_ar_bits_id = T56;
  assign T56 = T152;
  assign T152 = {1'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_ar_bits_region = T57;
  assign T57 = 4'h0;
  assign io_nasti_ar_bits_qos = T58;
  assign T58 = 4'h0;
  assign io_nasti_ar_bits_prot = T59;
  assign T59 = 3'h0;
  assign io_nasti_ar_bits_cache = T60;
  assign T60 = 4'h0;
  assign io_nasti_ar_bits_lock = T61;
  assign T61 = 1'h0;
  assign io_nasti_ar_bits_burst = T62;
  assign T62 = 2'h1;
  assign io_nasti_ar_bits_size = T63;
  assign T63 = T64;
  assign T64 = is_subblock ? T65 : 3'h3;
  assign T65 = T79 ? 3'h0 : T66;
  assign T66 = T78 ? 3'h0 : T67;
  assign T67 = T77 ? 3'h1 : T68;
  assign T68 = T76 ? 3'h1 : T69;
  assign T69 = T75 ? 3'h2 : T70;
  assign T70 = T74 ? 3'h3 : T71;
  assign T71 = T72 ? 3'h3 : 3'h7;
  assign T72 = T73 == 3'h7;
  assign T73 = io_tl_acquire_bits_union[4'h8:3'h6];
  assign T74 = T73 == 3'h3;
  assign T75 = T73 == 3'h2;
  assign T76 = T73 == 3'h5;
  assign T77 = T73 == 3'h1;
  assign T78 = T73 == 3'h4;
  assign T79 = T73 == 3'h0;
  assign io_nasti_ar_bits_len = T80;
  assign T80 = T153;
  assign T153 = {5'h0, T81};
  assign T81 = is_subblock ? 3'h0 : 3'h7;
  assign io_nasti_ar_bits_addr = T82;
  assign T82 = T83;
  assign T83 = {io_tl_acquire_bits_addr_block, T84};
  assign T84 = {io_tl_acquire_bits_addr_beat, T85};
  assign T85 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_ar_valid = T86;
  assign T86 = get_valid & roq_io_enq_ready;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_w_bits_user = T87;
  assign T87 = 1'h0;
  assign io_nasti_w_bits_strb = T88;
  assign T88 = T89;
  assign T89 = T103 ? T97 : T90;
  assign T90 = T92 ? T91 : 8'h0;
  assign T91 = io_tl_acquire_bits_union[4'h8:1'h1];
  assign T92 = T95 | T93;
  assign T93 = io_tl_acquire_bits_is_builtin_type & T94;
  assign T94 = io_tl_acquire_bits_a_type == 3'h2;
  assign T95 = io_tl_acquire_bits_is_builtin_type & T96;
  assign T96 = io_tl_acquire_bits_a_type == 3'h3;
  assign T97 = T98;
  assign T98 = 8'h0 - T154;
  assign T154 = {7'h0, T99};
  assign T99 = 1'h1;
  assign T103 = io_tl_acquire_bits_is_builtin_type & T104;
  assign T104 = io_tl_acquire_bits_a_type == 3'h4;
  assign io_nasti_w_bits_last = T105;
  assign T105 = T106;
  assign T106 = tl_wrap_out | T107;
  assign T107 = T108 & is_subblock;
  assign T108 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign tl_wrap_out = T112 & T109;
  assign T109 = tl_cnt_out == 3'h7;
  assign T155 = reset ? 3'h0 : T110;
  assign T110 = T112 ? T111 : tl_cnt_out;
  assign T111 = tl_cnt_out + 3'h1;
  assign T112 = T114 & is_multibeat;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T113;
  assign T113 = 3'h3 == io_tl_acquire_bits_a_type;
  assign T114 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign io_nasti_w_bits_data = T115;
  assign T115 = io_tl_acquire_bits_data;
  assign io_nasti_w_valid = T116;
  assign T116 = put_valid & aw_ready;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T156 = reset ? 1'h0 : T117;
  assign T117 = T123 ? 1'h0 : T118;
  assign T118 = T119 ? 1'h1 : w_inflight;
  assign T119 = T120 & is_multibeat;
  assign T120 = T122 & T121;
  assign T121 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T122 = w_inflight ^ 1'h1;
  assign T123 = w_inflight & tl_wrap_out;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign io_nasti_aw_bits_user = T124;
  assign T124 = 1'h0;
  assign io_nasti_aw_bits_id = T125;
  assign T125 = T157;
  assign T157 = {1'h0, io_tl_acquire_bits_client_xact_id};
  assign io_nasti_aw_bits_region = T126;
  assign T126 = 4'h0;
  assign io_nasti_aw_bits_qos = T127;
  assign T127 = 4'h0;
  assign io_nasti_aw_bits_prot = T128;
  assign T128 = 3'h0;
  assign io_nasti_aw_bits_cache = T129;
  assign T129 = 4'h0;
  assign io_nasti_aw_bits_lock = T130;
  assign T130 = 1'h0;
  assign io_nasti_aw_bits_burst = T131;
  assign T131 = 2'h1;
  assign io_nasti_aw_bits_size = T132;
  assign T132 = 3'h3;
  assign io_nasti_aw_bits_len = T133;
  assign T133 = T158;
  assign T158 = {5'h0, T134};
  assign T134 = is_multibeat ? 3'h7 : 3'h0;
  assign io_nasti_aw_bits_addr = T135;
  assign T135 = T136;
  assign T136 = {io_tl_acquire_bits_addr_block, T137};
  assign T137 = {io_tl_acquire_bits_addr_beat, T138};
  assign T138 = io_tl_acquire_bits_union[4'hb:4'h9];
  assign io_nasti_aw_valid = T139;
  assign T139 = T141 & T140;
  assign T140 = w_inflight ^ 1'h1;
  assign T141 = put_valid & io_nasti_w_ready;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_acquire_ready = T142;
  assign T142 = has_data ? T144 : T143;
  assign T143 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T144 = aw_ready & io_nasti_w_ready;
  ReorderQueue_1 roq(.clk(clk), .reset(reset),
       .io_enq_ready( roq_io_enq_ready ),
       .io_enq_valid( T48 ),
       .io_enq_bits_data_addr_beat( io_tl_acquire_bits_addr_beat ),
       .io_enq_bits_data_byteOff( T47 ),
       .io_enq_bits_data_subblock( is_subblock ),
       .io_enq_bits_tag( io_nasti_ar_bits_id ),
       .io_deq_valid( T33 ),
       .io_deq_tag( io_nasti_r_bits_id ),
       .io_deq_data_addr_beat( roq_io_deq_data_addr_beat ),
       .io_deq_data_byteOff( roq_io_deq_data_byteOff ),
       .io_deq_data_subblock( roq_io_deq_data_subblock )
       //.io_deq_matches(  )
  );
  Arbiter_5 gnt_arb(
       .io_in_1_ready( gnt_arb_io_in_1_ready ),
       .io_in_1_valid( io_nasti_b_valid ),
       .io_in_1_bits_addr_beat( T32 ),
       .io_in_1_bits_client_xact_id( T31 ),
       .io_in_1_bits_manager_xact_id( T30 ),
       .io_in_1_bits_is_builtin_type( T29 ),
       .io_in_1_bits_g_type( T28 ),
       .io_in_1_bits_data( T27 ),
       //.io_in_1_bits_client_id(  )
       .io_in_0_ready( gnt_arb_io_in_0_ready ),
       .io_in_0_valid( io_nasti_r_valid ),
       .io_in_0_bits_addr_beat( T18 ),
       .io_in_0_bits_client_xact_id( T17 ),
       .io_in_0_bits_manager_xact_id( T16 ),
       .io_in_0_bits_is_builtin_type( T15 ),
       .io_in_0_bits_g_type( T13 ),
       .io_in_0_bits_data( T10 ),
       //.io_in_0_bits_client_id(  )
       .io_out_ready( io_tl_grant_ready ),
       .io_out_valid( gnt_arb_io_out_valid ),
       .io_out_bits_addr_beat( gnt_arb_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( gnt_arb_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( gnt_arb_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( gnt_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( gnt_arb_io_out_bits_g_type ),
       .io_out_bits_data( gnt_arb_io_out_bits_data )
       //.io_out_bits_client_id(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign gnt_arb.io_in_1_bits_client_id = {1{$random}};
    assign gnt_arb.io_in_0_bits_client_id = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T5 <= 1'b1;
  if(!T6 && T5 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "NASTI read error");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "NASTI write error");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else if(T22) begin
      tl_cnt_in <= T21;
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else if(T38) begin
      nasti_cnt_out <= T37;
    end
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else if(T112) begin
      tl_cnt_out <= T111;
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else if(T123) begin
      w_inflight <= 1'h0;
    end else if(T119) begin
      w_inflight <= 1'h1;
    end
  end
endmodule

module ClientTileLinkIOWrapper_1(
    output io_in_acquire_ready,
    input  io_in_acquire_valid,
    input [25:0] io_in_acquire_bits_addr_block,
    input [2:0] io_in_acquire_bits_client_xact_id,
    input [1:0] io_in_acquire_bits_addr_beat,
    input  io_in_acquire_bits_is_builtin_type,
    input [2:0] io_in_acquire_bits_a_type,
    input [16:0] io_in_acquire_bits_union,
    input [127:0] io_in_acquire_bits_data,
    input  io_in_grant_ready,
    output io_in_grant_valid,
    output[1:0] io_in_grant_bits_addr_beat,
    output[2:0] io_in_grant_bits_client_xact_id,
    output io_in_grant_bits_manager_xact_id,
    output io_in_grant_bits_is_builtin_type,
    output[3:0] io_in_grant_bits_g_type,
    output[127:0] io_in_grant_bits_data,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[25:0] io_out_acquire_bits_addr_block,
    output[2:0] io_out_acquire_bits_client_xact_id,
    output[1:0] io_out_acquire_bits_addr_beat,
    output io_out_acquire_bits_is_builtin_type,
    output[2:0] io_out_acquire_bits_a_type,
    output[16:0] io_out_acquire_bits_union,
    output[127:0] io_out_acquire_bits_data,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_addr_beat,
    input [2:0] io_out_grant_bits_client_xact_id,
    input  io_out_grant_bits_manager_xact_id,
    input  io_out_grant_bits_is_builtin_type,
    input [3:0] io_out_grant_bits_g_type,
    input [127:0] io_out_grant_bits_data,
    output io_out_probe_ready,
    input  io_out_probe_valid,
    input [25:0] io_out_probe_bits_addr_block,
    input [1:0] io_out_probe_bits_p_type,
    input  io_out_release_ready,
    output io_out_release_valid
    //output[1:0] io_out_release_bits_addr_beat
    //output[25:0] io_out_release_bits_addr_block
    //output[2:0] io_out_release_bits_client_xact_id
    //output io_out_release_bits_voluntary
    //output[2:0] io_out_release_bits_r_type
    //output[127:0] io_out_release_bits_data
);



`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_out_release_bits_data = {4{$random}};
//  assign io_out_release_bits_r_type = {1{$random}};
//  assign io_out_release_bits_voluntary = {1{$random}};
//  assign io_out_release_bits_client_xact_id = {1{$random}};
//  assign io_out_release_bits_addr_block = {1{$random}};
//  assign io_out_release_bits_addr_beat = {1{$random}};
// synthesis translate_on
`endif
  assign io_out_release_valid = 1'h0;
  assign io_out_probe_ready = 1'h1;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_acquire_ready = io_out_acquire_ready;
endmodule

module ClientTileLinkEnqueuer(
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [25:0] io_inner_acquire_bits_addr_block,
    input [2:0] io_inner_acquire_bits_client_xact_id,
    input [1:0] io_inner_acquire_bits_addr_beat,
    input  io_inner_acquire_bits_is_builtin_type,
    input [2:0] io_inner_acquire_bits_a_type,
    input [16:0] io_inner_acquire_bits_union,
    input [127:0] io_inner_acquire_bits_data,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_addr_beat,
    output[2:0] io_inner_grant_bits_client_xact_id,
    output io_inner_grant_bits_manager_xact_id,
    output io_inner_grant_bits_is_builtin_type,
    output[3:0] io_inner_grant_bits_g_type,
    output[127:0] io_inner_grant_bits_data,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[25:0] io_inner_probe_bits_addr_block,
    output[1:0] io_inner_probe_bits_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_addr_beat,
    input [25:0] io_inner_release_bits_addr_block,
    input [2:0] io_inner_release_bits_client_xact_id,
    input  io_inner_release_bits_voluntary,
    input [2:0] io_inner_release_bits_r_type,
    input [127:0] io_inner_release_bits_data,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[25:0] io_outer_acquire_bits_addr_block,
    output[2:0] io_outer_acquire_bits_client_xact_id,
    output[1:0] io_outer_acquire_bits_addr_beat,
    output io_outer_acquire_bits_is_builtin_type,
    output[2:0] io_outer_acquire_bits_a_type,
    output[16:0] io_outer_acquire_bits_union,
    output[127:0] io_outer_acquire_bits_data,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_addr_beat,
    input [2:0] io_outer_grant_bits_client_xact_id,
    input  io_outer_grant_bits_manager_xact_id,
    input  io_outer_grant_bits_is_builtin_type,
    input [3:0] io_outer_grant_bits_g_type,
    input [127:0] io_outer_grant_bits_data,
    output io_outer_probe_ready,
    input  io_outer_probe_valid,
    input [25:0] io_outer_probe_bits_addr_block,
    input [1:0] io_outer_probe_bits_p_type,
    input  io_outer_release_ready,
    output io_outer_release_valid,
    output[1:0] io_outer_release_bits_addr_beat,
    output[25:0] io_outer_release_bits_addr_block,
    output[2:0] io_outer_release_bits_client_xact_id,
    output io_outer_release_bits_voluntary,
    output[2:0] io_outer_release_bits_r_type,
    output[127:0] io_outer_release_bits_data
);



  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_acquire_ready = io_outer_acquire_ready;
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [7:0] io_enq_bits_strb,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[7:0] io_deq_bits_strb,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T23;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T24;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T25;
  wire T8;
  wire T9;
  wire T10;
  wire[73:0] T11;
  reg [73:0] ram [7:0];
  wire[73:0] T12;
  wire[73:0] T13;
  wire[73:0] T14;
  wire[8:0] T15;
  wire[64:0] T16;
  wire[7:0] T17;
  wire T18;
  wire[63:0] T19;
  wire T20;
  wire empty;
  wire T21;
  wire T22;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T23 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T24 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T25 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T16, T15};
  assign T15 = {io_enq_bits_strb, io_enq_bits_user};
  assign T16 = {io_enq_bits_data, io_enq_bits_last};
  assign io_deq_bits_strb = T17;
  assign T17 = T11[4'h8:1'h1];
  assign io_deq_bits_last = T18;
  assign T18 = T11[4'h9:4'h9];
  assign io_deq_bits_data = T19;
  assign T19 = T11[7'h49:4'ha];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [63:0] io_enq_bits_data,
    input  io_enq_bits_last,
    input [3:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[63:0] io_deq_bits_data,
    output io_deq_bits_last,
    output[3:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[3:0] io_count
);

  wire[3:0] T0;
  wire[2:0] ptr_diff;
  reg [2:0] R1;
  wire[2:0] T25;
  wire[2:0] T2;
  wire[2:0] T3;
  wire do_deq;
  reg [2:0] R4;
  wire[2:0] T26;
  wire[2:0] T5;
  wire[2:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T27;
  wire T8;
  wire T9;
  wire T10;
  wire[71:0] T11;
  reg [71:0] ram [7:0];
  wire[71:0] T12;
  wire[71:0] T13;
  wire[71:0] T14;
  wire[5:0] T15;
  wire[4:0] T16;
  wire[65:0] T17;
  wire[3:0] T18;
  wire T19;
  wire[63:0] T20;
  wire[1:0] T21;
  wire T22;
  wire empty;
  wire T23;
  wire T24;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T25 = reset ? 3'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 3'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T26 = reset ? 3'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 3'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T27 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T17, T15};
  assign T15 = {io_enq_bits_last, T16};
  assign T16 = {io_enq_bits_id, io_enq_bits_user};
  assign T17 = {io_enq_bits_resp, io_enq_bits_data};
  assign io_deq_bits_id = T18;
  assign T18 = T11[3'h4:1'h1];
  assign io_deq_bits_last = T19;
  assign T19 = T11[3'h5:3'h5];
  assign io_deq_bits_data = T20;
  assign T20 = T11[7'h45:3'h6];
  assign io_deq_bits_resp = T21;
  assign T21 = T11[7'h47:7'h46];
  assign io_deq_valid = T22;
  assign T22 = empty ^ 1'h1;
  assign empty = ptr_match & T23;
  assign T23 = maybe_full ^ 1'h1;
  assign io_enq_ready = T24;
  assign T24 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 3'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 3'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_resp,
    input [3:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_resp,
    output[3:0] io_deq_bits_id,
    output io_deq_bits_user,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire T10;
  wire[6:0] T11;
  reg [6:0] ram [1:0];
  wire[6:0] T12;
  wire[6:0] T13;
  wire[6:0] T14;
  wire[4:0] T15;
  wire[3:0] T16;
  wire[1:0] T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_user = T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_resp, T15};
  assign T15 = {io_enq_bits_id, io_enq_bits_user};
  assign io_deq_bits_id = T16;
  assign T16 = T11[3'h4:1'h1];
  assign io_deq_bits_resp = T17;
  assign T17 = T11[3'h6:3'h5];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module RTC(input clk, input reset,
    input  io_aw_ready,
    output io_aw_valid,
    output[31:0] io_aw_bits_addr,
    output[7:0] io_aw_bits_len,
    output[2:0] io_aw_bits_size,
    output[1:0] io_aw_bits_burst,
    output io_aw_bits_lock,
    output[3:0] io_aw_bits_cache,
    output[2:0] io_aw_bits_prot,
    output[3:0] io_aw_bits_qos,
    output[3:0] io_aw_bits_region,
    output[3:0] io_aw_bits_id,
    output io_aw_bits_user,
    input  io_w_ready,
    output io_w_valid,
    output[63:0] io_w_bits_data,
    output io_w_bits_last,
    output[7:0] io_w_bits_strb,
    output io_w_bits_user,
    output io_b_ready,
    input  io_b_valid,
    input [1:0] io_b_bits_resp,
    input [3:0] io_b_bits_id,
    input  io_b_bits_user,
    input  io_ar_ready,
    output io_ar_valid,
    //output[31:0] io_ar_bits_addr
    //output[7:0] io_ar_bits_len
    //output[2:0] io_ar_bits_size
    //output[1:0] io_ar_bits_burst
    //output io_ar_bits_lock
    //output[3:0] io_ar_bits_cache
    //output[2:0] io_ar_bits_prot
    //output[3:0] io_ar_bits_qos
    //output[3:0] io_ar_bits_region
    //output[3:0] io_ar_bits_id
    //output io_ar_bits_user
    output io_r_ready,
    input  io_r_valid,
    input [1:0] io_r_bits_resp,
    input [63:0] io_r_bits_data,
    input  io_r_bits_last,
    input [3:0] io_r_bits_id,
    input  io_r_bits_user
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  reg  send_acked_0;
  wire T39;
  wire T3;
  wire T4;
  wire rtc_tick;
  reg [6:0] R5;
  wire[6:0] T40;
  wire[6:0] T6;
  wire[6:0] T7;
  wire T8;
  wire T9;
  wire[1:0] T10;
  wire T11;
  wire T41;
  wire T12;
  wire T13;
  wire T14;
  wire[7:0] T15;
  wire T16;
  wire[63:0] T17;
  reg [63:0] rtc;
  wire[63:0] T42;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  sending_data;
  wire T43;
  wire T20;
  wire T21;
  wire[3:0] T22;
  wire[3:0] T44;
  wire coreId;
  wire[3:0] T23;
  wire[3:0] T24;
  wire[2:0] T25;
  wire[3:0] T26;
  wire T27;
  wire[1:0] T28;
  wire[2:0] T29;
  wire[7:0] T30;
  wire[31:0] T31;
  wire[31:0] T45;
  reg [30:0] T32;
  reg  sending_addr;
  wire T46;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    send_acked_0 = {1{$random}};
    R5 = {1{$random}};
    rtc = {2{$random}};
    sending_data = {1{$random}};
    sending_addr = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_ar_bits_user = {1{$random}};
//  assign io_ar_bits_id = {1{$random}};
//  assign io_ar_bits_region = {1{$random}};
//  assign io_ar_bits_qos = {1{$random}};
//  assign io_ar_bits_prot = {1{$random}};
//  assign io_ar_bits_cache = {1{$random}};
//  assign io_ar_bits_lock = {1{$random}};
//  assign io_ar_bits_burst = {1{$random}};
//  assign io_ar_bits_size = {1{$random}};
//  assign io_ar_bits_len = {1{$random}};
//  assign io_ar_bits_addr = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T13 | send_acked_0;
  assign T39 = reset ? 1'h1 : T3;
  assign T3 = T8 ? 1'h1 : T4;
  assign T4 = rtc_tick ? 1'h0 : send_acked_0;
  assign rtc_tick = R5 == 7'h63;
  assign T40 = reset ? 7'h0 : T6;
  assign T6 = rtc_tick ? 7'h0 : T7;
  assign T7 = R5 + 7'h1;
  assign T8 = T12 & T9;
  assign T9 = T10[1'h0:1'h0];
  assign T10 = 1'h1 << T11;
  assign T11 = T41;
  assign T41 = io_b_bits_id[1'h0:1'h0];
  assign T12 = io_b_ready & io_b_valid;
  assign T13 = rtc_tick ^ 1'h1;
  assign io_r_ready = 1'h0;
  assign io_ar_valid = 1'h0;
  assign io_b_ready = 1'h1;
  assign io_w_bits_user = T14;
  assign T14 = 1'h0;
  assign io_w_bits_strb = T15;
  assign T15 = 8'hff;
  assign io_w_bits_last = T16;
  assign T16 = 1'h1;
  assign io_w_bits_data = T17;
  assign T17 = rtc;
  assign T42 = reset ? 64'h0 : T18;
  assign T18 = rtc_tick ? T19 : rtc;
  assign T19 = rtc + 64'h1;
  assign io_w_valid = sending_data;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = rtc_tick ? 1'h1 : sending_data;
  assign io_aw_bits_user = T21;
  assign T21 = 1'h0;
  assign io_aw_bits_id = T22;
  assign T22 = T44;
  assign T44 = {3'h0, coreId};
  assign coreId = 1'h0;
  assign io_aw_bits_region = T23;
  assign T23 = 4'h0;
  assign io_aw_bits_qos = T24;
  assign T24 = 4'h0;
  assign io_aw_bits_prot = T25;
  assign T25 = 3'h0;
  assign io_aw_bits_cache = T26;
  assign T26 = 4'h0;
  assign io_aw_bits_lock = T27;
  assign T27 = 1'h0;
  assign io_aw_bits_burst = T28;
  assign T28 = 2'h1;
  assign io_aw_bits_size = T29;
  assign T29 = 3'h3;
  assign io_aw_bits_len = T30;
  assign T30 = 8'h0;
  assign io_aw_bits_addr = T31;
  assign T31 = T45;
  assign T45 = {1'h0, T32};
  always @(*) case (coreId)
    0: T32 = 31'h4000b808;
    default: begin
      T32 = 31'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      T32 = {1{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign io_aw_valid = sending_addr;
  assign T46 = reset ? 1'h0 : T34;
  assign T34 = T38 ? 1'h0 : T35;
  assign T35 = T37 ? 1'h0 : T36;
  assign T36 = rtc_tick ? 1'h1 : sending_addr;
  assign T37 = io_aw_ready & io_aw_valid;
  assign T38 = io_w_ready & io_w_valid;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Not all clocks were updated for rtc tick");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      send_acked_0 <= 1'h1;
    end else if(T8) begin
      send_acked_0 <= 1'h1;
    end else if(rtc_tick) begin
      send_acked_0 <= 1'h0;
    end
    if(reset) begin
      R5 <= 7'h0;
    end else if(rtc_tick) begin
      R5 <= 7'h0;
    end else begin
      R5 <= T7;
    end
    if(reset) begin
      rtc <= 64'h0;
    end else if(rtc_tick) begin
      rtc <= T19;
    end
    if(reset) begin
      sending_data <= 1'h0;
    end else if(rtc_tick) begin
      sending_data <= 1'h1;
    end
    if(reset) begin
      sending_addr <= 1'h0;
    end else if(T38) begin
      sending_addr <= 1'h0;
    end else if(T37) begin
      sending_addr <= 1'h0;
    end else if(rtc_tick) begin
      sending_addr <= 1'h1;
    end
  end
endmodule

module SMIIONastiReadIOConverter_0(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [3:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[3:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [11:0] addr;
  wire[11:0] T22;
  wire[11:0] T23;
  wire[11:0] T24;
  wire[11:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  reg [3:0] id;
  wire[3:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0:1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'he:2'h3];
  assign T25 = addr + 12'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0:1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SMIIONastiWriteIOConverter_0(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [3:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[3:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [11:0] addr;
  wire[11:0] T39;
  wire[11:0] T40;
  wire[11:0] T41;
  wire[11:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[3:0] T46;
  reg [3:0] id;
  wire[3:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0:1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'he:2'h3];
  assign T42 = addr + 12'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= SMI size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [11:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [11:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[11:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[11:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SMIArbiter_0(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [11:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [11:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[11:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[11:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_0 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SMIIONastiIOConverter_0(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [3:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[3:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [3:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[3:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[11:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[3:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[11:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[3:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[11:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[11:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SMIIONastiReadIOConverter_0 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SMIIONastiWriteIOConverter_0 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SMIArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module SMIIONastiReadIOConverter_1(input clk, input reset,
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [3:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[3:0] io_r_bits_id,
    output io_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    //output[63:0] io_smi_req_bits_data
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire T0;
  reg [1:0] state;
  wire[1:0] T60;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  wire T6;
  reg  nWords;
  wire T61;
  wire[7:0] T7;
  wire[7:0] T62;
  wire T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[2:0] T13;
  wire T14;
  wire T15;
  reg  recvInd;
  wire T63;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire T21;
  reg [5:0] addr;
  wire[5:0] T22;
  wire[5:0] T23;
  wire[5:0] T24;
  wire[5:0] T25;
  wire T26;
  wire T27;
  wire T28;
  reg  sendDone;
  wire T64;
  wire T29;
  wire T30;
  wire T31;
  reg  sendInd;
  wire T65;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  reg [3:0] id;
  wire[3:0] T38;
  wire T39;
  wire T40;
  reg [7:0] nBeats;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  reg [63:0] buffer_0;
  wire[63:0] T66;
  wire[63:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[5:0] T49;
  reg [2:0] byteOff;
  wire[2:0] T50;
  wire[2:0] T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire[1:0] T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    nWords = {1{$random}};
    recvInd = {1{$random}};
    addr = {1{$random}};
    sendDone = {1{$random}};
    sendInd = {1{$random}};
    id = {1{$random}};
    nBeats = {1{$random}};
    buffer_0 = {2{$random}};
    byteOff = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_smi_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
  assign io_smi_resp_ready = T0;
  assign T0 = state == 2'h1;
  assign T60 = reset ? 2'h0 : T1;
  assign T1 = T21 ? T20 : T2;
  assign T2 = T5 ? 2'h2 : T3;
  assign T3 = T4 ? 2'h1 : state;
  assign T4 = io_ar_ready & io_ar_valid;
  assign T5 = T19 & T6;
  assign T6 = recvInd == nWords;
  assign T61 = T7[1'h0:1'h0];
  assign T7 = T14 ? T11 : T62;
  assign T62 = {7'h0, T8};
  assign T8 = T9 ? 1'h0 : nWords;
  assign T9 = T4 & T10;
  assign T10 = io_ar_bits_size < 3'h3;
  assign T11 = T12 - 8'h1;
  assign T12 = 1'h1 << T13;
  assign T13 = io_ar_bits_size - 3'h3;
  assign T14 = T4 & T15;
  assign T15 = T10 ^ 1'h1;
  assign T63 = reset ? 1'h0 : T16;
  assign T16 = T21 ? 1'h0 : T17;
  assign T17 = T19 ? T18 : recvInd;
  assign T18 = recvInd + 1'h1;
  assign T19 = io_smi_resp_ready & io_smi_resp_valid;
  assign T20 = io_r_bits_last ? 2'h0 : 2'h1;
  assign T21 = io_r_ready & io_r_valid;
  assign io_smi_req_bits_addr = addr;
  assign T22 = T26 ? T25 : T23;
  assign T23 = T4 ? T24 : addr;
  assign T24 = io_ar_bits_addr[4'h8:2'h3];
  assign T25 = addr + 6'h1;
  assign T26 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_req_bits_rw = 1'h0;
  assign io_smi_req_valid = T27;
  assign T27 = T35 & T28;
  assign T28 = sendDone ^ 1'h1;
  assign T64 = reset ? 1'h0 : T29;
  assign T29 = T21 ? 1'h0 : T30;
  assign T30 = T26 ? T31 : sendDone;
  assign T31 = sendInd == nWords;
  assign T65 = reset ? 1'h0 : T32;
  assign T32 = T21 ? 1'h0 : T33;
  assign T33 = T26 ? T34 : sendInd;
  assign T34 = sendInd + 1'h1;
  assign T35 = state == 2'h1;
  assign io_r_bits_user = T36;
  assign T36 = 1'h0;
  assign io_r_bits_id = T37;
  assign T37 = id;
  assign T38 = T4 ? io_ar_bits_id : id;
  assign io_r_bits_last = T39;
  assign T39 = T40;
  assign T40 = nBeats == 8'h0;
  assign T41 = T21 ? T43 : T42;
  assign T42 = T4 ? io_ar_bits_len : nBeats;
  assign T43 = nBeats - 8'h1;
  assign io_r_bits_data = T44;
  assign T44 = T45;
  assign T45 = buffer_0;
  assign T66 = reset ? 64'h0 : T46;
  assign T46 = T21 ? 64'h0 : T47;
  assign T47 = T53 ? T48 : buffer_0;
  assign T48 = io_smi_resp_bits >> T49;
  assign T49 = {byteOff, 3'h0};
  assign T50 = T14 ? 3'h0 : T51;
  assign T51 = T9 ? T52 : byteOff;
  assign T52 = io_ar_bits_addr[2'h2:1'h0];
  assign T53 = T19 & T54;
  assign T54 = T55[1'h0:1'h0];
  assign T55 = 1'h1 << T56;
  assign T56 = recvInd;
  assign io_r_bits_resp = T57;
  assign T57 = 2'h0;
  assign io_r_valid = T58;
  assign T58 = state == 2'h2;
  assign io_ar_ready = T59;
  assign T59 = state == 2'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T21) begin
      state <= T20;
    end else if(T5) begin
      state <= 2'h2;
    end else if(T4) begin
      state <= 2'h1;
    end
    nWords <= T61;
    if(reset) begin
      recvInd <= 1'h0;
    end else if(T21) begin
      recvInd <= 1'h0;
    end else if(T19) begin
      recvInd <= T18;
    end
    if(T26) begin
      addr <= T25;
    end else if(T4) begin
      addr <= T24;
    end
    if(reset) begin
      sendDone <= 1'h0;
    end else if(T21) begin
      sendDone <= 1'h0;
    end else if(T26) begin
      sendDone <= T31;
    end
    if(reset) begin
      sendInd <= 1'h0;
    end else if(T21) begin
      sendInd <= 1'h0;
    end else if(T26) begin
      sendInd <= T34;
    end
    if(T4) begin
      id <= io_ar_bits_id;
    end
    if(T21) begin
      nBeats <= T43;
    end else if(T4) begin
      nBeats <= io_ar_bits_len;
    end
    if(reset) begin
      buffer_0 <= 64'h0;
    end else if(T21) begin
      buffer_0 <= 64'h0;
    end else if(T53) begin
      buffer_0 <= T48;
    end
    if(T14) begin
      byteOff <= 3'h0;
    end else if(T9) begin
      byteOff <= T52;
    end
  end
endmodule

module SMIIONastiWriteIOConverter_1(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [3:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    output[1:0] io_b_bits_resp,
    output[3:0] io_b_bits_id,
    output io_b_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  reg [2:0] state;
  wire[2:0] T52;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  reg  last;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg  strb;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[255:0] T22;
  wire[255:0] T53;
  wire[255:0] T23;
  wire[255:0] T24;
  wire[7:0] T25;
  reg [2:0] size;
  wire[2:0] T26;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  reg [63:0] data;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [5:0] addr;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire[3:0] T46;
  reg [3:0] id;
  wire[3:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire T51;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    state = {1{$random}};
    last = {1{$random}};
    strb = {1{$random}};
    size = {1{$random}};
    data = {2{$random}};
    addr = {1{$random}};
    id = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T4 | T3;
  assign T3 = 3'h3 <= io_aw_bits_size;
  assign T4 = io_aw_valid ^ 1'h1;
  assign io_smi_resp_ready = T5;
  assign T5 = state == 3'h3;
  assign T52 = reset ? 3'h0 : T6;
  assign T6 = T35 ? 3'h0 : T7;
  assign T7 = T34 ? 3'h4 : T8;
  assign T8 = T16 ? T13 : T9;
  assign T9 = T12 ? 3'h2 : T10;
  assign T10 = T11 ? 3'h1 : state;
  assign T11 = io_aw_ready & io_aw_valid;
  assign T12 = io_w_ready & io_w_valid;
  assign T13 = last ? 3'h3 : 3'h1;
  assign T14 = T12 ? io_w_bits_last : T15;
  assign T15 = T11 ? 1'h0 : last;
  assign T16 = T33 & T17;
  assign T17 = strb == 1'h0;
  assign T18 = T28 ? 1'h0 : T19;
  assign T19 = T12 ? T20 : strb;
  assign T20 = T21;
  assign T21 = T22[1'h0:1'h0];
  assign T22 = T23 & T53;
  assign T53 = {248'h0, io_w_bits_strb};
  assign T23 = T24 - 256'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = 1'h1 << size;
  assign T26 = T11 ? io_aw_bits_size : size;
  assign T28 = T33 & T29;
  assign T29 = T32 & T30;
  assign T30 = io_smi_req_ready | T31;
  assign T31 = strb ^ 1'h1;
  assign T32 = T17 ^ 1'h1;
  assign T33 = state == 3'h2;
  assign T34 = io_smi_resp_ready & io_smi_resp_valid;
  assign T35 = io_b_ready & io_b_valid;
  assign io_smi_req_bits_data = data;
  assign T36 = T28 ? 64'h0 : T37;
  assign T37 = T12 ? io_w_bits_data : data;
  assign io_smi_req_bits_addr = addr;
  assign T39 = T28 ? T42 : T40;
  assign T40 = T11 ? T41 : addr;
  assign T41 = io_aw_bits_addr[4'h8:2'h3];
  assign T42 = addr + 6'h1;
  assign io_smi_req_bits_rw = 1'h1;
  assign io_smi_req_valid = T43;
  assign T43 = T44 & strb;
  assign T44 = state == 3'h2;
  assign io_b_bits_user = T45;
  assign T45 = 1'h0;
  assign io_b_bits_id = T46;
  assign T46 = id;
  assign T47 = T11 ? io_aw_bits_id : id;
  assign io_b_bits_resp = T48;
  assign T48 = 2'h0;
  assign io_b_valid = T49;
  assign T49 = state == 3'h4;
  assign io_w_ready = T50;
  assign T50 = state == 3'h1;
  assign io_aw_ready = T51;
  assign T51 = state == 3'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Nasti size must be >= SMI size");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      state <= 3'h0;
    end else if(T35) begin
      state <= 3'h0;
    end else if(T34) begin
      state <= 3'h4;
    end else if(T16) begin
      state <= T13;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T11) begin
      state <= 3'h1;
    end
    if(T12) begin
      last <= io_w_bits_last;
    end else if(T11) begin
      last <= 1'h0;
    end
    if(T28) begin
      strb <= 1'h0;
    end else if(T12) begin
      strb <= T20;
    end
    if(T11) begin
      size <= io_aw_bits_size;
    end
    if(T28) begin
      data <= 64'h0;
    end else if(T12) begin
      data <= io_w_bits_data;
    end
    if(T28) begin
      addr <= T42;
    end else if(T11) begin
      addr <= T41;
    end
    if(T11) begin
      id <= io_aw_bits_id;
    end
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_rw,
    input [5:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_rw,
    input [5:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_rw,
    output[5:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T27;
  wire T3;
  wire T4;
  wire[63:0] T5;
  wire T6;
  wire[5:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T27 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_data = T5;
  assign T5 = T6 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T6 = chosen;
  assign io_out_bits_addr = T7;
  assign T7 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_rw = T8;
  assign T8 = T6 ? io_in_1_bits_rw : io_in_0_bits_rw;
  assign io_out_valid = T9;
  assign T9 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = T18 | T12;
  assign T12 = T13 ^ 1'h1;
  assign T13 = T16 | T14;
  assign T14 = io_in_1_valid & T15;
  assign T15 = last_grant < 1'h1;
  assign T16 = io_in_0_valid & T17;
  assign T17 = last_grant < 1'h0;
  assign T18 = last_grant < 1'h0;
  assign io_in_1_ready = T19;
  assign T19 = T20 & io_out_ready;
  assign T20 = T24 | T21;
  assign T21 = T22 ^ 1'h1;
  assign T22 = T23 | io_in_0_valid;
  assign T23 = T16 | T14;
  assign T24 = T26 & T25;
  assign T25 = last_grant < 1'h1;
  assign T26 = T16 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module SMIArbiter_1(input clk, input reset,
    output io_in_1_req_ready,
    input  io_in_1_req_valid,
    input  io_in_1_req_bits_rw,
    input [5:0] io_in_1_req_bits_addr,
    input [63:0] io_in_1_req_bits_data,
    input  io_in_1_resp_ready,
    output io_in_1_resp_valid,
    output[63:0] io_in_1_resp_bits,
    output io_in_0_req_ready,
    input  io_in_0_req_valid,
    input  io_in_0_req_bits_rw,
    input [5:0] io_in_0_req_bits_addr,
    input [63:0] io_in_0_req_bits_data,
    input  io_in_0_resp_ready,
    output io_in_0_resp_valid,
    output[63:0] io_in_0_resp_bits,
    input  io_out_req_ready,
    output io_out_req_valid,
    output io_out_req_bits_rw,
    output[5:0] io_out_req_bits_addr,
    output[63:0] io_out_req_bits_data,
    output io_out_resp_ready,
    input  io_out_resp_valid,
    input [63:0] io_out_resp_bits
);

  wire T0;
  wire T1;
  reg  wait_resp;
  wire T15;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  choice;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire req_arb_io_in_1_ready;
  wire req_arb_io_in_0_ready;
  wire req_arb_io_out_valid;
  wire req_arb_io_out_bits_rw;
  wire[5:0] req_arb_io_out_bits_addr;
  wire[63:0] req_arb_io_out_bits_data;
  wire req_arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wait_resp = {1{$random}};
    choice = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_out_req_ready & T1;
  assign T1 = wait_resp ^ 1'h1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = T5 ? 1'h0 : T3;
  assign T3 = T4 ? 1'h1 : wait_resp;
  assign T4 = io_out_req_ready & io_out_req_valid;
  assign T5 = io_out_resp_ready & io_out_resp_valid;
  assign io_out_resp_ready = T6;
  assign T6 = T7 ? io_in_1_resp_ready : io_in_0_resp_ready;
  assign T7 = choice;
  assign T8 = T4 ? req_arb_io_chosen : choice;
  assign io_out_req_bits_data = req_arb_io_out_bits_data;
  assign io_out_req_bits_addr = req_arb_io_out_bits_addr;
  assign io_out_req_bits_rw = req_arb_io_out_bits_rw;
  assign io_out_req_valid = T9;
  assign T9 = req_arb_io_out_valid & T10;
  assign T10 = wait_resp ^ 1'h1;
  assign io_in_0_resp_bits = io_out_resp_bits;
  assign io_in_0_resp_valid = T11;
  assign T11 = io_out_resp_valid & T12;
  assign T12 = choice == 1'h0;
  assign io_in_0_req_ready = req_arb_io_in_0_ready;
  assign io_in_1_resp_bits = io_out_resp_bits;
  assign io_in_1_resp_valid = T13;
  assign T13 = io_out_resp_valid & T14;
  assign T14 = choice == 1'h1;
  assign io_in_1_req_ready = req_arb_io_in_1_ready;
  RRArbiter_1 req_arb(.clk(clk), .reset(reset),
       .io_in_1_ready( req_arb_io_in_1_ready ),
       .io_in_1_valid( io_in_1_req_valid ),
       .io_in_1_bits_rw( io_in_1_req_bits_rw ),
       .io_in_1_bits_addr( io_in_1_req_bits_addr ),
       .io_in_1_bits_data( io_in_1_req_bits_data ),
       .io_in_0_ready( req_arb_io_in_0_ready ),
       .io_in_0_valid( io_in_0_req_valid ),
       .io_in_0_bits_rw( io_in_0_req_bits_rw ),
       .io_in_0_bits_addr( io_in_0_req_bits_addr ),
       .io_in_0_bits_data( io_in_0_req_bits_data ),
       .io_out_ready( T0 ),
       .io_out_valid( req_arb_io_out_valid ),
       .io_out_bits_rw( req_arb_io_out_bits_rw ),
       .io_out_bits_addr( req_arb_io_out_bits_addr ),
       .io_out_bits_data( req_arb_io_out_bits_data ),
       .io_chosen( req_arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      wait_resp <= 1'h0;
    end else if(T5) begin
      wait_resp <= 1'h0;
    end else if(T4) begin
      wait_resp <= 1'h1;
    end
    if(T4) begin
      choice <= req_arb_io_chosen;
    end
  end
endmodule

module SMIIONastiIOConverter_1(input clk, input reset,
    output io_nasti_aw_ready,
    input  io_nasti_aw_valid,
    input [31:0] io_nasti_aw_bits_addr,
    input [7:0] io_nasti_aw_bits_len,
    input [2:0] io_nasti_aw_bits_size,
    input [1:0] io_nasti_aw_bits_burst,
    input  io_nasti_aw_bits_lock,
    input [3:0] io_nasti_aw_bits_cache,
    input [2:0] io_nasti_aw_bits_prot,
    input [3:0] io_nasti_aw_bits_qos,
    input [3:0] io_nasti_aw_bits_region,
    input [3:0] io_nasti_aw_bits_id,
    input  io_nasti_aw_bits_user,
    output io_nasti_w_ready,
    input  io_nasti_w_valid,
    input [63:0] io_nasti_w_bits_data,
    input  io_nasti_w_bits_last,
    input [7:0] io_nasti_w_bits_strb,
    input  io_nasti_w_bits_user,
    input  io_nasti_b_ready,
    output io_nasti_b_valid,
    output[1:0] io_nasti_b_bits_resp,
    output[3:0] io_nasti_b_bits_id,
    output io_nasti_b_bits_user,
    output io_nasti_ar_ready,
    input  io_nasti_ar_valid,
    input [31:0] io_nasti_ar_bits_addr,
    input [7:0] io_nasti_ar_bits_len,
    input [2:0] io_nasti_ar_bits_size,
    input [1:0] io_nasti_ar_bits_burst,
    input  io_nasti_ar_bits_lock,
    input [3:0] io_nasti_ar_bits_cache,
    input [2:0] io_nasti_ar_bits_prot,
    input [3:0] io_nasti_ar_bits_qos,
    input [3:0] io_nasti_ar_bits_region,
    input [3:0] io_nasti_ar_bits_id,
    input  io_nasti_ar_bits_user,
    input  io_nasti_r_ready,
    output io_nasti_r_valid,
    output[1:0] io_nasti_r_bits_resp,
    output[63:0] io_nasti_r_bits_data,
    output io_nasti_r_bits_last,
    output[3:0] io_nasti_r_bits_id,
    output io_nasti_r_bits_user,
    input  io_smi_req_ready,
    output io_smi_req_valid,
    output io_smi_req_bits_rw,
    output[5:0] io_smi_req_bits_addr,
    output[63:0] io_smi_req_bits_data,
    output io_smi_resp_ready,
    input  io_smi_resp_valid,
    input [63:0] io_smi_resp_bits
);

  wire reader_io_ar_ready;
  wire reader_io_r_valid;
  wire[1:0] reader_io_r_bits_resp;
  wire[63:0] reader_io_r_bits_data;
  wire reader_io_r_bits_last;
  wire[3:0] reader_io_r_bits_id;
  wire reader_io_r_bits_user;
  wire reader_io_smi_req_valid;
  wire reader_io_smi_req_bits_rw;
  wire[5:0] reader_io_smi_req_bits_addr;
  wire reader_io_smi_resp_ready;
  wire writer_io_aw_ready;
  wire writer_io_w_ready;
  wire writer_io_b_valid;
  wire[1:0] writer_io_b_bits_resp;
  wire[3:0] writer_io_b_bits_id;
  wire writer_io_b_bits_user;
  wire writer_io_smi_req_valid;
  wire writer_io_smi_req_bits_rw;
  wire[5:0] writer_io_smi_req_bits_addr;
  wire[63:0] writer_io_smi_req_bits_data;
  wire writer_io_smi_resp_ready;
  wire arb_io_in_1_req_ready;
  wire arb_io_in_1_resp_valid;
  wire[63:0] arb_io_in_1_resp_bits;
  wire arb_io_in_0_req_ready;
  wire arb_io_in_0_resp_valid;
  wire[63:0] arb_io_in_0_resp_bits;
  wire arb_io_out_req_valid;
  wire arb_io_out_req_bits_rw;
  wire[5:0] arb_io_out_req_bits_addr;
  wire[63:0] arb_io_out_req_bits_data;
  wire arb_io_out_resp_ready;


  assign io_smi_resp_ready = arb_io_out_resp_ready;
  assign io_smi_req_bits_data = arb_io_out_req_bits_data;
  assign io_smi_req_bits_addr = arb_io_out_req_bits_addr;
  assign io_smi_req_bits_rw = arb_io_out_req_bits_rw;
  assign io_smi_req_valid = arb_io_out_req_valid;
  assign io_nasti_r_bits_user = reader_io_r_bits_user;
  assign io_nasti_r_bits_id = reader_io_r_bits_id;
  assign io_nasti_r_bits_last = reader_io_r_bits_last;
  assign io_nasti_r_bits_data = reader_io_r_bits_data;
  assign io_nasti_r_bits_resp = reader_io_r_bits_resp;
  assign io_nasti_r_valid = reader_io_r_valid;
  assign io_nasti_ar_ready = reader_io_ar_ready;
  assign io_nasti_b_bits_user = writer_io_b_bits_user;
  assign io_nasti_b_bits_id = writer_io_b_bits_id;
  assign io_nasti_b_bits_resp = writer_io_b_bits_resp;
  assign io_nasti_b_valid = writer_io_b_valid;
  assign io_nasti_w_ready = writer_io_w_ready;
  assign io_nasti_aw_ready = writer_io_aw_ready;
  SMIIONastiReadIOConverter_1 reader(.clk(clk), .reset(reset),
       .io_ar_ready( reader_io_ar_ready ),
       .io_ar_valid( io_nasti_ar_valid ),
       .io_ar_bits_addr( io_nasti_ar_bits_addr ),
       .io_ar_bits_len( io_nasti_ar_bits_len ),
       .io_ar_bits_size( io_nasti_ar_bits_size ),
       .io_ar_bits_burst( io_nasti_ar_bits_burst ),
       .io_ar_bits_lock( io_nasti_ar_bits_lock ),
       .io_ar_bits_cache( io_nasti_ar_bits_cache ),
       .io_ar_bits_prot( io_nasti_ar_bits_prot ),
       .io_ar_bits_qos( io_nasti_ar_bits_qos ),
       .io_ar_bits_region( io_nasti_ar_bits_region ),
       .io_ar_bits_id( io_nasti_ar_bits_id ),
       .io_ar_bits_user( io_nasti_ar_bits_user ),
       .io_r_ready( io_nasti_r_ready ),
       .io_r_valid( reader_io_r_valid ),
       .io_r_bits_resp( reader_io_r_bits_resp ),
       .io_r_bits_data( reader_io_r_bits_data ),
       .io_r_bits_last( reader_io_r_bits_last ),
       .io_r_bits_id( reader_io_r_bits_id ),
       .io_r_bits_user( reader_io_r_bits_user ),
       .io_smi_req_ready( arb_io_in_0_req_ready ),
       .io_smi_req_valid( reader_io_smi_req_valid ),
       .io_smi_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_smi_req_bits_data(  )
       .io_smi_resp_ready( reader_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_0_resp_valid ),
       .io_smi_resp_bits( arb_io_in_0_resp_bits )
  );
  SMIIONastiWriteIOConverter_1 writer(.clk(clk), .reset(reset),
       .io_aw_ready( writer_io_aw_ready ),
       .io_aw_valid( io_nasti_aw_valid ),
       .io_aw_bits_addr( io_nasti_aw_bits_addr ),
       .io_aw_bits_len( io_nasti_aw_bits_len ),
       .io_aw_bits_size( io_nasti_aw_bits_size ),
       .io_aw_bits_burst( io_nasti_aw_bits_burst ),
       .io_aw_bits_lock( io_nasti_aw_bits_lock ),
       .io_aw_bits_cache( io_nasti_aw_bits_cache ),
       .io_aw_bits_prot( io_nasti_aw_bits_prot ),
       .io_aw_bits_qos( io_nasti_aw_bits_qos ),
       .io_aw_bits_region( io_nasti_aw_bits_region ),
       .io_aw_bits_id( io_nasti_aw_bits_id ),
       .io_aw_bits_user( io_nasti_aw_bits_user ),
       .io_w_ready( writer_io_w_ready ),
       .io_w_valid( io_nasti_w_valid ),
       .io_w_bits_data( io_nasti_w_bits_data ),
       .io_w_bits_last( io_nasti_w_bits_last ),
       .io_w_bits_strb( io_nasti_w_bits_strb ),
       .io_w_bits_user( io_nasti_w_bits_user ),
       .io_b_ready( io_nasti_b_ready ),
       .io_b_valid( writer_io_b_valid ),
       .io_b_bits_resp( writer_io_b_bits_resp ),
       .io_b_bits_id( writer_io_b_bits_id ),
       .io_b_bits_user( writer_io_b_bits_user ),
       .io_smi_req_ready( arb_io_in_1_req_ready ),
       .io_smi_req_valid( writer_io_smi_req_valid ),
       .io_smi_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( writer_io_smi_req_bits_data ),
       .io_smi_resp_ready( writer_io_smi_resp_ready ),
       .io_smi_resp_valid( arb_io_in_1_resp_valid ),
       .io_smi_resp_bits( arb_io_in_1_resp_bits )
  );
  SMIArbiter_1 arb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( arb_io_in_1_req_ready ),
       .io_in_1_req_valid( writer_io_smi_req_valid ),
       .io_in_1_req_bits_rw( writer_io_smi_req_bits_rw ),
       .io_in_1_req_bits_addr( writer_io_smi_req_bits_addr ),
       .io_in_1_req_bits_data( writer_io_smi_req_bits_data ),
       .io_in_1_resp_ready( writer_io_smi_resp_ready ),
       .io_in_1_resp_valid( arb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( arb_io_in_1_resp_bits ),
       .io_in_0_req_ready( arb_io_in_0_req_ready ),
       .io_in_0_req_valid( reader_io_smi_req_valid ),
       .io_in_0_req_bits_rw( reader_io_smi_req_bits_rw ),
       .io_in_0_req_bits_addr( reader_io_smi_req_bits_addr ),
       //.io_in_0_req_bits_data(  )
       .io_in_0_resp_ready( reader_io_smi_resp_ready ),
       .io_in_0_resp_valid( arb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( arb_io_in_0_resp_bits ),
       .io_out_req_ready( io_smi_req_ready ),
       .io_out_req_valid( arb_io_out_req_valid ),
       .io_out_req_bits_rw( arb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( arb_io_out_req_bits_addr ),
       .io_out_req_bits_data( arb_io_out_req_bits_data ),
       .io_out_resp_ready( arb_io_out_resp_ready ),
       .io_out_resp_valid( io_smi_resp_valid ),
       .io_out_resp_bits( io_smi_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign arb.io_in_0_req_bits_data = {2{$random}};
// synthesis translate_on
`endif
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [1:0] io_tiles_cached_0_release_bits_client_xact_id,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_uncached_acquire_ready,
    input  io_htif_uncached_acquire_valid,
    input [25:0] io_htif_uncached_acquire_bits_addr_block,
    input [1:0] io_htif_uncached_acquire_bits_client_xact_id,
    input [1:0] io_htif_uncached_acquire_bits_addr_beat,
    input  io_htif_uncached_acquire_bits_is_builtin_type,
    input [2:0] io_htif_uncached_acquire_bits_a_type,
    input [16:0] io_htif_uncached_acquire_bits_union,
    input [127:0] io_htif_uncached_acquire_bits_data,
    input  io_htif_uncached_grant_ready,
    output io_htif_uncached_grant_valid,
    output[1:0] io_htif_uncached_grant_bits_addr_beat,
    output[1:0] io_htif_uncached_grant_bits_client_xact_id,
    output[2:0] io_htif_uncached_grant_bits_manager_xact_id,
    output io_htif_uncached_grant_bits_is_builtin_type,
    output[3:0] io_htif_uncached_grant_bits_g_type,
    output[127:0] io_htif_uncached_grant_bits_data,
    input  io_incoherent_0,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[3:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [3:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[3:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [3:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
    input  io_csr_0_req_ready,
    output io_csr_0_req_valid,
    output io_csr_0_req_bits_rw,
    output[11:0] io_csr_0_req_bits_addr,
    output[63:0] io_csr_0_req_bits_data,
    output io_csr_0_resp_ready,
    input  io_csr_0_resp_valid,
    input [63:0] io_csr_0_resp_bits,
    input  io_scr_req_ready,
    output io_scr_req_valid,
    output io_scr_req_bits_rw,
    output[5:0] io_scr_req_bits_addr,
    output[63:0] io_scr_req_bits_data,
    output io_scr_resp_ready,
    input  io_scr_resp_valid,
    input [63:0] io_scr_resp_bits,
    input  io_mmio_aw_ready,
    output io_mmio_aw_valid,
    output[31:0] io_mmio_aw_bits_addr,
    output[7:0] io_mmio_aw_bits_len,
    output[2:0] io_mmio_aw_bits_size,
    output[1:0] io_mmio_aw_bits_burst,
    output io_mmio_aw_bits_lock,
    output[3:0] io_mmio_aw_bits_cache,
    output[2:0] io_mmio_aw_bits_prot,
    output[3:0] io_mmio_aw_bits_qos,
    output[3:0] io_mmio_aw_bits_region,
    output[3:0] io_mmio_aw_bits_id,
    output io_mmio_aw_bits_user,
    input  io_mmio_w_ready,
    output io_mmio_w_valid,
    output[63:0] io_mmio_w_bits_data,
    output io_mmio_w_bits_last,
    output[7:0] io_mmio_w_bits_strb,
    output io_mmio_w_bits_user,
    output io_mmio_b_ready,
    input  io_mmio_b_valid,
    input [1:0] io_mmio_b_bits_resp,
    input [3:0] io_mmio_b_bits_id,
    input  io_mmio_b_bits_user,
    input  io_mmio_ar_ready,
    output io_mmio_ar_valid,
    output[31:0] io_mmio_ar_bits_addr,
    output[7:0] io_mmio_ar_bits_len,
    output[2:0] io_mmio_ar_bits_size,
    output[1:0] io_mmio_ar_bits_burst,
    output io_mmio_ar_bits_lock,
    output[3:0] io_mmio_ar_bits_cache,
    output[2:0] io_mmio_ar_bits_prot,
    output[3:0] io_mmio_ar_bits_qos,
    output[3:0] io_mmio_ar_bits_region,
    output[3:0] io_mmio_ar_bits_id,
    output io_mmio_ar_bits_user,
    output io_mmio_r_ready,
    input  io_mmio_r_valid,
    input [1:0] io_mmio_r_bits_resp,
    input [63:0] io_mmio_r_bits_data,
    input  io_mmio_r_bits_last,
    input [3:0] io_mmio_r_bits_id,
    input  io_mmio_r_bits_user,
    input  io_deviceTree_aw_ready,
    output io_deviceTree_aw_valid,
    output[31:0] io_deviceTree_aw_bits_addr,
    output[7:0] io_deviceTree_aw_bits_len,
    output[2:0] io_deviceTree_aw_bits_size,
    output[1:0] io_deviceTree_aw_bits_burst,
    output io_deviceTree_aw_bits_lock,
    output[3:0] io_deviceTree_aw_bits_cache,
    output[2:0] io_deviceTree_aw_bits_prot,
    output[3:0] io_deviceTree_aw_bits_qos,
    output[3:0] io_deviceTree_aw_bits_region,
    output[3:0] io_deviceTree_aw_bits_id,
    output io_deviceTree_aw_bits_user,
    input  io_deviceTree_w_ready,
    output io_deviceTree_w_valid,
    output[63:0] io_deviceTree_w_bits_data,
    output io_deviceTree_w_bits_last,
    output[7:0] io_deviceTree_w_bits_strb,
    output io_deviceTree_w_bits_user,
    output io_deviceTree_b_ready,
    input  io_deviceTree_b_valid,
    input [1:0] io_deviceTree_b_bits_resp,
    input [3:0] io_deviceTree_b_bits_id,
    input  io_deviceTree_b_bits_user,
    input  io_deviceTree_ar_ready,
    output io_deviceTree_ar_valid,
    output[31:0] io_deviceTree_ar_bits_addr,
    output[7:0] io_deviceTree_ar_bits_len,
    output[2:0] io_deviceTree_ar_bits_size,
    output[1:0] io_deviceTree_ar_bits_burst,
    output io_deviceTree_ar_bits_lock,
    output[3:0] io_deviceTree_ar_bits_cache,
    output[2:0] io_deviceTree_ar_bits_prot,
    output[3:0] io_deviceTree_ar_bits_qos,
    output[3:0] io_deviceTree_ar_bits_region,
    output[3:0] io_deviceTree_ar_bits_id,
    output io_deviceTree_ar_bits_user,
    output io_deviceTree_r_ready,
    input  io_deviceTree_r_valid,
    input [1:0] io_deviceTree_r_bits_resp,
    input [63:0] io_deviceTree_r_bits_data,
    input  io_deviceTree_r_bits_last,
    input [3:0] io_deviceTree_r_bits_id,
    input  io_deviceTree_r_bits_user
    //output io_dma_req_ready
    //input  io_dma_req_valid
    //input [1:0] io_dma_req_bits_client_xact_id
    //input [1:0] io_dma_req_bits_cmd
    //input [31:0] io_dma_req_bits_source
    //input [31:0] io_dma_req_bits_dest
    //input [31:0] io_dma_req_bits_length
    //input  io_dma_resp_ready
    //output io_dma_resp_valid
    //output[1:0] io_dma_resp_bits_client_xact_id
    //output[1:0] io_dma_resp_bits_status
);

  wire ClientTileLinkIOWrapper_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_io_out_release_valid;
  wire ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_1_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  wire[1:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  wire[2:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_1_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_1_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_1_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_1_io_out_release_valid;
  wire ClientTileLinkIOWrapper_2_io_in_acquire_ready;
  wire ClientTileLinkIOWrapper_2_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat;
  wire[2:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOWrapper_2_io_in_grant_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOWrapper_2_io_out_acquire_bits_data;
  wire ClientTileLinkIOWrapper_2_io_out_grant_ready;
  wire ClientTileLinkIOWrapper_2_io_out_probe_ready;
  wire ClientTileLinkIOWrapper_2_io_out_release_valid;
  wire ClientTileLinkEnqueuer_io_inner_acquire_ready;
  wire ClientTileLinkEnqueuer_io_inner_grant_valid;
  wire[1:0] ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat;
  wire[2:0] ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id;
  wire ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id;
  wire ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkEnqueuer_io_inner_grant_bits_g_type;
  wire[127:0] ClientTileLinkEnqueuer_io_inner_grant_bits_data;
  wire ClientTileLinkEnqueuer_io_inner_probe_valid;
  wire[25:0] ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block;
  wire[1:0] ClientTileLinkEnqueuer_io_inner_probe_bits_p_type;
  wire ClientTileLinkEnqueuer_io_inner_release_ready;
  wire ClientTileLinkEnqueuer_io_outer_acquire_valid;
  wire[25:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat;
  wire ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type;
  wire[16:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_union;
  wire[127:0] ClientTileLinkEnqueuer_io_outer_acquire_bits_data;
  wire ClientTileLinkEnqueuer_io_outer_grant_ready;
  wire ClientTileLinkEnqueuer_io_outer_probe_ready;
  wire ClientTileLinkEnqueuer_io_outer_release_valid;
  wire[1:0] ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat;
  wire[25:0] ClientTileLinkEnqueuer_io_outer_release_bits_addr_block;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id;
  wire ClientTileLinkEnqueuer_io_outer_release_bits_voluntary;
  wire[2:0] ClientTileLinkEnqueuer_io_outer_release_bits_r_type;
  wire[127:0] ClientTileLinkEnqueuer_io_outer_release_bits_data;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[31:0] Queue_io_deq_bits_addr;
  wire[7:0] Queue_io_deq_bits_len;
  wire[2:0] Queue_io_deq_bits_size;
  wire[1:0] Queue_io_deq_bits_burst;
  wire Queue_io_deq_bits_lock;
  wire[3:0] Queue_io_deq_bits_cache;
  wire[2:0] Queue_io_deq_bits_prot;
  wire[3:0] Queue_io_deq_bits_qos;
  wire[3:0] Queue_io_deq_bits_region;
  wire[3:0] Queue_io_deq_bits_id;
  wire Queue_io_deq_bits_user;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[31:0] Queue_1_io_deq_bits_addr;
  wire[7:0] Queue_1_io_deq_bits_len;
  wire[2:0] Queue_1_io_deq_bits_size;
  wire[1:0] Queue_1_io_deq_bits_burst;
  wire Queue_1_io_deq_bits_lock;
  wire[3:0] Queue_1_io_deq_bits_cache;
  wire[2:0] Queue_1_io_deq_bits_prot;
  wire[3:0] Queue_1_io_deq_bits_qos;
  wire[3:0] Queue_1_io_deq_bits_region;
  wire[3:0] Queue_1_io_deq_bits_id;
  wire Queue_1_io_deq_bits_user;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[63:0] Queue_2_io_deq_bits_data;
  wire Queue_2_io_deq_bits_last;
  wire[7:0] Queue_2_io_deq_bits_strb;
  wire Queue_2_io_deq_bits_user;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[1:0] Queue_3_io_deq_bits_resp;
  wire[63:0] Queue_3_io_deq_bits_data;
  wire Queue_3_io_deq_bits_last;
  wire[3:0] Queue_3_io_deq_bits_id;
  wire Queue_3_io_deq_bits_user;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[1:0] Queue_4_io_deq_bits_resp;
  wire[3:0] Queue_4_io_deq_bits_id;
  wire Queue_4_io_deq_bits_user;
  wire rtc_io_aw_valid;
  wire[31:0] rtc_io_aw_bits_addr;
  wire[7:0] rtc_io_aw_bits_len;
  wire[2:0] rtc_io_aw_bits_size;
  wire[1:0] rtc_io_aw_bits_burst;
  wire rtc_io_aw_bits_lock;
  wire[3:0] rtc_io_aw_bits_cache;
  wire[2:0] rtc_io_aw_bits_prot;
  wire[3:0] rtc_io_aw_bits_qos;
  wire[3:0] rtc_io_aw_bits_region;
  wire[3:0] rtc_io_aw_bits_id;
  wire rtc_io_aw_bits_user;
  wire rtc_io_w_valid;
  wire[63:0] rtc_io_w_bits_data;
  wire rtc_io_w_bits_last;
  wire[7:0] rtc_io_w_bits_strb;
  wire rtc_io_w_bits_user;
  wire rtc_io_b_ready;
  wire rtc_io_ar_valid;
  wire rtc_io_r_ready;
  wire ClientTileLinkIOUnwrapper_io_in_acquire_ready;
  wire ClientTileLinkIOUnwrapper_io_in_grant_valid;
  wire[1:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat;
  wire[2:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id;
  wire ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type;
  wire[3:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type;
  wire[127:0] ClientTileLinkIOUnwrapper_io_in_grant_bits_data;
  wire ClientTileLinkIOUnwrapper_io_in_probe_valid;
  wire ClientTileLinkIOUnwrapper_io_in_release_ready;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_valid;
  wire[25:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block;
  wire[2:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id;
  wire[1:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat;
  wire ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type;
  wire[2:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type;
  wire[16:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_union;
  wire[127:0] ClientTileLinkIOUnwrapper_io_out_acquire_bits_data;
  wire ClientTileLinkIOUnwrapper_io_out_grant_ready;
  wire TileLinkIONarrower_io_in_acquire_ready;
  wire TileLinkIONarrower_io_in_grant_valid;
  wire[1:0] TileLinkIONarrower_io_in_grant_bits_addr_beat;
  wire[2:0] TileLinkIONarrower_io_in_grant_bits_client_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_manager_xact_id;
  wire TileLinkIONarrower_io_in_grant_bits_is_builtin_type;
  wire[3:0] TileLinkIONarrower_io_in_grant_bits_g_type;
  wire[127:0] TileLinkIONarrower_io_in_grant_bits_data;
  wire TileLinkIONarrower_io_out_acquire_valid;
  wire[25:0] TileLinkIONarrower_io_out_acquire_bits_addr_block;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_client_xact_id;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_addr_beat;
  wire TileLinkIONarrower_io_out_acquire_bits_is_builtin_type;
  wire[2:0] TileLinkIONarrower_io_out_acquire_bits_a_type;
  wire[11:0] TileLinkIONarrower_io_out_acquire_bits_union;
  wire[63:0] TileLinkIONarrower_io_out_acquire_bits_data;
  wire TileLinkIONarrower_io_out_grant_ready;
  wire NastiIOTileLinkIOConverter_io_tl_acquire_ready;
  wire NastiIOTileLinkIOConverter_io_tl_grant_valid;
  wire[2:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat;
  wire[2:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id;
  wire NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type;
  wire[3:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type;
  wire[63:0] NastiIOTileLinkIOConverter_io_tl_grant_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_region;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_aw_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_aw_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_w_valid;
  wire[63:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_data;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_last;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_w_bits_strb;
  wire NastiIOTileLinkIOConverter_io_nasti_w_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_b_ready;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_valid;
  wire[31:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr;
  wire[7:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_len;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_size;
  wire[1:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache;
  wire[2:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_region;
  wire[3:0] NastiIOTileLinkIOConverter_io_nasti_ar_bits_id;
  wire NastiIOTileLinkIOConverter_io_nasti_ar_bits_user;
  wire NastiIOTileLinkIOConverter_io_nasti_r_ready;
  wire L2BroadcastHub_io_inner_acquire_ready;
  wire L2BroadcastHub_io_inner_grant_valid;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_addr_beat;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_xact_id;
  wire[2:0] L2BroadcastHub_io_inner_grant_bits_manager_xact_id;
  wire L2BroadcastHub_io_inner_grant_bits_is_builtin_type;
  wire[3:0] L2BroadcastHub_io_inner_grant_bits_g_type;
  wire[127:0] L2BroadcastHub_io_inner_grant_bits_data;
  wire[1:0] L2BroadcastHub_io_inner_grant_bits_client_id;
  wire L2BroadcastHub_io_inner_finish_ready;
  wire L2BroadcastHub_io_inner_probe_valid;
  wire[25:0] L2BroadcastHub_io_inner_probe_bits_addr_block;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_p_type;
  wire[1:0] L2BroadcastHub_io_inner_probe_bits_client_id;
  wire L2BroadcastHub_io_inner_release_ready;
  wire L2BroadcastHub_io_outer_acquire_valid;
  wire[25:0] L2BroadcastHub_io_outer_acquire_bits_addr_block;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_client_xact_id;
  wire[1:0] L2BroadcastHub_io_outer_acquire_bits_addr_beat;
  wire L2BroadcastHub_io_outer_acquire_bits_is_builtin_type;
  wire[2:0] L2BroadcastHub_io_outer_acquire_bits_a_type;
  wire[16:0] L2BroadcastHub_io_outer_acquire_bits_union;
  wire[127:0] L2BroadcastHub_io_outer_acquire_bits_data;
  wire L2BroadcastHub_io_outer_grant_ready;
  wire SMIIONastiIOConverter_io_nasti_aw_ready;
  wire SMIIONastiIOConverter_io_nasti_w_ready;
  wire SMIIONastiIOConverter_io_nasti_b_valid;
  wire[1:0] SMIIONastiIOConverter_io_nasti_b_bits_resp;
  wire[3:0] SMIIONastiIOConverter_io_nasti_b_bits_id;
  wire SMIIONastiIOConverter_io_nasti_b_bits_user;
  wire SMIIONastiIOConverter_io_nasti_ar_ready;
  wire SMIIONastiIOConverter_io_nasti_r_valid;
  wire[1:0] SMIIONastiIOConverter_io_nasti_r_bits_resp;
  wire[63:0] SMIIONastiIOConverter_io_nasti_r_bits_data;
  wire SMIIONastiIOConverter_io_nasti_r_bits_last;
  wire[3:0] SMIIONastiIOConverter_io_nasti_r_bits_id;
  wire SMIIONastiIOConverter_io_nasti_r_bits_user;
  wire SMIIONastiIOConverter_io_smi_req_valid;
  wire SMIIONastiIOConverter_io_smi_req_bits_rw;
  wire[11:0] SMIIONastiIOConverter_io_smi_req_bits_addr;
  wire[63:0] SMIIONastiIOConverter_io_smi_req_bits_data;
  wire SMIIONastiIOConverter_io_smi_resp_ready;
  wire conv_io_nasti_aw_ready;
  wire conv_io_nasti_w_ready;
  wire conv_io_nasti_b_valid;
  wire[1:0] conv_io_nasti_b_bits_resp;
  wire[3:0] conv_io_nasti_b_bits_id;
  wire conv_io_nasti_b_bits_user;
  wire conv_io_nasti_ar_ready;
  wire conv_io_nasti_r_valid;
  wire[1:0] conv_io_nasti_r_bits_resp;
  wire[63:0] conv_io_nasti_r_bits_data;
  wire conv_io_nasti_r_bits_last;
  wire[3:0] conv_io_nasti_r_bits_id;
  wire conv_io_nasti_r_bits_user;
  wire conv_io_smi_req_valid;
  wire conv_io_smi_req_bits_rw;
  wire[5:0] conv_io_smi_req_bits_addr;
  wire[63:0] conv_io_smi_req_bits_data;
  wire conv_io_smi_resp_ready;
  wire l1tol2net_io_clients_2_acquire_ready;
  wire l1tol2net_io_clients_2_grant_valid;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_2_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_2_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_2_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_2_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_2_grant_bits_data;
  wire l1tol2net_io_clients_2_probe_valid;
  wire[25:0] l1tol2net_io_clients_2_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_2_probe_bits_p_type;
  wire l1tol2net_io_clients_2_release_ready;
  wire l1tol2net_io_clients_1_acquire_ready;
  wire l1tol2net_io_clients_1_grant_valid;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_1_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_1_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_1_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_1_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_1_grant_bits_data;
  wire l1tol2net_io_clients_1_probe_valid;
  wire[25:0] l1tol2net_io_clients_1_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_1_probe_bits_p_type;
  wire l1tol2net_io_clients_1_release_ready;
  wire l1tol2net_io_clients_0_acquire_ready;
  wire l1tol2net_io_clients_0_grant_valid;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_addr_beat;
  wire[1:0] l1tol2net_io_clients_0_grant_bits_client_xact_id;
  wire[2:0] l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  wire l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  wire[3:0] l1tol2net_io_clients_0_grant_bits_g_type;
  wire[127:0] l1tol2net_io_clients_0_grant_bits_data;
  wire l1tol2net_io_clients_0_probe_valid;
  wire[25:0] l1tol2net_io_clients_0_probe_bits_addr_block;
  wire[1:0] l1tol2net_io_clients_0_probe_bits_p_type;
  wire l1tol2net_io_clients_0_release_ready;
  wire l1tol2net_io_managers_0_acquire_valid;
  wire[25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire[2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire[16:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire[127:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire[1:0] l1tol2net_io_managers_0_acquire_bits_client_id;
  wire l1tol2net_io_managers_0_grant_ready;
  wire l1tol2net_io_managers_0_finish_valid;
  wire[2:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire l1tol2net_io_managers_0_probe_ready;
  wire l1tol2net_io_managers_0_release_valid;
  wire[1:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire[25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire l1tol2net_io_managers_0_release_bits_voluntary;
  wire[2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire[127:0] l1tol2net_io_managers_0_release_bits_data;
  wire[1:0] l1tol2net_io_managers_0_release_bits_client_id;
  wire interconnect_io_masters_1_aw_ready;
  wire interconnect_io_masters_1_w_ready;
  wire interconnect_io_masters_1_b_valid;
  wire[1:0] interconnect_io_masters_1_b_bits_resp;
  wire[3:0] interconnect_io_masters_1_b_bits_id;
  wire interconnect_io_masters_1_b_bits_user;
  wire interconnect_io_masters_1_ar_ready;
  wire interconnect_io_masters_1_r_valid;
  wire[1:0] interconnect_io_masters_1_r_bits_resp;
  wire[63:0] interconnect_io_masters_1_r_bits_data;
  wire interconnect_io_masters_1_r_bits_last;
  wire[3:0] interconnect_io_masters_1_r_bits_id;
  wire interconnect_io_masters_1_r_bits_user;
  wire interconnect_io_masters_0_aw_ready;
  wire interconnect_io_masters_0_w_ready;
  wire interconnect_io_masters_0_b_valid;
  wire[1:0] interconnect_io_masters_0_b_bits_resp;
  wire[3:0] interconnect_io_masters_0_b_bits_id;
  wire interconnect_io_masters_0_b_bits_user;
  wire interconnect_io_masters_0_ar_ready;
  wire interconnect_io_masters_0_r_valid;
  wire[1:0] interconnect_io_masters_0_r_bits_resp;
  wire[63:0] interconnect_io_masters_0_r_bits_data;
  wire interconnect_io_masters_0_r_bits_last;
  wire[3:0] interconnect_io_masters_0_r_bits_id;
  wire interconnect_io_masters_0_r_bits_user;
  wire interconnect_io_slaves_4_aw_valid;
  wire[31:0] interconnect_io_slaves_4_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_4_aw_bits_len;
  wire[2:0] interconnect_io_slaves_4_aw_bits_size;
  wire[1:0] interconnect_io_slaves_4_aw_bits_burst;
  wire interconnect_io_slaves_4_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_4_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_4_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_4_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_4_aw_bits_region;
  wire[3:0] interconnect_io_slaves_4_aw_bits_id;
  wire interconnect_io_slaves_4_aw_bits_user;
  wire interconnect_io_slaves_4_w_valid;
  wire[63:0] interconnect_io_slaves_4_w_bits_data;
  wire interconnect_io_slaves_4_w_bits_last;
  wire[7:0] interconnect_io_slaves_4_w_bits_strb;
  wire interconnect_io_slaves_4_w_bits_user;
  wire interconnect_io_slaves_4_b_ready;
  wire interconnect_io_slaves_4_ar_valid;
  wire[31:0] interconnect_io_slaves_4_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_4_ar_bits_len;
  wire[2:0] interconnect_io_slaves_4_ar_bits_size;
  wire[1:0] interconnect_io_slaves_4_ar_bits_burst;
  wire interconnect_io_slaves_4_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_4_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_4_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_4_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_4_ar_bits_region;
  wire[3:0] interconnect_io_slaves_4_ar_bits_id;
  wire interconnect_io_slaves_4_ar_bits_user;
  wire interconnect_io_slaves_4_r_ready;
  wire interconnect_io_slaves_3_aw_valid;
  wire[31:0] interconnect_io_slaves_3_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_3_aw_bits_len;
  wire[2:0] interconnect_io_slaves_3_aw_bits_size;
  wire[1:0] interconnect_io_slaves_3_aw_bits_burst;
  wire interconnect_io_slaves_3_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_3_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_3_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_3_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_3_aw_bits_region;
  wire[3:0] interconnect_io_slaves_3_aw_bits_id;
  wire interconnect_io_slaves_3_aw_bits_user;
  wire interconnect_io_slaves_3_w_valid;
  wire[63:0] interconnect_io_slaves_3_w_bits_data;
  wire interconnect_io_slaves_3_w_bits_last;
  wire[7:0] interconnect_io_slaves_3_w_bits_strb;
  wire interconnect_io_slaves_3_w_bits_user;
  wire interconnect_io_slaves_3_b_ready;
  wire interconnect_io_slaves_3_ar_valid;
  wire[31:0] interconnect_io_slaves_3_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_3_ar_bits_len;
  wire[2:0] interconnect_io_slaves_3_ar_bits_size;
  wire[1:0] interconnect_io_slaves_3_ar_bits_burst;
  wire interconnect_io_slaves_3_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_3_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_3_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_3_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_3_ar_bits_region;
  wire[3:0] interconnect_io_slaves_3_ar_bits_id;
  wire interconnect_io_slaves_3_ar_bits_user;
  wire interconnect_io_slaves_3_r_ready;
  wire interconnect_io_slaves_2_aw_valid;
  wire[31:0] interconnect_io_slaves_2_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_2_aw_bits_len;
  wire[2:0] interconnect_io_slaves_2_aw_bits_size;
  wire[1:0] interconnect_io_slaves_2_aw_bits_burst;
  wire interconnect_io_slaves_2_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_2_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_2_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_2_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_2_aw_bits_region;
  wire[3:0] interconnect_io_slaves_2_aw_bits_id;
  wire interconnect_io_slaves_2_aw_bits_user;
  wire interconnect_io_slaves_2_w_valid;
  wire[63:0] interconnect_io_slaves_2_w_bits_data;
  wire interconnect_io_slaves_2_w_bits_last;
  wire[7:0] interconnect_io_slaves_2_w_bits_strb;
  wire interconnect_io_slaves_2_w_bits_user;
  wire interconnect_io_slaves_2_b_ready;
  wire interconnect_io_slaves_2_ar_valid;
  wire[31:0] interconnect_io_slaves_2_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_2_ar_bits_len;
  wire[2:0] interconnect_io_slaves_2_ar_bits_size;
  wire[1:0] interconnect_io_slaves_2_ar_bits_burst;
  wire interconnect_io_slaves_2_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_2_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_2_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_2_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_2_ar_bits_region;
  wire[3:0] interconnect_io_slaves_2_ar_bits_id;
  wire interconnect_io_slaves_2_ar_bits_user;
  wire interconnect_io_slaves_2_r_ready;
  wire interconnect_io_slaves_1_aw_valid;
  wire[31:0] interconnect_io_slaves_1_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_1_aw_bits_len;
  wire[2:0] interconnect_io_slaves_1_aw_bits_size;
  wire[1:0] interconnect_io_slaves_1_aw_bits_burst;
  wire interconnect_io_slaves_1_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_1_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_1_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_1_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_1_aw_bits_region;
  wire[3:0] interconnect_io_slaves_1_aw_bits_id;
  wire interconnect_io_slaves_1_aw_bits_user;
  wire interconnect_io_slaves_1_w_valid;
  wire[63:0] interconnect_io_slaves_1_w_bits_data;
  wire interconnect_io_slaves_1_w_bits_last;
  wire[7:0] interconnect_io_slaves_1_w_bits_strb;
  wire interconnect_io_slaves_1_w_bits_user;
  wire interconnect_io_slaves_1_b_ready;
  wire interconnect_io_slaves_1_ar_valid;
  wire[31:0] interconnect_io_slaves_1_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_1_ar_bits_len;
  wire[2:0] interconnect_io_slaves_1_ar_bits_size;
  wire[1:0] interconnect_io_slaves_1_ar_bits_burst;
  wire interconnect_io_slaves_1_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_1_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_1_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_1_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_1_ar_bits_region;
  wire[3:0] interconnect_io_slaves_1_ar_bits_id;
  wire interconnect_io_slaves_1_ar_bits_user;
  wire interconnect_io_slaves_1_r_ready;
  wire interconnect_io_slaves_0_aw_valid;
  wire[31:0] interconnect_io_slaves_0_aw_bits_addr;
  wire[7:0] interconnect_io_slaves_0_aw_bits_len;
  wire[2:0] interconnect_io_slaves_0_aw_bits_size;
  wire[1:0] interconnect_io_slaves_0_aw_bits_burst;
  wire interconnect_io_slaves_0_aw_bits_lock;
  wire[3:0] interconnect_io_slaves_0_aw_bits_cache;
  wire[2:0] interconnect_io_slaves_0_aw_bits_prot;
  wire[3:0] interconnect_io_slaves_0_aw_bits_qos;
  wire[3:0] interconnect_io_slaves_0_aw_bits_region;
  wire[3:0] interconnect_io_slaves_0_aw_bits_id;
  wire interconnect_io_slaves_0_aw_bits_user;
  wire interconnect_io_slaves_0_w_valid;
  wire[63:0] interconnect_io_slaves_0_w_bits_data;
  wire interconnect_io_slaves_0_w_bits_last;
  wire[7:0] interconnect_io_slaves_0_w_bits_strb;
  wire interconnect_io_slaves_0_w_bits_user;
  wire interconnect_io_slaves_0_b_ready;
  wire interconnect_io_slaves_0_ar_valid;
  wire[31:0] interconnect_io_slaves_0_ar_bits_addr;
  wire[7:0] interconnect_io_slaves_0_ar_bits_len;
  wire[2:0] interconnect_io_slaves_0_ar_bits_size;
  wire[1:0] interconnect_io_slaves_0_ar_bits_burst;
  wire interconnect_io_slaves_0_ar_bits_lock;
  wire[3:0] interconnect_io_slaves_0_ar_bits_cache;
  wire[2:0] interconnect_io_slaves_0_ar_bits_prot;
  wire[3:0] interconnect_io_slaves_0_ar_bits_qos;
  wire[3:0] interconnect_io_slaves_0_ar_bits_region;
  wire[3:0] interconnect_io_slaves_0_ar_bits_id;
  wire interconnect_io_slaves_0_ar_bits_user;
  wire interconnect_io_slaves_0_r_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_dma_resp_bits_status = {1{$random}};
//  assign io_dma_resp_bits_client_xact_id = {1{$random}};
//  assign io_dma_resp_valid = {1{$random}};
//  assign io_dma_req_ready = {1{$random}};
//  assign io_mem_backup_req_bits = {1{$random}};
//  assign io_mem_backup_req_valid = {1{$random}};
// synthesis translate_on
`endif
  assign io_deviceTree_r_ready = interconnect_io_slaves_1_r_ready;
  assign io_deviceTree_ar_bits_user = interconnect_io_slaves_1_ar_bits_user;
  assign io_deviceTree_ar_bits_id = interconnect_io_slaves_1_ar_bits_id;
  assign io_deviceTree_ar_bits_region = interconnect_io_slaves_1_ar_bits_region;
  assign io_deviceTree_ar_bits_qos = interconnect_io_slaves_1_ar_bits_qos;
  assign io_deviceTree_ar_bits_prot = interconnect_io_slaves_1_ar_bits_prot;
  assign io_deviceTree_ar_bits_cache = interconnect_io_slaves_1_ar_bits_cache;
  assign io_deviceTree_ar_bits_lock = interconnect_io_slaves_1_ar_bits_lock;
  assign io_deviceTree_ar_bits_burst = interconnect_io_slaves_1_ar_bits_burst;
  assign io_deviceTree_ar_bits_size = interconnect_io_slaves_1_ar_bits_size;
  assign io_deviceTree_ar_bits_len = interconnect_io_slaves_1_ar_bits_len;
  assign io_deviceTree_ar_bits_addr = interconnect_io_slaves_1_ar_bits_addr;
  assign io_deviceTree_ar_valid = interconnect_io_slaves_1_ar_valid;
  assign io_deviceTree_b_ready = interconnect_io_slaves_1_b_ready;
  assign io_deviceTree_w_bits_user = interconnect_io_slaves_1_w_bits_user;
  assign io_deviceTree_w_bits_strb = interconnect_io_slaves_1_w_bits_strb;
  assign io_deviceTree_w_bits_last = interconnect_io_slaves_1_w_bits_last;
  assign io_deviceTree_w_bits_data = interconnect_io_slaves_1_w_bits_data;
  assign io_deviceTree_w_valid = interconnect_io_slaves_1_w_valid;
  assign io_deviceTree_aw_bits_user = interconnect_io_slaves_1_aw_bits_user;
  assign io_deviceTree_aw_bits_id = interconnect_io_slaves_1_aw_bits_id;
  assign io_deviceTree_aw_bits_region = interconnect_io_slaves_1_aw_bits_region;
  assign io_deviceTree_aw_bits_qos = interconnect_io_slaves_1_aw_bits_qos;
  assign io_deviceTree_aw_bits_prot = interconnect_io_slaves_1_aw_bits_prot;
  assign io_deviceTree_aw_bits_cache = interconnect_io_slaves_1_aw_bits_cache;
  assign io_deviceTree_aw_bits_lock = interconnect_io_slaves_1_aw_bits_lock;
  assign io_deviceTree_aw_bits_burst = interconnect_io_slaves_1_aw_bits_burst;
  assign io_deviceTree_aw_bits_size = interconnect_io_slaves_1_aw_bits_size;
  assign io_deviceTree_aw_bits_len = interconnect_io_slaves_1_aw_bits_len;
  assign io_deviceTree_aw_bits_addr = interconnect_io_slaves_1_aw_bits_addr;
  assign io_deviceTree_aw_valid = interconnect_io_slaves_1_aw_valid;
  assign io_mmio_r_ready = interconnect_io_slaves_4_r_ready;
  assign io_mmio_ar_bits_user = interconnect_io_slaves_4_ar_bits_user;
  assign io_mmio_ar_bits_id = interconnect_io_slaves_4_ar_bits_id;
  assign io_mmio_ar_bits_region = interconnect_io_slaves_4_ar_bits_region;
  assign io_mmio_ar_bits_qos = interconnect_io_slaves_4_ar_bits_qos;
  assign io_mmio_ar_bits_prot = interconnect_io_slaves_4_ar_bits_prot;
  assign io_mmio_ar_bits_cache = interconnect_io_slaves_4_ar_bits_cache;
  assign io_mmio_ar_bits_lock = interconnect_io_slaves_4_ar_bits_lock;
  assign io_mmio_ar_bits_burst = interconnect_io_slaves_4_ar_bits_burst;
  assign io_mmio_ar_bits_size = interconnect_io_slaves_4_ar_bits_size;
  assign io_mmio_ar_bits_len = interconnect_io_slaves_4_ar_bits_len;
  assign io_mmio_ar_bits_addr = interconnect_io_slaves_4_ar_bits_addr;
  assign io_mmio_ar_valid = interconnect_io_slaves_4_ar_valid;
  assign io_mmio_b_ready = interconnect_io_slaves_4_b_ready;
  assign io_mmio_w_bits_user = interconnect_io_slaves_4_w_bits_user;
  assign io_mmio_w_bits_strb = interconnect_io_slaves_4_w_bits_strb;
  assign io_mmio_w_bits_last = interconnect_io_slaves_4_w_bits_last;
  assign io_mmio_w_bits_data = interconnect_io_slaves_4_w_bits_data;
  assign io_mmio_w_valid = interconnect_io_slaves_4_w_valid;
  assign io_mmio_aw_bits_user = interconnect_io_slaves_4_aw_bits_user;
  assign io_mmio_aw_bits_id = interconnect_io_slaves_4_aw_bits_id;
  assign io_mmio_aw_bits_region = interconnect_io_slaves_4_aw_bits_region;
  assign io_mmio_aw_bits_qos = interconnect_io_slaves_4_aw_bits_qos;
  assign io_mmio_aw_bits_prot = interconnect_io_slaves_4_aw_bits_prot;
  assign io_mmio_aw_bits_cache = interconnect_io_slaves_4_aw_bits_cache;
  assign io_mmio_aw_bits_lock = interconnect_io_slaves_4_aw_bits_lock;
  assign io_mmio_aw_bits_burst = interconnect_io_slaves_4_aw_bits_burst;
  assign io_mmio_aw_bits_size = interconnect_io_slaves_4_aw_bits_size;
  assign io_mmio_aw_bits_len = interconnect_io_slaves_4_aw_bits_len;
  assign io_mmio_aw_bits_addr = interconnect_io_slaves_4_aw_bits_addr;
  assign io_mmio_aw_valid = interconnect_io_slaves_4_aw_valid;
  assign io_scr_resp_ready = conv_io_smi_resp_ready;
  assign io_scr_req_bits_data = conv_io_smi_req_bits_data;
  assign io_scr_req_bits_addr = conv_io_smi_req_bits_addr;
  assign io_scr_req_bits_rw = conv_io_smi_req_bits_rw;
  assign io_scr_req_valid = conv_io_smi_req_valid;
  assign io_csr_0_resp_ready = SMIIONastiIOConverter_io_smi_resp_ready;
  assign io_csr_0_req_bits_data = SMIIONastiIOConverter_io_smi_req_bits_data;
  assign io_csr_0_req_bits_addr = SMIIONastiIOConverter_io_smi_req_bits_addr;
  assign io_csr_0_req_bits_rw = SMIIONastiIOConverter_io_smi_req_bits_rw;
  assign io_csr_0_req_valid = SMIIONastiIOConverter_io_smi_req_valid;
  assign io_mem_0_r_ready = interconnect_io_slaves_0_r_ready;
  assign io_mem_0_ar_bits_user = interconnect_io_slaves_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = interconnect_io_slaves_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = interconnect_io_slaves_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = interconnect_io_slaves_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = interconnect_io_slaves_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = interconnect_io_slaves_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = interconnect_io_slaves_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = interconnect_io_slaves_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = interconnect_io_slaves_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = interconnect_io_slaves_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = interconnect_io_slaves_0_ar_bits_addr;
  assign io_mem_0_ar_valid = interconnect_io_slaves_0_ar_valid;
  assign io_mem_0_b_ready = interconnect_io_slaves_0_b_ready;
  assign io_mem_0_w_bits_user = interconnect_io_slaves_0_w_bits_user;
  assign io_mem_0_w_bits_strb = interconnect_io_slaves_0_w_bits_strb;
  assign io_mem_0_w_bits_last = interconnect_io_slaves_0_w_bits_last;
  assign io_mem_0_w_bits_data = interconnect_io_slaves_0_w_bits_data;
  assign io_mem_0_w_valid = interconnect_io_slaves_0_w_valid;
  assign io_mem_0_aw_bits_user = interconnect_io_slaves_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = interconnect_io_slaves_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = interconnect_io_slaves_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = interconnect_io_slaves_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = interconnect_io_slaves_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = interconnect_io_slaves_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = interconnect_io_slaves_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = interconnect_io_slaves_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = interconnect_io_slaves_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = interconnect_io_slaves_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = interconnect_io_slaves_0_aw_bits_addr;
  assign io_mem_0_aw_valid = interconnect_io_slaves_0_aw_valid;
  assign io_htif_uncached_grant_bits_data = ClientTileLinkIOWrapper_1_io_in_grant_bits_data;
  assign io_htif_uncached_grant_bits_g_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type;
  assign io_htif_uncached_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type;
  assign io_htif_uncached_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id;
  assign io_htif_uncached_grant_bits_client_xact_id = ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id;
  assign io_htif_uncached_grant_bits_addr_beat = ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat;
  assign io_htif_uncached_grant_valid = ClientTileLinkIOWrapper_1_io_in_grant_valid;
  assign io_htif_uncached_acquire_ready = ClientTileLinkIOWrapper_1_io_in_acquire_ready;
  assign io_tiles_uncached_0_grant_bits_data = ClientTileLinkIOWrapper_io_in_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = ClientTileLinkIOWrapper_io_in_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = ClientTileLinkIOWrapper_io_in_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = ClientTileLinkIOWrapper_io_in_acquire_ready;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_0_acquire_ready;
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_in_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_in_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  ClientTileLinkIOWrapper_0 ClientTileLinkIOWrapper_1(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_1_io_in_acquire_ready ),
       .io_in_acquire_valid( io_htif_uncached_acquire_valid ),
       .io_in_acquire_bits_addr_block( io_htif_uncached_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( io_htif_uncached_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( io_htif_uncached_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( io_htif_uncached_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( io_htif_uncached_acquire_bits_a_type ),
       .io_in_acquire_bits_union( io_htif_uncached_acquire_bits_union ),
       .io_in_acquire_bits_data( io_htif_uncached_acquire_bits_data ),
       .io_in_grant_ready( io_htif_uncached_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_1_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_1_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_1_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_1_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_1_io_in_grant_bits_data ),
       .io_out_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_out_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_out_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_out_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_out_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_out_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_out_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  RocketChipTileLinkArbiter l1tol2net(.clk(clk), .reset(reset),
       .io_clients_2_acquire_ready( l1tol2net_io_clients_2_acquire_ready ),
       .io_clients_2_acquire_valid( ClientTileLinkIOWrapper_1_io_out_acquire_valid ),
       .io_clients_2_acquire_bits_addr_block( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_block ),
       .io_clients_2_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_1_io_out_acquire_bits_client_xact_id ),
       .io_clients_2_acquire_bits_addr_beat( ClientTileLinkIOWrapper_1_io_out_acquire_bits_addr_beat ),
       .io_clients_2_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_is_builtin_type ),
       .io_clients_2_acquire_bits_a_type( ClientTileLinkIOWrapper_1_io_out_acquire_bits_a_type ),
       .io_clients_2_acquire_bits_union( ClientTileLinkIOWrapper_1_io_out_acquire_bits_union ),
       .io_clients_2_acquire_bits_data( ClientTileLinkIOWrapper_1_io_out_acquire_bits_data ),
       .io_clients_2_grant_ready( ClientTileLinkIOWrapper_1_io_out_grant_ready ),
       .io_clients_2_grant_valid( l1tol2net_io_clients_2_grant_valid ),
       .io_clients_2_grant_bits_addr_beat( l1tol2net_io_clients_2_grant_bits_addr_beat ),
       .io_clients_2_grant_bits_client_xact_id( l1tol2net_io_clients_2_grant_bits_client_xact_id ),
       .io_clients_2_grant_bits_manager_xact_id( l1tol2net_io_clients_2_grant_bits_manager_xact_id ),
       .io_clients_2_grant_bits_is_builtin_type( l1tol2net_io_clients_2_grant_bits_is_builtin_type ),
       .io_clients_2_grant_bits_g_type( l1tol2net_io_clients_2_grant_bits_g_type ),
       .io_clients_2_grant_bits_data( l1tol2net_io_clients_2_grant_bits_data ),
       .io_clients_2_probe_ready( ClientTileLinkIOWrapper_1_io_out_probe_ready ),
       .io_clients_2_probe_valid( l1tol2net_io_clients_2_probe_valid ),
       .io_clients_2_probe_bits_addr_block( l1tol2net_io_clients_2_probe_bits_addr_block ),
       .io_clients_2_probe_bits_p_type( l1tol2net_io_clients_2_probe_bits_p_type ),
       .io_clients_2_release_ready( l1tol2net_io_clients_2_release_ready ),
       .io_clients_2_release_valid( ClientTileLinkIOWrapper_1_io_out_release_valid ),
       //.io_clients_2_release_bits_addr_beat(  )
       //.io_clients_2_release_bits_addr_block(  )
       //.io_clients_2_release_bits_client_xact_id(  )
       //.io_clients_2_release_bits_voluntary(  )
       //.io_clients_2_release_bits_r_type(  )
       //.io_clients_2_release_bits_data(  )
       .io_clients_1_acquire_ready( l1tol2net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( ClientTileLinkIOWrapper_io_out_acquire_valid ),
       .io_clients_1_acquire_bits_addr_block( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_block ),
       .io_clients_1_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_io_out_acquire_bits_client_xact_id ),
       .io_clients_1_acquire_bits_addr_beat( ClientTileLinkIOWrapper_io_out_acquire_bits_addr_beat ),
       .io_clients_1_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_io_out_acquire_bits_is_builtin_type ),
       .io_clients_1_acquire_bits_a_type( ClientTileLinkIOWrapper_io_out_acquire_bits_a_type ),
       .io_clients_1_acquire_bits_union( ClientTileLinkIOWrapper_io_out_acquire_bits_union ),
       .io_clients_1_acquire_bits_data( ClientTileLinkIOWrapper_io_out_acquire_bits_data ),
       .io_clients_1_grant_ready( ClientTileLinkIOWrapper_io_out_grant_ready ),
       .io_clients_1_grant_valid( l1tol2net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_addr_beat( l1tol2net_io_clients_1_grant_bits_addr_beat ),
       .io_clients_1_grant_bits_client_xact_id( l1tol2net_io_clients_1_grant_bits_client_xact_id ),
       .io_clients_1_grant_bits_manager_xact_id( l1tol2net_io_clients_1_grant_bits_manager_xact_id ),
       .io_clients_1_grant_bits_is_builtin_type( l1tol2net_io_clients_1_grant_bits_is_builtin_type ),
       .io_clients_1_grant_bits_g_type( l1tol2net_io_clients_1_grant_bits_g_type ),
       .io_clients_1_grant_bits_data( l1tol2net_io_clients_1_grant_bits_data ),
       .io_clients_1_probe_ready( ClientTileLinkIOWrapper_io_out_probe_ready ),
       .io_clients_1_probe_valid( l1tol2net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_addr_block( l1tol2net_io_clients_1_probe_bits_addr_block ),
       .io_clients_1_probe_bits_p_type( l1tol2net_io_clients_1_probe_bits_p_type ),
       .io_clients_1_release_ready( l1tol2net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( ClientTileLinkIOWrapper_io_out_release_valid ),
       //.io_clients_1_release_bits_addr_beat(  )
       //.io_clients_1_release_bits_addr_block(  )
       //.io_clients_1_release_bits_client_xact_id(  )
       //.io_clients_1_release_bits_voluntary(  )
       //.io_clients_1_release_bits_r_type(  )
       //.io_clients_1_release_bits_data(  )
       .io_clients_0_acquire_ready( l1tol2net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_clients_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_clients_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_clients_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_clients_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_clients_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_clients_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_clients_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_clients_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_clients_0_grant_valid( l1tol2net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_addr_beat( l1tol2net_io_clients_0_grant_bits_addr_beat ),
       .io_clients_0_grant_bits_client_xact_id( l1tol2net_io_clients_0_grant_bits_client_xact_id ),
       .io_clients_0_grant_bits_manager_xact_id( l1tol2net_io_clients_0_grant_bits_manager_xact_id ),
       .io_clients_0_grant_bits_is_builtin_type( l1tol2net_io_clients_0_grant_bits_is_builtin_type ),
       .io_clients_0_grant_bits_g_type( l1tol2net_io_clients_0_grant_bits_g_type ),
       .io_clients_0_grant_bits_data( l1tol2net_io_clients_0_grant_bits_data ),
       .io_clients_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_clients_0_probe_valid( l1tol2net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_addr_block( l1tol2net_io_clients_0_probe_bits_addr_block ),
       .io_clients_0_probe_bits_p_type( l1tol2net_io_clients_0_probe_bits_p_type ),
       .io_clients_0_release_ready( l1tol2net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_clients_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_clients_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_clients_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_clients_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_clients_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_clients_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_managers_0_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_managers_0_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_managers_0_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_managers_0_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_managers_0_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_managers_0_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_managers_0_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_managers_0_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_managers_0_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_managers_0_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_managers_0_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_managers_0_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_managers_0_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_managers_0_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_managers_0_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_managers_0_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_managers_0_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_managers_0_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_managers_0_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_managers_0_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_managers_0_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_managers_0_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_managers_0_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_managers_0_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_managers_0_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_managers_0_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_managers_0_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_managers_0_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_managers_0_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_managers_0_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_managers_0_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_managers_0_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_managers_0_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_managers_0_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_managers_0_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_managers_0_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign l1tol2net.io_clients_2_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_2_release_bits_data = {4{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_beat = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_addr_block = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_client_xact_id = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_voluntary = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_r_type = {1{$random}};
    assign l1tol2net.io_clients_1_release_bits_data = {4{$random}};
// synthesis translate_on
`endif
  L2BroadcastHub L2BroadcastHub(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2BroadcastHub_io_inner_acquire_ready ),
       .io_inner_acquire_valid( l1tol2net_io_managers_0_acquire_valid ),
       .io_inner_acquire_bits_addr_block( l1tol2net_io_managers_0_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( l1tol2net_io_managers_0_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( l1tol2net_io_managers_0_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( l1tol2net_io_managers_0_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( l1tol2net_io_managers_0_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( l1tol2net_io_managers_0_acquire_bits_union ),
       .io_inner_acquire_bits_data( l1tol2net_io_managers_0_acquire_bits_data ),
       .io_inner_acquire_bits_client_id( l1tol2net_io_managers_0_acquire_bits_client_id ),
       .io_inner_grant_ready( l1tol2net_io_managers_0_grant_ready ),
       .io_inner_grant_valid( L2BroadcastHub_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( L2BroadcastHub_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( L2BroadcastHub_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( L2BroadcastHub_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( L2BroadcastHub_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( L2BroadcastHub_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( L2BroadcastHub_io_inner_grant_bits_data ),
       .io_inner_grant_bits_client_id( L2BroadcastHub_io_inner_grant_bits_client_id ),
       .io_inner_finish_ready( L2BroadcastHub_io_inner_finish_ready ),
       .io_inner_finish_valid( l1tol2net_io_managers_0_finish_valid ),
       .io_inner_finish_bits_manager_xact_id( l1tol2net_io_managers_0_finish_bits_manager_xact_id ),
       .io_inner_probe_ready( l1tol2net_io_managers_0_probe_ready ),
       .io_inner_probe_valid( L2BroadcastHub_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( L2BroadcastHub_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( L2BroadcastHub_io_inner_probe_bits_p_type ),
       .io_inner_probe_bits_client_id( L2BroadcastHub_io_inner_probe_bits_client_id ),
       .io_inner_release_ready( L2BroadcastHub_io_inner_release_ready ),
       .io_inner_release_valid( l1tol2net_io_managers_0_release_valid ),
       .io_inner_release_bits_addr_beat( l1tol2net_io_managers_0_release_bits_addr_beat ),
       .io_inner_release_bits_addr_block( l1tol2net_io_managers_0_release_bits_addr_block ),
       .io_inner_release_bits_client_xact_id( l1tol2net_io_managers_0_release_bits_client_xact_id ),
       .io_inner_release_bits_voluntary( l1tol2net_io_managers_0_release_bits_voluntary ),
       .io_inner_release_bits_r_type( l1tol2net_io_managers_0_release_bits_r_type ),
       .io_inner_release_bits_data( l1tol2net_io_managers_0_release_bits_data ),
       .io_inner_release_bits_client_id( l1tol2net_io_managers_0_release_bits_client_id ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_outer_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_outer_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data )
  );
  NastiRecursiveInterconnect_1 interconnect(.clk(clk), .reset(reset),
       .io_masters_1_aw_ready( interconnect_io_masters_1_aw_ready ),
       .io_masters_1_aw_valid( rtc_io_aw_valid ),
       .io_masters_1_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_masters_1_aw_bits_len( rtc_io_aw_bits_len ),
       .io_masters_1_aw_bits_size( rtc_io_aw_bits_size ),
       .io_masters_1_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_masters_1_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_masters_1_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_masters_1_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_masters_1_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_masters_1_aw_bits_region( rtc_io_aw_bits_region ),
       .io_masters_1_aw_bits_id( rtc_io_aw_bits_id ),
       .io_masters_1_aw_bits_user( rtc_io_aw_bits_user ),
       .io_masters_1_w_ready( interconnect_io_masters_1_w_ready ),
       .io_masters_1_w_valid( rtc_io_w_valid ),
       .io_masters_1_w_bits_data( rtc_io_w_bits_data ),
       .io_masters_1_w_bits_last( rtc_io_w_bits_last ),
       .io_masters_1_w_bits_strb( rtc_io_w_bits_strb ),
       .io_masters_1_w_bits_user( rtc_io_w_bits_user ),
       .io_masters_1_b_ready( rtc_io_b_ready ),
       .io_masters_1_b_valid( interconnect_io_masters_1_b_valid ),
       .io_masters_1_b_bits_resp( interconnect_io_masters_1_b_bits_resp ),
       .io_masters_1_b_bits_id( interconnect_io_masters_1_b_bits_id ),
       .io_masters_1_b_bits_user( interconnect_io_masters_1_b_bits_user ),
       .io_masters_1_ar_ready( interconnect_io_masters_1_ar_ready ),
       .io_masters_1_ar_valid( rtc_io_ar_valid ),
       //.io_masters_1_ar_bits_addr(  )
       //.io_masters_1_ar_bits_len(  )
       //.io_masters_1_ar_bits_size(  )
       //.io_masters_1_ar_bits_burst(  )
       //.io_masters_1_ar_bits_lock(  )
       //.io_masters_1_ar_bits_cache(  )
       //.io_masters_1_ar_bits_prot(  )
       //.io_masters_1_ar_bits_qos(  )
       //.io_masters_1_ar_bits_region(  )
       //.io_masters_1_ar_bits_id(  )
       //.io_masters_1_ar_bits_user(  )
       .io_masters_1_r_ready( rtc_io_r_ready ),
       .io_masters_1_r_valid( interconnect_io_masters_1_r_valid ),
       .io_masters_1_r_bits_resp( interconnect_io_masters_1_r_bits_resp ),
       .io_masters_1_r_bits_data( interconnect_io_masters_1_r_bits_data ),
       .io_masters_1_r_bits_last( interconnect_io_masters_1_r_bits_last ),
       .io_masters_1_r_bits_id( interconnect_io_masters_1_r_bits_id ),
       .io_masters_1_r_bits_user( interconnect_io_masters_1_r_bits_user ),
       .io_masters_0_aw_ready( interconnect_io_masters_0_aw_ready ),
       .io_masters_0_aw_valid( Queue_1_io_deq_valid ),
       .io_masters_0_aw_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_masters_0_aw_bits_len( Queue_1_io_deq_bits_len ),
       .io_masters_0_aw_bits_size( Queue_1_io_deq_bits_size ),
       .io_masters_0_aw_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_masters_0_aw_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_masters_0_aw_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_masters_0_aw_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_masters_0_aw_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_masters_0_aw_bits_region( Queue_1_io_deq_bits_region ),
       .io_masters_0_aw_bits_id( Queue_1_io_deq_bits_id ),
       .io_masters_0_aw_bits_user( Queue_1_io_deq_bits_user ),
       .io_masters_0_w_ready( interconnect_io_masters_0_w_ready ),
       .io_masters_0_w_valid( Queue_2_io_deq_valid ),
       .io_masters_0_w_bits_data( Queue_2_io_deq_bits_data ),
       .io_masters_0_w_bits_last( Queue_2_io_deq_bits_last ),
       .io_masters_0_w_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_masters_0_w_bits_user( Queue_2_io_deq_bits_user ),
       .io_masters_0_b_ready( Queue_4_io_enq_ready ),
       .io_masters_0_b_valid( interconnect_io_masters_0_b_valid ),
       .io_masters_0_b_bits_resp( interconnect_io_masters_0_b_bits_resp ),
       .io_masters_0_b_bits_id( interconnect_io_masters_0_b_bits_id ),
       .io_masters_0_b_bits_user( interconnect_io_masters_0_b_bits_user ),
       .io_masters_0_ar_ready( interconnect_io_masters_0_ar_ready ),
       .io_masters_0_ar_valid( Queue_io_deq_valid ),
       .io_masters_0_ar_bits_addr( Queue_io_deq_bits_addr ),
       .io_masters_0_ar_bits_len( Queue_io_deq_bits_len ),
       .io_masters_0_ar_bits_size( Queue_io_deq_bits_size ),
       .io_masters_0_ar_bits_burst( Queue_io_deq_bits_burst ),
       .io_masters_0_ar_bits_lock( Queue_io_deq_bits_lock ),
       .io_masters_0_ar_bits_cache( Queue_io_deq_bits_cache ),
       .io_masters_0_ar_bits_prot( Queue_io_deq_bits_prot ),
       .io_masters_0_ar_bits_qos( Queue_io_deq_bits_qos ),
       .io_masters_0_ar_bits_region( Queue_io_deq_bits_region ),
       .io_masters_0_ar_bits_id( Queue_io_deq_bits_id ),
       .io_masters_0_ar_bits_user( Queue_io_deq_bits_user ),
       .io_masters_0_r_ready( Queue_3_io_enq_ready ),
       .io_masters_0_r_valid( interconnect_io_masters_0_r_valid ),
       .io_masters_0_r_bits_resp( interconnect_io_masters_0_r_bits_resp ),
       .io_masters_0_r_bits_data( interconnect_io_masters_0_r_bits_data ),
       .io_masters_0_r_bits_last( interconnect_io_masters_0_r_bits_last ),
       .io_masters_0_r_bits_id( interconnect_io_masters_0_r_bits_id ),
       .io_masters_0_r_bits_user( interconnect_io_masters_0_r_bits_user ),
       .io_slaves_4_aw_ready( io_mmio_aw_ready ),
       .io_slaves_4_aw_valid( interconnect_io_slaves_4_aw_valid ),
       .io_slaves_4_aw_bits_addr( interconnect_io_slaves_4_aw_bits_addr ),
       .io_slaves_4_aw_bits_len( interconnect_io_slaves_4_aw_bits_len ),
       .io_slaves_4_aw_bits_size( interconnect_io_slaves_4_aw_bits_size ),
       .io_slaves_4_aw_bits_burst( interconnect_io_slaves_4_aw_bits_burst ),
       .io_slaves_4_aw_bits_lock( interconnect_io_slaves_4_aw_bits_lock ),
       .io_slaves_4_aw_bits_cache( interconnect_io_slaves_4_aw_bits_cache ),
       .io_slaves_4_aw_bits_prot( interconnect_io_slaves_4_aw_bits_prot ),
       .io_slaves_4_aw_bits_qos( interconnect_io_slaves_4_aw_bits_qos ),
       .io_slaves_4_aw_bits_region( interconnect_io_slaves_4_aw_bits_region ),
       .io_slaves_4_aw_bits_id( interconnect_io_slaves_4_aw_bits_id ),
       .io_slaves_4_aw_bits_user( interconnect_io_slaves_4_aw_bits_user ),
       .io_slaves_4_w_ready( io_mmio_w_ready ),
       .io_slaves_4_w_valid( interconnect_io_slaves_4_w_valid ),
       .io_slaves_4_w_bits_data( interconnect_io_slaves_4_w_bits_data ),
       .io_slaves_4_w_bits_last( interconnect_io_slaves_4_w_bits_last ),
       .io_slaves_4_w_bits_strb( interconnect_io_slaves_4_w_bits_strb ),
       .io_slaves_4_w_bits_user( interconnect_io_slaves_4_w_bits_user ),
       .io_slaves_4_b_ready( interconnect_io_slaves_4_b_ready ),
       .io_slaves_4_b_valid( io_mmio_b_valid ),
       .io_slaves_4_b_bits_resp( io_mmio_b_bits_resp ),
       .io_slaves_4_b_bits_id( io_mmio_b_bits_id ),
       .io_slaves_4_b_bits_user( io_mmio_b_bits_user ),
       .io_slaves_4_ar_ready( io_mmio_ar_ready ),
       .io_slaves_4_ar_valid( interconnect_io_slaves_4_ar_valid ),
       .io_slaves_4_ar_bits_addr( interconnect_io_slaves_4_ar_bits_addr ),
       .io_slaves_4_ar_bits_len( interconnect_io_slaves_4_ar_bits_len ),
       .io_slaves_4_ar_bits_size( interconnect_io_slaves_4_ar_bits_size ),
       .io_slaves_4_ar_bits_burst( interconnect_io_slaves_4_ar_bits_burst ),
       .io_slaves_4_ar_bits_lock( interconnect_io_slaves_4_ar_bits_lock ),
       .io_slaves_4_ar_bits_cache( interconnect_io_slaves_4_ar_bits_cache ),
       .io_slaves_4_ar_bits_prot( interconnect_io_slaves_4_ar_bits_prot ),
       .io_slaves_4_ar_bits_qos( interconnect_io_slaves_4_ar_bits_qos ),
       .io_slaves_4_ar_bits_region( interconnect_io_slaves_4_ar_bits_region ),
       .io_slaves_4_ar_bits_id( interconnect_io_slaves_4_ar_bits_id ),
       .io_slaves_4_ar_bits_user( interconnect_io_slaves_4_ar_bits_user ),
       .io_slaves_4_r_ready( interconnect_io_slaves_4_r_ready ),
       .io_slaves_4_r_valid( io_mmio_r_valid ),
       .io_slaves_4_r_bits_resp( io_mmio_r_bits_resp ),
       .io_slaves_4_r_bits_data( io_mmio_r_bits_data ),
       .io_slaves_4_r_bits_last( io_mmio_r_bits_last ),
       .io_slaves_4_r_bits_id( io_mmio_r_bits_id ),
       .io_slaves_4_r_bits_user( io_mmio_r_bits_user ),
       .io_slaves_3_aw_ready( conv_io_nasti_aw_ready ),
       .io_slaves_3_aw_valid( interconnect_io_slaves_3_aw_valid ),
       .io_slaves_3_aw_bits_addr( interconnect_io_slaves_3_aw_bits_addr ),
       .io_slaves_3_aw_bits_len( interconnect_io_slaves_3_aw_bits_len ),
       .io_slaves_3_aw_bits_size( interconnect_io_slaves_3_aw_bits_size ),
       .io_slaves_3_aw_bits_burst( interconnect_io_slaves_3_aw_bits_burst ),
       .io_slaves_3_aw_bits_lock( interconnect_io_slaves_3_aw_bits_lock ),
       .io_slaves_3_aw_bits_cache( interconnect_io_slaves_3_aw_bits_cache ),
       .io_slaves_3_aw_bits_prot( interconnect_io_slaves_3_aw_bits_prot ),
       .io_slaves_3_aw_bits_qos( interconnect_io_slaves_3_aw_bits_qos ),
       .io_slaves_3_aw_bits_region( interconnect_io_slaves_3_aw_bits_region ),
       .io_slaves_3_aw_bits_id( interconnect_io_slaves_3_aw_bits_id ),
       .io_slaves_3_aw_bits_user( interconnect_io_slaves_3_aw_bits_user ),
       .io_slaves_3_w_ready( conv_io_nasti_w_ready ),
       .io_slaves_3_w_valid( interconnect_io_slaves_3_w_valid ),
       .io_slaves_3_w_bits_data( interconnect_io_slaves_3_w_bits_data ),
       .io_slaves_3_w_bits_last( interconnect_io_slaves_3_w_bits_last ),
       .io_slaves_3_w_bits_strb( interconnect_io_slaves_3_w_bits_strb ),
       .io_slaves_3_w_bits_user( interconnect_io_slaves_3_w_bits_user ),
       .io_slaves_3_b_ready( interconnect_io_slaves_3_b_ready ),
       .io_slaves_3_b_valid( conv_io_nasti_b_valid ),
       .io_slaves_3_b_bits_resp( conv_io_nasti_b_bits_resp ),
       .io_slaves_3_b_bits_id( conv_io_nasti_b_bits_id ),
       .io_slaves_3_b_bits_user( conv_io_nasti_b_bits_user ),
       .io_slaves_3_ar_ready( conv_io_nasti_ar_ready ),
       .io_slaves_3_ar_valid( interconnect_io_slaves_3_ar_valid ),
       .io_slaves_3_ar_bits_addr( interconnect_io_slaves_3_ar_bits_addr ),
       .io_slaves_3_ar_bits_len( interconnect_io_slaves_3_ar_bits_len ),
       .io_slaves_3_ar_bits_size( interconnect_io_slaves_3_ar_bits_size ),
       .io_slaves_3_ar_bits_burst( interconnect_io_slaves_3_ar_bits_burst ),
       .io_slaves_3_ar_bits_lock( interconnect_io_slaves_3_ar_bits_lock ),
       .io_slaves_3_ar_bits_cache( interconnect_io_slaves_3_ar_bits_cache ),
       .io_slaves_3_ar_bits_prot( interconnect_io_slaves_3_ar_bits_prot ),
       .io_slaves_3_ar_bits_qos( interconnect_io_slaves_3_ar_bits_qos ),
       .io_slaves_3_ar_bits_region( interconnect_io_slaves_3_ar_bits_region ),
       .io_slaves_3_ar_bits_id( interconnect_io_slaves_3_ar_bits_id ),
       .io_slaves_3_ar_bits_user( interconnect_io_slaves_3_ar_bits_user ),
       .io_slaves_3_r_ready( interconnect_io_slaves_3_r_ready ),
       .io_slaves_3_r_valid( conv_io_nasti_r_valid ),
       .io_slaves_3_r_bits_resp( conv_io_nasti_r_bits_resp ),
       .io_slaves_3_r_bits_data( conv_io_nasti_r_bits_data ),
       .io_slaves_3_r_bits_last( conv_io_nasti_r_bits_last ),
       .io_slaves_3_r_bits_id( conv_io_nasti_r_bits_id ),
       .io_slaves_3_r_bits_user( conv_io_nasti_r_bits_user ),
       .io_slaves_2_aw_ready( SMIIONastiIOConverter_io_nasti_aw_ready ),
       .io_slaves_2_aw_valid( interconnect_io_slaves_2_aw_valid ),
       .io_slaves_2_aw_bits_addr( interconnect_io_slaves_2_aw_bits_addr ),
       .io_slaves_2_aw_bits_len( interconnect_io_slaves_2_aw_bits_len ),
       .io_slaves_2_aw_bits_size( interconnect_io_slaves_2_aw_bits_size ),
       .io_slaves_2_aw_bits_burst( interconnect_io_slaves_2_aw_bits_burst ),
       .io_slaves_2_aw_bits_lock( interconnect_io_slaves_2_aw_bits_lock ),
       .io_slaves_2_aw_bits_cache( interconnect_io_slaves_2_aw_bits_cache ),
       .io_slaves_2_aw_bits_prot( interconnect_io_slaves_2_aw_bits_prot ),
       .io_slaves_2_aw_bits_qos( interconnect_io_slaves_2_aw_bits_qos ),
       .io_slaves_2_aw_bits_region( interconnect_io_slaves_2_aw_bits_region ),
       .io_slaves_2_aw_bits_id( interconnect_io_slaves_2_aw_bits_id ),
       .io_slaves_2_aw_bits_user( interconnect_io_slaves_2_aw_bits_user ),
       .io_slaves_2_w_ready( SMIIONastiIOConverter_io_nasti_w_ready ),
       .io_slaves_2_w_valid( interconnect_io_slaves_2_w_valid ),
       .io_slaves_2_w_bits_data( interconnect_io_slaves_2_w_bits_data ),
       .io_slaves_2_w_bits_last( interconnect_io_slaves_2_w_bits_last ),
       .io_slaves_2_w_bits_strb( interconnect_io_slaves_2_w_bits_strb ),
       .io_slaves_2_w_bits_user( interconnect_io_slaves_2_w_bits_user ),
       .io_slaves_2_b_ready( interconnect_io_slaves_2_b_ready ),
       .io_slaves_2_b_valid( SMIIONastiIOConverter_io_nasti_b_valid ),
       .io_slaves_2_b_bits_resp( SMIIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_slaves_2_b_bits_id( SMIIONastiIOConverter_io_nasti_b_bits_id ),
       .io_slaves_2_b_bits_user( SMIIONastiIOConverter_io_nasti_b_bits_user ),
       .io_slaves_2_ar_ready( SMIIONastiIOConverter_io_nasti_ar_ready ),
       .io_slaves_2_ar_valid( interconnect_io_slaves_2_ar_valid ),
       .io_slaves_2_ar_bits_addr( interconnect_io_slaves_2_ar_bits_addr ),
       .io_slaves_2_ar_bits_len( interconnect_io_slaves_2_ar_bits_len ),
       .io_slaves_2_ar_bits_size( interconnect_io_slaves_2_ar_bits_size ),
       .io_slaves_2_ar_bits_burst( interconnect_io_slaves_2_ar_bits_burst ),
       .io_slaves_2_ar_bits_lock( interconnect_io_slaves_2_ar_bits_lock ),
       .io_slaves_2_ar_bits_cache( interconnect_io_slaves_2_ar_bits_cache ),
       .io_slaves_2_ar_bits_prot( interconnect_io_slaves_2_ar_bits_prot ),
       .io_slaves_2_ar_bits_qos( interconnect_io_slaves_2_ar_bits_qos ),
       .io_slaves_2_ar_bits_region( interconnect_io_slaves_2_ar_bits_region ),
       .io_slaves_2_ar_bits_id( interconnect_io_slaves_2_ar_bits_id ),
       .io_slaves_2_ar_bits_user( interconnect_io_slaves_2_ar_bits_user ),
       .io_slaves_2_r_ready( interconnect_io_slaves_2_r_ready ),
       .io_slaves_2_r_valid( SMIIONastiIOConverter_io_nasti_r_valid ),
       .io_slaves_2_r_bits_resp( SMIIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_slaves_2_r_bits_data( SMIIONastiIOConverter_io_nasti_r_bits_data ),
       .io_slaves_2_r_bits_last( SMIIONastiIOConverter_io_nasti_r_bits_last ),
       .io_slaves_2_r_bits_id( SMIIONastiIOConverter_io_nasti_r_bits_id ),
       .io_slaves_2_r_bits_user( SMIIONastiIOConverter_io_nasti_r_bits_user ),
       .io_slaves_1_aw_ready( io_deviceTree_aw_ready ),
       .io_slaves_1_aw_valid( interconnect_io_slaves_1_aw_valid ),
       .io_slaves_1_aw_bits_addr( interconnect_io_slaves_1_aw_bits_addr ),
       .io_slaves_1_aw_bits_len( interconnect_io_slaves_1_aw_bits_len ),
       .io_slaves_1_aw_bits_size( interconnect_io_slaves_1_aw_bits_size ),
       .io_slaves_1_aw_bits_burst( interconnect_io_slaves_1_aw_bits_burst ),
       .io_slaves_1_aw_bits_lock( interconnect_io_slaves_1_aw_bits_lock ),
       .io_slaves_1_aw_bits_cache( interconnect_io_slaves_1_aw_bits_cache ),
       .io_slaves_1_aw_bits_prot( interconnect_io_slaves_1_aw_bits_prot ),
       .io_slaves_1_aw_bits_qos( interconnect_io_slaves_1_aw_bits_qos ),
       .io_slaves_1_aw_bits_region( interconnect_io_slaves_1_aw_bits_region ),
       .io_slaves_1_aw_bits_id( interconnect_io_slaves_1_aw_bits_id ),
       .io_slaves_1_aw_bits_user( interconnect_io_slaves_1_aw_bits_user ),
       .io_slaves_1_w_ready( io_deviceTree_w_ready ),
       .io_slaves_1_w_valid( interconnect_io_slaves_1_w_valid ),
       .io_slaves_1_w_bits_data( interconnect_io_slaves_1_w_bits_data ),
       .io_slaves_1_w_bits_last( interconnect_io_slaves_1_w_bits_last ),
       .io_slaves_1_w_bits_strb( interconnect_io_slaves_1_w_bits_strb ),
       .io_slaves_1_w_bits_user( interconnect_io_slaves_1_w_bits_user ),
       .io_slaves_1_b_ready( interconnect_io_slaves_1_b_ready ),
       .io_slaves_1_b_valid( io_deviceTree_b_valid ),
       .io_slaves_1_b_bits_resp( io_deviceTree_b_bits_resp ),
       .io_slaves_1_b_bits_id( io_deviceTree_b_bits_id ),
       .io_slaves_1_b_bits_user( io_deviceTree_b_bits_user ),
       .io_slaves_1_ar_ready( io_deviceTree_ar_ready ),
       .io_slaves_1_ar_valid( interconnect_io_slaves_1_ar_valid ),
       .io_slaves_1_ar_bits_addr( interconnect_io_slaves_1_ar_bits_addr ),
       .io_slaves_1_ar_bits_len( interconnect_io_slaves_1_ar_bits_len ),
       .io_slaves_1_ar_bits_size( interconnect_io_slaves_1_ar_bits_size ),
       .io_slaves_1_ar_bits_burst( interconnect_io_slaves_1_ar_bits_burst ),
       .io_slaves_1_ar_bits_lock( interconnect_io_slaves_1_ar_bits_lock ),
       .io_slaves_1_ar_bits_cache( interconnect_io_slaves_1_ar_bits_cache ),
       .io_slaves_1_ar_bits_prot( interconnect_io_slaves_1_ar_bits_prot ),
       .io_slaves_1_ar_bits_qos( interconnect_io_slaves_1_ar_bits_qos ),
       .io_slaves_1_ar_bits_region( interconnect_io_slaves_1_ar_bits_region ),
       .io_slaves_1_ar_bits_id( interconnect_io_slaves_1_ar_bits_id ),
       .io_slaves_1_ar_bits_user( interconnect_io_slaves_1_ar_bits_user ),
       .io_slaves_1_r_ready( interconnect_io_slaves_1_r_ready ),
       .io_slaves_1_r_valid( io_deviceTree_r_valid ),
       .io_slaves_1_r_bits_resp( io_deviceTree_r_bits_resp ),
       .io_slaves_1_r_bits_data( io_deviceTree_r_bits_data ),
       .io_slaves_1_r_bits_last( io_deviceTree_r_bits_last ),
       .io_slaves_1_r_bits_id( io_deviceTree_r_bits_id ),
       .io_slaves_1_r_bits_user( io_deviceTree_r_bits_user ),
       .io_slaves_0_aw_ready( io_mem_0_aw_ready ),
       .io_slaves_0_aw_valid( interconnect_io_slaves_0_aw_valid ),
       .io_slaves_0_aw_bits_addr( interconnect_io_slaves_0_aw_bits_addr ),
       .io_slaves_0_aw_bits_len( interconnect_io_slaves_0_aw_bits_len ),
       .io_slaves_0_aw_bits_size( interconnect_io_slaves_0_aw_bits_size ),
       .io_slaves_0_aw_bits_burst( interconnect_io_slaves_0_aw_bits_burst ),
       .io_slaves_0_aw_bits_lock( interconnect_io_slaves_0_aw_bits_lock ),
       .io_slaves_0_aw_bits_cache( interconnect_io_slaves_0_aw_bits_cache ),
       .io_slaves_0_aw_bits_prot( interconnect_io_slaves_0_aw_bits_prot ),
       .io_slaves_0_aw_bits_qos( interconnect_io_slaves_0_aw_bits_qos ),
       .io_slaves_0_aw_bits_region( interconnect_io_slaves_0_aw_bits_region ),
       .io_slaves_0_aw_bits_id( interconnect_io_slaves_0_aw_bits_id ),
       .io_slaves_0_aw_bits_user( interconnect_io_slaves_0_aw_bits_user ),
       .io_slaves_0_w_ready( io_mem_0_w_ready ),
       .io_slaves_0_w_valid( interconnect_io_slaves_0_w_valid ),
       .io_slaves_0_w_bits_data( interconnect_io_slaves_0_w_bits_data ),
       .io_slaves_0_w_bits_last( interconnect_io_slaves_0_w_bits_last ),
       .io_slaves_0_w_bits_strb( interconnect_io_slaves_0_w_bits_strb ),
       .io_slaves_0_w_bits_user( interconnect_io_slaves_0_w_bits_user ),
       .io_slaves_0_b_ready( interconnect_io_slaves_0_b_ready ),
       .io_slaves_0_b_valid( io_mem_0_b_valid ),
       .io_slaves_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_slaves_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_slaves_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_slaves_0_ar_ready( io_mem_0_ar_ready ),
       .io_slaves_0_ar_valid( interconnect_io_slaves_0_ar_valid ),
       .io_slaves_0_ar_bits_addr( interconnect_io_slaves_0_ar_bits_addr ),
       .io_slaves_0_ar_bits_len( interconnect_io_slaves_0_ar_bits_len ),
       .io_slaves_0_ar_bits_size( interconnect_io_slaves_0_ar_bits_size ),
       .io_slaves_0_ar_bits_burst( interconnect_io_slaves_0_ar_bits_burst ),
       .io_slaves_0_ar_bits_lock( interconnect_io_slaves_0_ar_bits_lock ),
       .io_slaves_0_ar_bits_cache( interconnect_io_slaves_0_ar_bits_cache ),
       .io_slaves_0_ar_bits_prot( interconnect_io_slaves_0_ar_bits_prot ),
       .io_slaves_0_ar_bits_qos( interconnect_io_slaves_0_ar_bits_qos ),
       .io_slaves_0_ar_bits_region( interconnect_io_slaves_0_ar_bits_region ),
       .io_slaves_0_ar_bits_id( interconnect_io_slaves_0_ar_bits_id ),
       .io_slaves_0_ar_bits_user( interconnect_io_slaves_0_ar_bits_user ),
       .io_slaves_0_r_ready( interconnect_io_slaves_0_r_ready ),
       .io_slaves_0_r_valid( io_mem_0_r_valid ),
       .io_slaves_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_slaves_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_slaves_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_slaves_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_slaves_0_r_bits_user( io_mem_0_r_bits_user )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign interconnect.io_masters_1_ar_bits_addr = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_len = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_size = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_burst = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_lock = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_cache = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_prot = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_qos = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_region = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_id = {1{$random}};
    assign interconnect.io_masters_1_ar_bits_user = {1{$random}};
// synthesis translate_on
`endif
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper(.clk(clk), .reset(reset),
       .io_in_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkEnqueuer_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkEnqueuer_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkEnqueuer_io_outer_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkEnqueuer_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_in_probe_ready( ClientTileLinkEnqueuer_io_outer_probe_ready ),
       .io_in_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_in_probe_bits_addr_block(  )
       //.io_in_probe_bits_p_type(  )
       .io_in_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_in_release_valid( ClientTileLinkEnqueuer_io_outer_release_valid ),
       .io_in_release_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat ),
       .io_in_release_bits_addr_block( ClientTileLinkEnqueuer_io_outer_release_bits_addr_block ),
       .io_in_release_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id ),
       .io_in_release_bits_voluntary( ClientTileLinkEnqueuer_io_outer_release_bits_voluntary ),
       .io_in_release_bits_r_type( ClientTileLinkEnqueuer_io_outer_release_bits_r_type ),
       .io_in_release_bits_data( ClientTileLinkEnqueuer_io_outer_release_bits_data ),
       .io_out_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_out_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_out_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_out_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data )
  );
  TileLinkIONarrower TileLinkIONarrower(.clk(clk), .reset(reset),
       .io_in_acquire_ready( TileLinkIONarrower_io_in_acquire_ready ),
       .io_in_acquire_valid( ClientTileLinkIOUnwrapper_io_out_acquire_valid ),
       .io_in_acquire_bits_addr_block( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_out_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( ClientTileLinkIOUnwrapper_io_out_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( ClientTileLinkIOUnwrapper_io_out_acquire_bits_a_type ),
       .io_in_acquire_bits_union( ClientTileLinkIOUnwrapper_io_out_acquire_bits_union ),
       .io_in_acquire_bits_data( ClientTileLinkIOUnwrapper_io_out_acquire_bits_data ),
       .io_in_grant_ready( ClientTileLinkIOUnwrapper_io_out_grant_ready ),
       .io_in_grant_valid( TileLinkIONarrower_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( TileLinkIONarrower_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( TileLinkIONarrower_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( TileLinkIONarrower_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( TileLinkIONarrower_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( TileLinkIONarrower_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( TileLinkIONarrower_io_in_grant_bits_data ),
       .io_out_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_out_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_out_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_out_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_out_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_out_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data )
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter(.clk(clk), .reset(reset),
       .io_tl_acquire_ready( NastiIOTileLinkIOConverter_io_tl_acquire_ready ),
       .io_tl_acquire_valid( TileLinkIONarrower_io_out_acquire_valid ),
       .io_tl_acquire_bits_addr_block( TileLinkIONarrower_io_out_acquire_bits_addr_block ),
       .io_tl_acquire_bits_client_xact_id( TileLinkIONarrower_io_out_acquire_bits_client_xact_id ),
       .io_tl_acquire_bits_addr_beat( TileLinkIONarrower_io_out_acquire_bits_addr_beat ),
       .io_tl_acquire_bits_is_builtin_type( TileLinkIONarrower_io_out_acquire_bits_is_builtin_type ),
       .io_tl_acquire_bits_a_type( TileLinkIONarrower_io_out_acquire_bits_a_type ),
       .io_tl_acquire_bits_union( TileLinkIONarrower_io_out_acquire_bits_union ),
       .io_tl_acquire_bits_data( TileLinkIONarrower_io_out_acquire_bits_data ),
       .io_tl_grant_ready( TileLinkIONarrower_io_out_grant_ready ),
       .io_tl_grant_valid( NastiIOTileLinkIOConverter_io_tl_grant_valid ),
       .io_tl_grant_bits_addr_beat( NastiIOTileLinkIOConverter_io_tl_grant_bits_addr_beat ),
       .io_tl_grant_bits_client_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_client_xact_id ),
       .io_tl_grant_bits_manager_xact_id( NastiIOTileLinkIOConverter_io_tl_grant_bits_manager_xact_id ),
       .io_tl_grant_bits_is_builtin_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_is_builtin_type ),
       .io_tl_grant_bits_g_type( NastiIOTileLinkIOConverter_io_tl_grant_bits_g_type ),
       .io_tl_grant_bits_data( NastiIOTileLinkIOConverter_io_tl_grant_bits_data ),
       .io_nasti_aw_ready( Queue_1_io_enq_ready ),
       .io_nasti_aw_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_nasti_aw_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_nasti_aw_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_nasti_aw_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_nasti_aw_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_nasti_aw_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_nasti_aw_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_nasti_aw_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_nasti_aw_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_nasti_aw_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_nasti_aw_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_nasti_aw_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_nasti_w_ready( Queue_2_io_enq_ready ),
       .io_nasti_w_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_nasti_w_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_nasti_w_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_nasti_w_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_nasti_w_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_nasti_b_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_nasti_b_valid( Queue_4_io_deq_valid ),
       .io_nasti_b_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_nasti_b_bits_id( Queue_4_io_deq_bits_id ),
       .io_nasti_b_bits_user( Queue_4_io_deq_bits_user ),
       .io_nasti_ar_ready( Queue_io_enq_ready ),
       .io_nasti_ar_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_nasti_ar_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_nasti_ar_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_nasti_ar_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_nasti_ar_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_nasti_ar_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_nasti_ar_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_nasti_ar_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_nasti_ar_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_nasti_ar_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_nasti_ar_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_nasti_ar_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_nasti_r_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_nasti_r_valid( Queue_3_io_deq_valid ),
       .io_nasti_r_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_nasti_r_bits_data( Queue_3_io_deq_bits_data ),
       .io_nasti_r_bits_last( Queue_3_io_deq_bits_last ),
       .io_nasti_r_bits_id( Queue_3_io_deq_bits_id ),
       .io_nasti_r_bits_user( Queue_3_io_deq_bits_user )
  );
  ClientTileLinkIOWrapper_1 ClientTileLinkIOWrapper_2(
       .io_in_acquire_ready( ClientTileLinkIOWrapper_2_io_in_acquire_ready ),
       .io_in_acquire_valid( L2BroadcastHub_io_outer_acquire_valid ),
       .io_in_acquire_bits_addr_block( L2BroadcastHub_io_outer_acquire_bits_addr_block ),
       .io_in_acquire_bits_client_xact_id( L2BroadcastHub_io_outer_acquire_bits_client_xact_id ),
       .io_in_acquire_bits_addr_beat( L2BroadcastHub_io_outer_acquire_bits_addr_beat ),
       .io_in_acquire_bits_is_builtin_type( L2BroadcastHub_io_outer_acquire_bits_is_builtin_type ),
       .io_in_acquire_bits_a_type( L2BroadcastHub_io_outer_acquire_bits_a_type ),
       .io_in_acquire_bits_union( L2BroadcastHub_io_outer_acquire_bits_union ),
       .io_in_acquire_bits_data( L2BroadcastHub_io_outer_acquire_bits_data ),
       .io_in_grant_ready( L2BroadcastHub_io_outer_grant_ready ),
       .io_in_grant_valid( ClientTileLinkIOWrapper_2_io_in_grant_valid ),
       .io_in_grant_bits_addr_beat( ClientTileLinkIOWrapper_2_io_in_grant_bits_addr_beat ),
       .io_in_grant_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_client_xact_id ),
       .io_in_grant_bits_manager_xact_id( ClientTileLinkIOWrapper_2_io_in_grant_bits_manager_xact_id ),
       .io_in_grant_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_is_builtin_type ),
       .io_in_grant_bits_g_type( ClientTileLinkIOWrapper_2_io_in_grant_bits_g_type ),
       .io_in_grant_bits_data( ClientTileLinkIOWrapper_2_io_in_grant_bits_data ),
       .io_out_acquire_ready( ClientTileLinkEnqueuer_io_inner_acquire_ready ),
       .io_out_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_out_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_out_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_out_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_out_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_out_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_out_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_out_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_out_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_out_grant_valid( ClientTileLinkEnqueuer_io_inner_grant_valid ),
       .io_out_grant_bits_addr_beat( ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat ),
       .io_out_grant_bits_client_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id ),
       .io_out_grant_bits_manager_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id ),
       .io_out_grant_bits_is_builtin_type( ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type ),
       .io_out_grant_bits_g_type( ClientTileLinkEnqueuer_io_inner_grant_bits_g_type ),
       .io_out_grant_bits_data( ClientTileLinkEnqueuer_io_inner_grant_bits_data ),
       .io_out_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_out_probe_valid( ClientTileLinkEnqueuer_io_inner_probe_valid ),
       .io_out_probe_bits_addr_block( ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block ),
       .io_out_probe_bits_p_type( ClientTileLinkEnqueuer_io_inner_probe_bits_p_type ),
       .io_out_release_ready( ClientTileLinkEnqueuer_io_inner_release_ready ),
       .io_out_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid )
       //.io_out_release_bits_addr_beat(  )
       //.io_out_release_bits_addr_block(  )
       //.io_out_release_bits_client_xact_id(  )
       //.io_out_release_bits_voluntary(  )
       //.io_out_release_bits_r_type(  )
       //.io_out_release_bits_data(  )
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer(
       .io_inner_acquire_ready( ClientTileLinkEnqueuer_io_inner_acquire_ready ),
       .io_inner_acquire_valid( ClientTileLinkIOWrapper_2_io_out_acquire_valid ),
       .io_inner_acquire_bits_addr_block( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_block ),
       .io_inner_acquire_bits_client_xact_id( ClientTileLinkIOWrapper_2_io_out_acquire_bits_client_xact_id ),
       .io_inner_acquire_bits_addr_beat( ClientTileLinkIOWrapper_2_io_out_acquire_bits_addr_beat ),
       .io_inner_acquire_bits_is_builtin_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_is_builtin_type ),
       .io_inner_acquire_bits_a_type( ClientTileLinkIOWrapper_2_io_out_acquire_bits_a_type ),
       .io_inner_acquire_bits_union( ClientTileLinkIOWrapper_2_io_out_acquire_bits_union ),
       .io_inner_acquire_bits_data( ClientTileLinkIOWrapper_2_io_out_acquire_bits_data ),
       .io_inner_grant_ready( ClientTileLinkIOWrapper_2_io_out_grant_ready ),
       .io_inner_grant_valid( ClientTileLinkEnqueuer_io_inner_grant_valid ),
       .io_inner_grant_bits_addr_beat( ClientTileLinkEnqueuer_io_inner_grant_bits_addr_beat ),
       .io_inner_grant_bits_client_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_client_xact_id ),
       .io_inner_grant_bits_manager_xact_id( ClientTileLinkEnqueuer_io_inner_grant_bits_manager_xact_id ),
       .io_inner_grant_bits_is_builtin_type( ClientTileLinkEnqueuer_io_inner_grant_bits_is_builtin_type ),
       .io_inner_grant_bits_g_type( ClientTileLinkEnqueuer_io_inner_grant_bits_g_type ),
       .io_inner_grant_bits_data( ClientTileLinkEnqueuer_io_inner_grant_bits_data ),
       .io_inner_probe_ready( ClientTileLinkIOWrapper_2_io_out_probe_ready ),
       .io_inner_probe_valid( ClientTileLinkEnqueuer_io_inner_probe_valid ),
       .io_inner_probe_bits_addr_block( ClientTileLinkEnqueuer_io_inner_probe_bits_addr_block ),
       .io_inner_probe_bits_p_type( ClientTileLinkEnqueuer_io_inner_probe_bits_p_type ),
       .io_inner_release_ready( ClientTileLinkEnqueuer_io_inner_release_ready ),
       .io_inner_release_valid( ClientTileLinkIOWrapper_2_io_out_release_valid ),
       //.io_inner_release_bits_addr_beat(  )
       //.io_inner_release_bits_addr_block(  )
       //.io_inner_release_bits_client_xact_id(  )
       //.io_inner_release_bits_voluntary(  )
       //.io_inner_release_bits_r_type(  )
       //.io_inner_release_bits_data(  )
       .io_outer_acquire_ready( ClientTileLinkIOUnwrapper_io_in_acquire_ready ),
       .io_outer_acquire_valid( ClientTileLinkEnqueuer_io_outer_acquire_valid ),
       .io_outer_acquire_bits_addr_block( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_block ),
       .io_outer_acquire_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_acquire_bits_client_xact_id ),
       .io_outer_acquire_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_acquire_bits_addr_beat ),
       .io_outer_acquire_bits_is_builtin_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_is_builtin_type ),
       .io_outer_acquire_bits_a_type( ClientTileLinkEnqueuer_io_outer_acquire_bits_a_type ),
       .io_outer_acquire_bits_union( ClientTileLinkEnqueuer_io_outer_acquire_bits_union ),
       .io_outer_acquire_bits_data( ClientTileLinkEnqueuer_io_outer_acquire_bits_data ),
       .io_outer_grant_ready( ClientTileLinkEnqueuer_io_outer_grant_ready ),
       .io_outer_grant_valid( ClientTileLinkIOUnwrapper_io_in_grant_valid ),
       .io_outer_grant_bits_addr_beat( ClientTileLinkIOUnwrapper_io_in_grant_bits_addr_beat ),
       .io_outer_grant_bits_client_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_client_xact_id ),
       .io_outer_grant_bits_manager_xact_id( ClientTileLinkIOUnwrapper_io_in_grant_bits_manager_xact_id ),
       .io_outer_grant_bits_is_builtin_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_is_builtin_type ),
       .io_outer_grant_bits_g_type( ClientTileLinkIOUnwrapper_io_in_grant_bits_g_type ),
       .io_outer_grant_bits_data( ClientTileLinkIOUnwrapper_io_in_grant_bits_data ),
       .io_outer_probe_ready( ClientTileLinkEnqueuer_io_outer_probe_ready ),
       .io_outer_probe_valid( ClientTileLinkIOUnwrapper_io_in_probe_valid ),
       //.io_outer_probe_bits_addr_block(  )
       //.io_outer_probe_bits_p_type(  )
       .io_outer_release_ready( ClientTileLinkIOUnwrapper_io_in_release_ready ),
       .io_outer_release_valid( ClientTileLinkEnqueuer_io_outer_release_valid ),
       .io_outer_release_bits_addr_beat( ClientTileLinkEnqueuer_io_outer_release_bits_addr_beat ),
       .io_outer_release_bits_addr_block( ClientTileLinkEnqueuer_io_outer_release_bits_addr_block ),
       .io_outer_release_bits_client_xact_id( ClientTileLinkEnqueuer_io_outer_release_bits_client_xact_id ),
       .io_outer_release_bits_voluntary( ClientTileLinkEnqueuer_io_outer_release_bits_voluntary ),
       .io_outer_release_bits_r_type( ClientTileLinkEnqueuer_io_outer_release_bits_r_type ),
       .io_outer_release_bits_data( ClientTileLinkEnqueuer_io_outer_release_bits_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign ClientTileLinkEnqueuer.io_inner_release_bits_addr_beat = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_addr_block = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_client_xact_id = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_voluntary = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_r_type = {1{$random}};
    assign ClientTileLinkEnqueuer.io_inner_release_bits_data = {4{$random}};
    assign ClientTileLinkEnqueuer.io_outer_probe_bits_addr_block = {1{$random}};
    assign ClientTileLinkEnqueuer.io_outer_probe_bits_p_type = {1{$random}};
// synthesis translate_on
`endif
  Queue_2 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_ar_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_ar_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_ar_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_ar_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_ar_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_ar_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_ar_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_ar_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_ar_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_ar_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_ar_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_ar_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_ar_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_io_deq_bits_len ),
       .io_deq_bits_size( Queue_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_io_deq_bits_region ),
       .io_deq_bits_id( Queue_io_deq_bits_id ),
       .io_deq_bits_user( Queue_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_2 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_aw_valid ),
       .io_enq_bits_addr( NastiIOTileLinkIOConverter_io_nasti_aw_bits_addr ),
       .io_enq_bits_len( NastiIOTileLinkIOConverter_io_nasti_aw_bits_len ),
       .io_enq_bits_size( NastiIOTileLinkIOConverter_io_nasti_aw_bits_size ),
       .io_enq_bits_burst( NastiIOTileLinkIOConverter_io_nasti_aw_bits_burst ),
       .io_enq_bits_lock( NastiIOTileLinkIOConverter_io_nasti_aw_bits_lock ),
       .io_enq_bits_cache( NastiIOTileLinkIOConverter_io_nasti_aw_bits_cache ),
       .io_enq_bits_prot( NastiIOTileLinkIOConverter_io_nasti_aw_bits_prot ),
       .io_enq_bits_qos( NastiIOTileLinkIOConverter_io_nasti_aw_bits_qos ),
       .io_enq_bits_region( NastiIOTileLinkIOConverter_io_nasti_aw_bits_region ),
       .io_enq_bits_id( NastiIOTileLinkIOConverter_io_nasti_aw_bits_id ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_aw_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_aw_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_addr( Queue_1_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_1_io_deq_bits_len ),
       .io_deq_bits_size( Queue_1_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_1_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_1_io_deq_bits_lock ),
       .io_deq_bits_cache( Queue_1_io_deq_bits_cache ),
       .io_deq_bits_prot( Queue_1_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_1_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_1_io_deq_bits_region ),
       .io_deq_bits_id( Queue_1_io_deq_bits_id ),
       .io_deq_bits_user( Queue_1_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( NastiIOTileLinkIOConverter_io_nasti_w_valid ),
       .io_enq_bits_data( NastiIOTileLinkIOConverter_io_nasti_w_bits_data ),
       .io_enq_bits_last( NastiIOTileLinkIOConverter_io_nasti_w_bits_last ),
       .io_enq_bits_strb( NastiIOTileLinkIOConverter_io_nasti_w_bits_strb ),
       .io_enq_bits_user( NastiIOTileLinkIOConverter_io_nasti_w_bits_user ),
       .io_deq_ready( interconnect_io_masters_0_w_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_data( Queue_2_io_deq_bits_data ),
       .io_deq_bits_last( Queue_2_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_2_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_2_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( interconnect_io_masters_0_r_valid ),
       .io_enq_bits_resp( interconnect_io_masters_0_r_bits_resp ),
       .io_enq_bits_data( interconnect_io_masters_0_r_bits_data ),
       .io_enq_bits_last( interconnect_io_masters_0_r_bits_last ),
       .io_enq_bits_id( interconnect_io_masters_0_r_bits_id ),
       .io_enq_bits_user( interconnect_io_masters_0_r_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_r_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_resp( Queue_3_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_3_io_deq_bits_data ),
       .io_deq_bits_last( Queue_3_io_deq_bits_last ),
       .io_deq_bits_id( Queue_3_io_deq_bits_id ),
       .io_deq_bits_user( Queue_3_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( interconnect_io_masters_0_b_valid ),
       .io_enq_bits_resp( interconnect_io_masters_0_b_bits_resp ),
       .io_enq_bits_id( interconnect_io_masters_0_b_bits_id ),
       .io_enq_bits_user( interconnect_io_masters_0_b_bits_user ),
       .io_deq_ready( NastiIOTileLinkIOConverter_io_nasti_b_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_resp( Queue_4_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_4_io_deq_bits_id ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  RTC rtc(.clk(clk), .reset(reset),
       .io_aw_ready( interconnect_io_masters_1_aw_ready ),
       .io_aw_valid( rtc_io_aw_valid ),
       .io_aw_bits_addr( rtc_io_aw_bits_addr ),
       .io_aw_bits_len( rtc_io_aw_bits_len ),
       .io_aw_bits_size( rtc_io_aw_bits_size ),
       .io_aw_bits_burst( rtc_io_aw_bits_burst ),
       .io_aw_bits_lock( rtc_io_aw_bits_lock ),
       .io_aw_bits_cache( rtc_io_aw_bits_cache ),
       .io_aw_bits_prot( rtc_io_aw_bits_prot ),
       .io_aw_bits_qos( rtc_io_aw_bits_qos ),
       .io_aw_bits_region( rtc_io_aw_bits_region ),
       .io_aw_bits_id( rtc_io_aw_bits_id ),
       .io_aw_bits_user( rtc_io_aw_bits_user ),
       .io_w_ready( interconnect_io_masters_1_w_ready ),
       .io_w_valid( rtc_io_w_valid ),
       .io_w_bits_data( rtc_io_w_bits_data ),
       .io_w_bits_last( rtc_io_w_bits_last ),
       .io_w_bits_strb( rtc_io_w_bits_strb ),
       .io_w_bits_user( rtc_io_w_bits_user ),
       .io_b_ready( rtc_io_b_ready ),
       .io_b_valid( interconnect_io_masters_1_b_valid ),
       .io_b_bits_resp( interconnect_io_masters_1_b_bits_resp ),
       .io_b_bits_id( interconnect_io_masters_1_b_bits_id ),
       .io_b_bits_user( interconnect_io_masters_1_b_bits_user ),
       .io_ar_ready( interconnect_io_masters_1_ar_ready ),
       .io_ar_valid( rtc_io_ar_valid ),
       //.io_ar_bits_addr(  )
       //.io_ar_bits_len(  )
       //.io_ar_bits_size(  )
       //.io_ar_bits_burst(  )
       //.io_ar_bits_lock(  )
       //.io_ar_bits_cache(  )
       //.io_ar_bits_prot(  )
       //.io_ar_bits_qos(  )
       //.io_ar_bits_region(  )
       //.io_ar_bits_id(  )
       //.io_ar_bits_user(  )
       .io_r_ready( rtc_io_r_ready ),
       .io_r_valid( interconnect_io_masters_1_r_valid ),
       .io_r_bits_resp( interconnect_io_masters_1_r_bits_resp ),
       .io_r_bits_data( interconnect_io_masters_1_r_bits_data ),
       .io_r_bits_last( interconnect_io_masters_1_r_bits_last ),
       .io_r_bits_id( interconnect_io_masters_1_r_bits_id ),
       .io_r_bits_user( interconnect_io_masters_1_r_bits_user )
  );
  SMIIONastiIOConverter_0 SMIIONastiIOConverter(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( SMIIONastiIOConverter_io_nasti_aw_ready ),
       .io_nasti_aw_valid( interconnect_io_slaves_2_aw_valid ),
       .io_nasti_aw_bits_addr( interconnect_io_slaves_2_aw_bits_addr ),
       .io_nasti_aw_bits_len( interconnect_io_slaves_2_aw_bits_len ),
       .io_nasti_aw_bits_size( interconnect_io_slaves_2_aw_bits_size ),
       .io_nasti_aw_bits_burst( interconnect_io_slaves_2_aw_bits_burst ),
       .io_nasti_aw_bits_lock( interconnect_io_slaves_2_aw_bits_lock ),
       .io_nasti_aw_bits_cache( interconnect_io_slaves_2_aw_bits_cache ),
       .io_nasti_aw_bits_prot( interconnect_io_slaves_2_aw_bits_prot ),
       .io_nasti_aw_bits_qos( interconnect_io_slaves_2_aw_bits_qos ),
       .io_nasti_aw_bits_region( interconnect_io_slaves_2_aw_bits_region ),
       .io_nasti_aw_bits_id( interconnect_io_slaves_2_aw_bits_id ),
       .io_nasti_aw_bits_user( interconnect_io_slaves_2_aw_bits_user ),
       .io_nasti_w_ready( SMIIONastiIOConverter_io_nasti_w_ready ),
       .io_nasti_w_valid( interconnect_io_slaves_2_w_valid ),
       .io_nasti_w_bits_data( interconnect_io_slaves_2_w_bits_data ),
       .io_nasti_w_bits_last( interconnect_io_slaves_2_w_bits_last ),
       .io_nasti_w_bits_strb( interconnect_io_slaves_2_w_bits_strb ),
       .io_nasti_w_bits_user( interconnect_io_slaves_2_w_bits_user ),
       .io_nasti_b_ready( interconnect_io_slaves_2_b_ready ),
       .io_nasti_b_valid( SMIIONastiIOConverter_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( SMIIONastiIOConverter_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( SMIIONastiIOConverter_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( SMIIONastiIOConverter_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( SMIIONastiIOConverter_io_nasti_ar_ready ),
       .io_nasti_ar_valid( interconnect_io_slaves_2_ar_valid ),
       .io_nasti_ar_bits_addr( interconnect_io_slaves_2_ar_bits_addr ),
       .io_nasti_ar_bits_len( interconnect_io_slaves_2_ar_bits_len ),
       .io_nasti_ar_bits_size( interconnect_io_slaves_2_ar_bits_size ),
       .io_nasti_ar_bits_burst( interconnect_io_slaves_2_ar_bits_burst ),
       .io_nasti_ar_bits_lock( interconnect_io_slaves_2_ar_bits_lock ),
       .io_nasti_ar_bits_cache( interconnect_io_slaves_2_ar_bits_cache ),
       .io_nasti_ar_bits_prot( interconnect_io_slaves_2_ar_bits_prot ),
       .io_nasti_ar_bits_qos( interconnect_io_slaves_2_ar_bits_qos ),
       .io_nasti_ar_bits_region( interconnect_io_slaves_2_ar_bits_region ),
       .io_nasti_ar_bits_id( interconnect_io_slaves_2_ar_bits_id ),
       .io_nasti_ar_bits_user( interconnect_io_slaves_2_ar_bits_user ),
       .io_nasti_r_ready( interconnect_io_slaves_2_r_ready ),
       .io_nasti_r_valid( SMIIONastiIOConverter_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( SMIIONastiIOConverter_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( SMIIONastiIOConverter_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( SMIIONastiIOConverter_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( SMIIONastiIOConverter_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( SMIIONastiIOConverter_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_csr_0_req_ready ),
       .io_smi_req_valid( SMIIONastiIOConverter_io_smi_req_valid ),
       .io_smi_req_bits_rw( SMIIONastiIOConverter_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( SMIIONastiIOConverter_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( SMIIONastiIOConverter_io_smi_req_bits_data ),
       .io_smi_resp_ready( SMIIONastiIOConverter_io_smi_resp_ready ),
       .io_smi_resp_valid( io_csr_0_resp_valid ),
       .io_smi_resp_bits( io_csr_0_resp_bits )
  );
  SMIIONastiIOConverter_1 conv(.clk(clk), .reset(reset),
       .io_nasti_aw_ready( conv_io_nasti_aw_ready ),
       .io_nasti_aw_valid( interconnect_io_slaves_3_aw_valid ),
       .io_nasti_aw_bits_addr( interconnect_io_slaves_3_aw_bits_addr ),
       .io_nasti_aw_bits_len( interconnect_io_slaves_3_aw_bits_len ),
       .io_nasti_aw_bits_size( interconnect_io_slaves_3_aw_bits_size ),
       .io_nasti_aw_bits_burst( interconnect_io_slaves_3_aw_bits_burst ),
       .io_nasti_aw_bits_lock( interconnect_io_slaves_3_aw_bits_lock ),
       .io_nasti_aw_bits_cache( interconnect_io_slaves_3_aw_bits_cache ),
       .io_nasti_aw_bits_prot( interconnect_io_slaves_3_aw_bits_prot ),
       .io_nasti_aw_bits_qos( interconnect_io_slaves_3_aw_bits_qos ),
       .io_nasti_aw_bits_region( interconnect_io_slaves_3_aw_bits_region ),
       .io_nasti_aw_bits_id( interconnect_io_slaves_3_aw_bits_id ),
       .io_nasti_aw_bits_user( interconnect_io_slaves_3_aw_bits_user ),
       .io_nasti_w_ready( conv_io_nasti_w_ready ),
       .io_nasti_w_valid( interconnect_io_slaves_3_w_valid ),
       .io_nasti_w_bits_data( interconnect_io_slaves_3_w_bits_data ),
       .io_nasti_w_bits_last( interconnect_io_slaves_3_w_bits_last ),
       .io_nasti_w_bits_strb( interconnect_io_slaves_3_w_bits_strb ),
       .io_nasti_w_bits_user( interconnect_io_slaves_3_w_bits_user ),
       .io_nasti_b_ready( interconnect_io_slaves_3_b_ready ),
       .io_nasti_b_valid( conv_io_nasti_b_valid ),
       .io_nasti_b_bits_resp( conv_io_nasti_b_bits_resp ),
       .io_nasti_b_bits_id( conv_io_nasti_b_bits_id ),
       .io_nasti_b_bits_user( conv_io_nasti_b_bits_user ),
       .io_nasti_ar_ready( conv_io_nasti_ar_ready ),
       .io_nasti_ar_valid( interconnect_io_slaves_3_ar_valid ),
       .io_nasti_ar_bits_addr( interconnect_io_slaves_3_ar_bits_addr ),
       .io_nasti_ar_bits_len( interconnect_io_slaves_3_ar_bits_len ),
       .io_nasti_ar_bits_size( interconnect_io_slaves_3_ar_bits_size ),
       .io_nasti_ar_bits_burst( interconnect_io_slaves_3_ar_bits_burst ),
       .io_nasti_ar_bits_lock( interconnect_io_slaves_3_ar_bits_lock ),
       .io_nasti_ar_bits_cache( interconnect_io_slaves_3_ar_bits_cache ),
       .io_nasti_ar_bits_prot( interconnect_io_slaves_3_ar_bits_prot ),
       .io_nasti_ar_bits_qos( interconnect_io_slaves_3_ar_bits_qos ),
       .io_nasti_ar_bits_region( interconnect_io_slaves_3_ar_bits_region ),
       .io_nasti_ar_bits_id( interconnect_io_slaves_3_ar_bits_id ),
       .io_nasti_ar_bits_user( interconnect_io_slaves_3_ar_bits_user ),
       .io_nasti_r_ready( interconnect_io_slaves_3_r_ready ),
       .io_nasti_r_valid( conv_io_nasti_r_valid ),
       .io_nasti_r_bits_resp( conv_io_nasti_r_bits_resp ),
       .io_nasti_r_bits_data( conv_io_nasti_r_bits_data ),
       .io_nasti_r_bits_last( conv_io_nasti_r_bits_last ),
       .io_nasti_r_bits_id( conv_io_nasti_r_bits_id ),
       .io_nasti_r_bits_user( conv_io_nasti_r_bits_user ),
       .io_smi_req_ready( io_scr_req_ready ),
       .io_smi_req_valid( conv_io_smi_req_valid ),
       .io_smi_req_bits_rw( conv_io_smi_req_bits_rw ),
       .io_smi_req_bits_addr( conv_io_smi_req_bits_addr ),
       .io_smi_req_bits_data( conv_io_smi_req_bits_data ),
       .io_smi_resp_ready( conv_io_smi_resp_ready ),
       .io_smi_resp_valid( io_scr_resp_valid ),
       .io_smi_resp_bits( io_scr_resp_bits )
  );
endmodule

module SCRFile(input clk, input reset,
    output io_smi_req_ready,
    input  io_smi_req_valid,
    input  io_smi_req_bits_rw,
    input [5:0] io_smi_req_bits_addr,
    input [63:0] io_smi_req_bits_data,
    input  io_smi_resp_ready,
    output io_smi_resp_valid,
    output[63:0] io_smi_resp_bits,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[63:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T8;
  wire[5:0] T9;
  reg [5:0] read_addr;
  wire[5:0] T135;
  wire[5:0] T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T13;
  wire T14;
  wire[63:0] T15;
  wire[63:0] T16;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T17;
  wire[63:0] T18;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T19;
  wire T20;
  wire T21;
  wire[63:0] T22;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T25;
  wire[63:0] T26;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T27;
  wire T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T31;
  wire[63:0] T32;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T41;
  wire[63:0] T42;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T43;
  wire T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T47;
  wire[63:0] T48;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T49;
  wire T50;
  wire T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T55;
  wire[63:0] T56;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T57;
  wire T58;
  wire[63:0] T59;
  wire[63:0] T60;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T61;
  wire[63:0] T62;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  wire[63:0] T72;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T73;
  wire[63:0] T74;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T75;
  wire T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T79;
  wire[63:0] T80;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T81;
  wire T82;
  wire T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T87;
  wire[63:0] T88;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T89;
  wire T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T93;
  wire[63:0] T94;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[63:0] T99;
  wire[63:0] T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T103;
  wire[63:0] T104;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T105;
  wire T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T109;
  wire[63:0] T110;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T111;
  wire T112;
  wire T113;
  wire[63:0] T114;
  wire[63:0] T115;
  wire[63:0] T116;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T117;
  wire[63:0] T118;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T119;
  wire T120;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T123;
  wire[63:0] T124;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  reg  resp_valid;
  wire T136;
  wire T131;
  wire T132;
  wire T133;
  wire T134;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    read_addr = {1{$random}};
    resp_valid = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_scr_wdata = io_smi_req_bits_data;
  assign io_scr_waddr = io_smi_req_bits_addr;
  assign io_scr_wen = T0;
  assign T0 = T1 & io_smi_req_bits_rw;
  assign T1 = io_smi_req_ready & io_smi_req_valid;
  assign io_smi_resp_bits = T2;
  assign T2 = T130 ? T68 : T3;
  assign T3 = T67 ? T37 : T4;
  assign T4 = T36 ? T22 : T5;
  assign T5 = T21 ? T15 : T6;
  assign T6 = T14 ? T12 : T7;
  assign T7 = T8 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h400;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = read_addr;
  assign T135 = reset ? 6'h0 : T10;
  assign T10 = T11 ? io_smi_req_bits_addr : read_addr;
  assign T11 = io_smi_req_ready & io_smi_req_valid;
  assign T12 = T13 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T13 = T9[1'h0:1'h0];
  assign T14 = T9[1'h1:1'h1];
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign T22 = T35 ? T29 : T23;
  assign T23 = T28 ? T26 : T24;
  assign T24 = T25 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T25 = T9[1'h0:1'h0];
  assign T26 = T27 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T27 = T9[1'h0:1'h0];
  assign T28 = T9[1'h1:1'h1];
  assign T29 = T34 ? T32 : T30;
  assign T30 = T31 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T31 = T9[1'h0:1'h0];
  assign T32 = T33 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T33 = T9[1'h0:1'h0];
  assign T34 = T9[1'h1:1'h1];
  assign T35 = T9[2'h2:2'h2];
  assign T36 = T9[2'h3:2'h3];
  assign T37 = T66 ? T52 : T38;
  assign T38 = T51 ? T45 : T39;
  assign T39 = T44 ? T42 : T40;
  assign T40 = T41 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T41 = T9[1'h0:1'h0];
  assign T42 = T43 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T43 = T9[1'h0:1'h0];
  assign T44 = T9[1'h1:1'h1];
  assign T45 = T50 ? T48 : T46;
  assign T46 = T47 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T47 = T9[1'h0:1'h0];
  assign T48 = T49 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T49 = T9[1'h0:1'h0];
  assign T50 = T9[1'h1:1'h1];
  assign T51 = T9[2'h2:2'h2];
  assign T52 = T65 ? T59 : T53;
  assign T53 = T58 ? T56 : T54;
  assign T54 = T55 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T55 = T9[1'h0:1'h0];
  assign T56 = T57 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T57 = T9[1'h0:1'h0];
  assign T58 = T9[1'h1:1'h1];
  assign T59 = T64 ? T62 : T60;
  assign T60 = T61 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T61 = T9[1'h0:1'h0];
  assign T62 = T63 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T63 = T9[1'h0:1'h0];
  assign T64 = T9[1'h1:1'h1];
  assign T65 = T9[2'h2:2'h2];
  assign T66 = T9[2'h3:2'h3];
  assign T67 = T9[3'h4:3'h4];
  assign T68 = T129 ? T99 : T69;
  assign T69 = T98 ? T84 : T70;
  assign T70 = T83 ? T77 : T71;
  assign T71 = T76 ? T74 : T72;
  assign T72 = T73 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T73 = T9[1'h0:1'h0];
  assign T74 = T75 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T75 = T9[1'h0:1'h0];
  assign T76 = T9[1'h1:1'h1];
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T79 = T9[1'h0:1'h0];
  assign T80 = T81 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T81 = T9[1'h0:1'h0];
  assign T82 = T9[1'h1:1'h1];
  assign T83 = T9[2'h2:2'h2];
  assign T84 = T97 ? T91 : T85;
  assign T85 = T90 ? T88 : T86;
  assign T86 = T87 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T87 = T9[1'h0:1'h0];
  assign T88 = T89 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T89 = T9[1'h0:1'h0];
  assign T90 = T9[1'h1:1'h1];
  assign T91 = T96 ? T94 : T92;
  assign T92 = T93 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T93 = T9[1'h0:1'h0];
  assign T94 = T95 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T95 = T9[1'h0:1'h0];
  assign T96 = T9[1'h1:1'h1];
  assign T97 = T9[2'h2:2'h2];
  assign T98 = T9[2'h3:2'h3];
  assign T99 = T128 ? T114 : T100;
  assign T100 = T113 ? T107 : T101;
  assign T101 = T106 ? T104 : T102;
  assign T102 = T103 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T103 = T9[1'h0:1'h0];
  assign T104 = T105 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T105 = T9[1'h0:1'h0];
  assign T106 = T9[1'h1:1'h1];
  assign T107 = T112 ? T110 : T108;
  assign T108 = T109 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T109 = T9[1'h0:1'h0];
  assign T110 = T111 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T111 = T9[1'h0:1'h0];
  assign T112 = T9[1'h1:1'h1];
  assign T113 = T9[2'h2:2'h2];
  assign T114 = T127 ? T121 : T115;
  assign T115 = T120 ? T118 : T116;
  assign T116 = T117 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T117 = T9[1'h0:1'h0];
  assign T118 = T119 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T119 = T9[1'h0:1'h0];
  assign T120 = T9[1'h1:1'h1];
  assign T121 = T126 ? T124 : T122;
  assign T122 = T123 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T123 = T9[1'h0:1'h0];
  assign T124 = T125 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T125 = T9[1'h0:1'h0];
  assign T126 = T9[1'h1:1'h1];
  assign T127 = T9[2'h2:2'h2];
  assign T128 = T9[2'h3:2'h3];
  assign T129 = T9[3'h4:3'h4];
  assign T130 = T9[3'h5:3'h5];
  assign io_smi_resp_valid = resp_valid;
  assign T136 = reset ? 1'h0 : T131;
  assign T131 = T133 ? 1'h0 : T132;
  assign T132 = T11 ? 1'h1 : resp_valid;
  assign T133 = io_smi_resp_ready & io_smi_resp_valid;
  assign io_smi_req_ready = T134;
  assign T134 = resp_valid ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      read_addr <= 6'h0;
    end else if(T11) begin
      read_addr <= io_smi_req_bits_addr;
    end
    if(reset) begin
      resp_valid <= 1'h0;
    end else if(T133) begin
      resp_valid <= 1'h0;
    end else if(T11) begin
      resp_valid <= 1'h1;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_addr,
    input [7:0] io_enq_bits_len,
    input [2:0] io_enq_bits_size,
    input [1:0] io_enq_bits_burst,
    input  io_enq_bits_lock,
    input [3:0] io_enq_bits_cache,
    input [2:0] io_enq_bits_prot,
    input [3:0] io_enq_bits_qos,
    input [3:0] io_enq_bits_region,
    input [3:0] io_enq_bits_id,
    input  io_enq_bits_user,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_addr,
    output[7:0] io_deq_bits_len,
    output[2:0] io_deq_bits_size,
    output[1:0] io_deq_bits_burst,
    output io_deq_bits_lock,
    output[3:0] io_deq_bits_cache,
    output[2:0] io_deq_bits_prot,
    output[3:0] io_deq_bits_qos,
    output[3:0] io_deq_bits_region,
    output[3:0] io_deq_bits_id,
    output io_deq_bits_user,
    output io_count
);

  wire T29;
  wire[1:0] T0;
  reg  full;
  wire T30;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire T3;
  wire[65:0] T4;
  reg [65:0] ram [0:0];
  wire[65:0] T5;
  wire[65:0] T6;
  wire[65:0] T7;
  wire[19:0] T8;
  wire[8:0] T9;
  wire[4:0] T10;
  wire[10:0] T11;
  wire[6:0] T12;
  wire[45:0] T13;
  wire[5:0] T14;
  wire[2:0] T15;
  wire[39:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[2:0] T20;
  wire[3:0] T21;
  wire T22;
  wire[1:0] T23;
  wire[2:0] T24;
  wire[7:0] T25;
  wire[31:0] T26;
  wire T27;
  wire empty;
  wire T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T29;
  assign T29 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T30 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_user = T3;
  assign T3 = T4[1'h0:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {T13, T8};
  assign T8 = {T11, T9};
  assign T9 = {io_enq_bits_region, T10};
  assign T10 = {io_enq_bits_id, io_enq_bits_user};
  assign T11 = {io_enq_bits_cache, T12};
  assign T12 = {io_enq_bits_prot, io_enq_bits_qos};
  assign T13 = {T16, T14};
  assign T14 = {io_enq_bits_size, T15};
  assign T15 = {io_enq_bits_burst, io_enq_bits_lock};
  assign T16 = {io_enq_bits_addr, io_enq_bits_len};
  assign io_deq_bits_id = T17;
  assign T17 = T4[3'h4:1'h1];
  assign io_deq_bits_region = T18;
  assign T18 = T4[4'h8:3'h5];
  assign io_deq_bits_qos = T19;
  assign T19 = T4[4'hc:4'h9];
  assign io_deq_bits_prot = T20;
  assign T20 = T4[4'hf:4'hd];
  assign io_deq_bits_cache = T21;
  assign T21 = T4[5'h13:5'h10];
  assign io_deq_bits_lock = T22;
  assign T22 = T4[5'h14:5'h14];
  assign io_deq_bits_burst = T23;
  assign T23 = T4[5'h16:5'h15];
  assign io_deq_bits_size = T24;
  assign T24 = T4[5'h19:5'h17];
  assign io_deq_bits_len = T25;
  assign T25 = T4[6'h21:5'h1a];
  assign io_deq_bits_addr = T26;
  assign T26 = T4[7'h41:6'h22];
  assign io_deq_valid = T27;
  assign T27 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module NastiROM(input clk, input reset,
    output io_aw_ready,
    input  io_aw_valid,
    input [31:0] io_aw_bits_addr,
    input [7:0] io_aw_bits_len,
    input [2:0] io_aw_bits_size,
    input [1:0] io_aw_bits_burst,
    input  io_aw_bits_lock,
    input [3:0] io_aw_bits_cache,
    input [2:0] io_aw_bits_prot,
    input [3:0] io_aw_bits_qos,
    input [3:0] io_aw_bits_region,
    input [3:0] io_aw_bits_id,
    input  io_aw_bits_user,
    output io_w_ready,
    input  io_w_valid,
    input [63:0] io_w_bits_data,
    input  io_w_bits_last,
    input [7:0] io_w_bits_strb,
    input  io_w_bits_user,
    input  io_b_ready,
    output io_b_valid,
    //output[1:0] io_b_bits_resp
    //output[3:0] io_b_bits_id
    //output io_b_bits_user
    output io_ar_ready,
    input  io_ar_valid,
    input [31:0] io_ar_bits_addr,
    input [7:0] io_ar_bits_len,
    input [2:0] io_ar_bits_size,
    input [1:0] io_ar_bits_burst,
    input  io_ar_bits_lock,
    input [3:0] io_ar_bits_cache,
    input [2:0] io_ar_bits_prot,
    input [3:0] io_ar_bits_qos,
    input [3:0] io_ar_bits_region,
    input [3:0] io_ar_bits_id,
    input  io_ar_bits_user,
    input  io_r_ready,
    output io_r_valid,
    output[1:0] io_r_bits_resp,
    output[63:0] io_r_bits_data,
    output io_r_bits_last,
    output[3:0] io_r_bits_id,
    output io_r_bits_user
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg[0:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire[3:0] T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] rdata;
  wire[7:0] T13;
  wire[7:0] T14;
  wire[63:0] T15;
  wire[15:0] T16;
  wire[15:0] T17;
  wire[63:0] T18;
  wire[31:0] T19;
  wire[31:0] T20;
  reg [63:0] rdata_word;
  wire[6:0] T22;
  wire[31:0] T23;
  wire T24;
  wire[31:0] T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[31:0] T52;
  wire T28;
  wire T29;
  wire T30;
  wire[3:0] T31;
  wire[3:0] T32;
  wire T33;
  wire[1:0] T34;
  wire[15:0] T35;
  wire T36;
  wire[47:0] T37;
  wire[47:0] T38;
  wire[47:0] T39;
  wire[47:0] T53;
  wire T40;
  wire T41;
  wire T42;
  wire[7:0] T43;
  wire T44;
  wire[55:0] T45;
  wire[55:0] T46;
  wire[55:0] T47;
  wire[55:0] T54;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire[31:0] Queue_io_deq_bits_addr;
  wire[7:0] Queue_io_deq_bits_len;
  wire[2:0] Queue_io_deq_bits_size;
  wire[3:0] Queue_io_deq_bits_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T4 = 1'b0;
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_b_bits_user = {1{$random}};
//  assign io_b_bits_id = {1{$random}};
//  assign io_b_bits_resp = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = io_aw_valid | io_w_valid;
  assign T5 = T6 | reset;
  assign T6 = T8 | T7;
  assign T7 = Queue_io_deq_bits_len == 8'h0;
  assign T8 = Queue_io_deq_valid ^ 1'h1;
  assign io_r_bits_user = T9;
  assign T9 = 1'h0;
  assign io_r_bits_id = T10;
  assign T10 = Queue_io_deq_bits_id;
  assign io_r_bits_last = T11;
  assign T11 = 1'h1;
  assign io_r_bits_data = T12;
  assign T12 = rdata;
  assign rdata = {T45, T13};
  assign T13 = T44 ? T43 : T14;
  assign T14 = T15[3'h7:1'h0];
  assign T15 = {T37, T16};
  assign T16 = T36 ? T35 : T17;
  assign T17 = T18[4'hf:1'h0];
  assign T18 = {T25, T19};
  assign T19 = T24 ? T23 : T20;
  assign T20 = rdata_word[5'h1f:1'h0];
  always @(*) case (T22)
    0: rdata_word = 64'hb020000edfe0dd0;
    1: rdata_word = 64'hc001000038000000;
    2: rdata_word = 64'h1100000028000000;
    3: rdata_word = 64'h10000000;
    4: rdata_word = 64'h880100004b000000;
    5: rdata_word = 64'h0;
    6: rdata_word = 64'h0;
    7: rdata_word = 64'h1000000;
    8: rdata_word = 64'h400000003000000;
    9: rdata_word = 64'h200000000000000;
    10: rdata_word = 64'h400000003000000;
    11: rdata_word = 64'h20000000f000000;
    12: rdata_word = 64'hc00000003000000;
    13: rdata_word = 64'h6b636f521b000000;
    14: rdata_word = 64'h706968432d7465;
    15: rdata_word = 64'h6f6d656d01000000;
    16: rdata_word = 64'h30407972;
    17: rdata_word = 64'h700000003000000;
    18: rdata_word = 64'h6f6d656d21000000;
    19: rdata_word = 64'h300000000007972;
    20: rdata_word = 64'h2d00000010000000;
    21: rdata_word = 64'h0;
    22: rdata_word = 64'h4000000000;
    23: rdata_word = 64'h100000002000000;
    24: rdata_word = 64'h73757063;
    25: rdata_word = 64'h400000003000000;
    26: rdata_word = 64'h200000000000000;
    27: rdata_word = 64'h400000003000000;
    28: rdata_word = 64'h20000000f000000;
    29: rdata_word = 64'h4075706301000000;
    30: rdata_word = 64'h3030303830303034;
    31: rdata_word = 64'h300000000000000;
    32: rdata_word = 64'h2100000004000000;
    33: rdata_word = 64'h300000000757063;
    34: rdata_word = 64'h3100000006000000;
    35: rdata_word = 64'h7663736972;
    36: rdata_word = 64'h500000003000000;
    37: rdata_word = 64'h343676723c000000;
    38: rdata_word = 64'h300000000000000;
    39: rdata_word = 64'h2d00000008000000;
    40: rdata_word = 64'h80004000000000;
    41: rdata_word = 64'h200000002000000;
    42: rdata_word = 64'h4072637301000000;
    43: rdata_word = 64'h3030303031303034;
    44: rdata_word = 64'h300000000000000;
    45: rdata_word = 64'h2100000004000000;
    46: rdata_word = 64'h300000000726373;
    47: rdata_word = 64'h3100000006000000;
    48: rdata_word = 64'h7663736972;
    49: rdata_word = 64'h400000003000000;
    50: rdata_word = 64'h300000040000000;
    51: rdata_word = 64'h1000000003000000;
    52: rdata_word = 64'h2d000000;
    53: rdata_word = 64'h140;
    54: rdata_word = 64'h200000000020000;
    55: rdata_word = 64'h900000002000000;
    56: rdata_word = 64'h7373657264646123;
    57: rdata_word = 64'h2300736c6c65632d;
    58: rdata_word = 64'h6c65632d657a6973;
    59: rdata_word = 64'h6c65646f6d00736c;
    60: rdata_word = 64'h5f65636976656400;
    61: rdata_word = 64'h6765720065707974;
    62: rdata_word = 64'h697461706d6f6300;
    63: rdata_word = 64'h61736900656c62;
    64: rdata_word = 64'h69746365746f7270;
    65: rdata_word = 64'h6e6f;
    66: rdata_word = 64'h0;
    default: begin
      rdata_word = 64'bx;
`ifndef SYNTHESIS
// synthesis translate_off
      rdata_word = {2{$random}};
// synthesis translate_on
`endif
    end
  endcase
  assign T22 = Queue_io_deq_bits_addr[4'h9:2'h3];
  assign T23 = rdata_word[6'h3f:6'h20];
  assign T24 = Queue_io_deq_bits_addr[2'h2:2'h2];
  assign T25 = T33 ? T27 : T26;
  assign T26 = rdata_word[6'h3f:6'h20];
  assign T27 = 32'h0 - T52;
  assign T52 = {31'h0, T28};
  assign T28 = T30 & T29;
  assign T29 = T19[5'h1f:5'h1f];
  assign T30 = $signed(1'h0) <= $signed(T31);
  assign T31 = T32;
  assign T32 = {1'h1, Queue_io_deq_bits_size};
  assign T33 = T34 == 2'h2;
  assign T34 = T32[1'h1:1'h0];
  assign T35 = T18[5'h1f:5'h10];
  assign T36 = Queue_io_deq_bits_addr[1'h1:1'h1];
  assign T37 = T42 ? T39 : T38;
  assign T38 = T18[6'h3f:5'h10];
  assign T39 = 48'h0 - T53;
  assign T53 = {47'h0, T40};
  assign T40 = T30 & T41;
  assign T41 = T16[4'hf:4'hf];
  assign T42 = T34 == 2'h1;
  assign T43 = T15[4'hf:4'h8];
  assign T44 = Queue_io_deq_bits_addr[1'h0:1'h0];
  assign T45 = T50 ? T47 : T46;
  assign T46 = T15[6'h3f:4'h8];
  assign T47 = 56'h0 - T54;
  assign T54 = {55'h0, T48};
  assign T48 = T30 & T49;
  assign T49 = T13[3'h7:3'h7];
  assign T50 = T34 == 2'h0;
  assign io_r_bits_resp = T51;
  assign T51 = 2'h0;
  assign io_r_valid = Queue_io_deq_valid;
  assign io_ar_ready = Queue_io_enq_ready;
  assign io_b_valid = 1'h0;
  assign io_w_ready = 1'h0;
  assign io_aw_ready = 1'h0;
  Queue_7 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( io_ar_valid ),
       .io_enq_bits_addr( io_ar_bits_addr ),
       .io_enq_bits_len( io_ar_bits_len ),
       .io_enq_bits_size( io_ar_bits_size ),
       .io_enq_bits_burst( io_ar_bits_burst ),
       .io_enq_bits_lock( io_ar_bits_lock ),
       .io_enq_bits_cache( io_ar_bits_cache ),
       .io_enq_bits_prot( io_ar_bits_prot ),
       .io_enq_bits_qos( io_ar_bits_qos ),
       .io_enq_bits_region( io_ar_bits_region ),
       .io_enq_bits_id( io_ar_bits_id ),
       .io_enq_bits_user( io_ar_bits_user ),
       .io_deq_ready( io_r_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_io_deq_bits_len ),
       .io_deq_bits_size( Queue_io_deq_bits_size ),
       //.io_deq_bits_burst(  )
       //.io_deq_bits_lock(  )
       //.io_deq_bits_cache(  )
       //.io_deq_bits_prot(  )
       //.io_deq_bits_qos(  )
       //.io_deq_bits_region(  )
       .io_deq_bits_id( Queue_io_deq_bits_id )
       //.io_deq_bits_user(  )
       //.io_count(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T4 <= 1'b1;
  if(!T5 && T4 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't burst-read from NastiROM");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "Can't write to NastiROM");
    $finish;
  end
// synthesis translate_on
`endif
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[3:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [3:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[3:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [3:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user,
    output io_tiles_cached_0_acquire_ready,
    input  io_tiles_cached_0_acquire_valid,
    input [25:0] io_tiles_cached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_cached_0_acquire_bits_addr_beat,
    input  io_tiles_cached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_cached_0_acquire_bits_a_type,
    input [16:0] io_tiles_cached_0_acquire_bits_union,
    input [127:0] io_tiles_cached_0_acquire_bits_data,
    input  io_tiles_cached_0_grant_ready,
    output io_tiles_cached_0_grant_valid,
    output[1:0] io_tiles_cached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_cached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
    output io_tiles_cached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_cached_0_grant_bits_g_type,
    output[127:0] io_tiles_cached_0_grant_bits_data,
    input  io_tiles_cached_0_probe_ready,
    output io_tiles_cached_0_probe_valid,
    output[25:0] io_tiles_cached_0_probe_bits_addr_block,
    output[1:0] io_tiles_cached_0_probe_bits_p_type,
    output io_tiles_cached_0_release_ready,
    input  io_tiles_cached_0_release_valid,
    input [1:0] io_tiles_cached_0_release_bits_addr_beat,
    input [25:0] io_tiles_cached_0_release_bits_addr_block,
    input [1:0] io_tiles_cached_0_release_bits_client_xact_id,
    input  io_tiles_cached_0_release_bits_voluntary,
    input [2:0] io_tiles_cached_0_release_bits_r_type,
    input [127:0] io_tiles_cached_0_release_bits_data,
    output io_tiles_uncached_0_acquire_ready,
    input  io_tiles_uncached_0_acquire_valid,
    input [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
    input [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
    input [1:0] io_tiles_uncached_0_acquire_bits_addr_beat,
    input  io_tiles_uncached_0_acquire_bits_is_builtin_type,
    input [2:0] io_tiles_uncached_0_acquire_bits_a_type,
    input [16:0] io_tiles_uncached_0_acquire_bits_union,
    input [127:0] io_tiles_uncached_0_acquire_bits_data,
    input  io_tiles_uncached_0_grant_ready,
    output io_tiles_uncached_0_grant_valid,
    output[1:0] io_tiles_uncached_0_grant_bits_addr_beat,
    output[1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
    output[2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
    output io_tiles_uncached_0_grant_bits_is_builtin_type,
    output[3:0] io_tiles_uncached_0_grant_bits_g_type,
    output[127:0] io_tiles_uncached_0_grant_bits_data,
    output io_htif_0_reset,
    output io_htif_0_id,
    input  io_htif_0_csr_req_ready,
    output io_htif_0_csr_req_valid,
    output io_htif_0_csr_req_bits_rw,
    output[11:0] io_htif_0_csr_req_bits_addr,
    output[63:0] io_htif_0_csr_req_bits_data,
    output io_htif_0_csr_resp_ready,
    input  io_htif_0_csr_resp_valid,
    input [63:0] io_htif_0_csr_resp_bits,
    input  io_htif_0_debug_stats_csr,
    //input  io_mem_backup_ctrl_en
    //input  io_mem_backup_ctrl_in_valid
    //input  io_mem_backup_ctrl_out_ready
    //output io_mem_backup_ctrl_out_valid
    input  io_mmio_aw_ready,
    output io_mmio_aw_valid,
    output[31:0] io_mmio_aw_bits_addr,
    output[7:0] io_mmio_aw_bits_len,
    output[2:0] io_mmio_aw_bits_size,
    output[1:0] io_mmio_aw_bits_burst,
    output io_mmio_aw_bits_lock,
    output[3:0] io_mmio_aw_bits_cache,
    output[2:0] io_mmio_aw_bits_prot,
    output[3:0] io_mmio_aw_bits_qos,
    output[3:0] io_mmio_aw_bits_region,
    output[3:0] io_mmio_aw_bits_id,
    output io_mmio_aw_bits_user,
    input  io_mmio_w_ready,
    output io_mmio_w_valid,
    output[63:0] io_mmio_w_bits_data,
    output io_mmio_w_bits_last,
    output[7:0] io_mmio_w_bits_strb,
    output io_mmio_w_bits_user,
    output io_mmio_b_ready,
    input  io_mmio_b_valid,
    input [1:0] io_mmio_b_bits_resp,
    input [3:0] io_mmio_b_bits_id,
    input  io_mmio_b_bits_user,
    input  io_mmio_ar_ready,
    output io_mmio_ar_valid,
    output[31:0] io_mmio_ar_bits_addr,
    output[7:0] io_mmio_ar_bits_len,
    output[2:0] io_mmio_ar_bits_size,
    output[1:0] io_mmio_ar_bits_burst,
    output io_mmio_ar_bits_lock,
    output[3:0] io_mmio_ar_bits_cache,
    output[2:0] io_mmio_ar_bits_prot,
    output[3:0] io_mmio_ar_bits_qos,
    output[3:0] io_mmio_ar_bits_region,
    output[3:0] io_mmio_ar_bits_id,
    output io_mmio_ar_bits_user,
    output io_mmio_r_ready,
    input  io_mmio_r_valid,
    input [1:0] io_mmio_r_bits_resp,
    input [63:0] io_mmio_r_bits_data,
    input  io_mmio_r_bits_last,
    input [3:0] io_mmio_r_bits_id,
    input  io_mmio_r_bits_user
    //output io_dma_0_req_ready
    //input  io_dma_0_req_valid
    //input [1:0] io_dma_0_req_bits_client_xact_id
    //input [1:0] io_dma_0_req_bits_cmd
    //input [31:0] io_dma_0_req_bits_source
    //input [31:0] io_dma_0_req_bits_dest
    //input [31:0] io_dma_0_req_bits_length
    //input  io_dma_0_resp_ready
    //output io_dma_0_resp_valid
    //output[1:0] io_dma_0_resp_bits_client_xact_id
    //output[1:0] io_dma_0_resp_bits_status
);

  wire htif_io_host_in_ready;
  wire htif_io_host_out_valid;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_debug_stats_csr;
  wire htif_io_cpu_0_reset;
  wire htif_io_cpu_0_id;
  wire htif_io_cpu_0_csr_req_valid;
  wire htif_io_cpu_0_csr_req_bits_rw;
  wire[11:0] htif_io_cpu_0_csr_req_bits_addr;
  wire[63:0] htif_io_cpu_0_csr_req_bits_data;
  wire htif_io_cpu_0_csr_resp_ready;
  wire htif_io_mem_acquire_valid;
  wire[25:0] htif_io_mem_acquire_bits_addr_block;
  wire[1:0] htif_io_mem_acquire_bits_client_xact_id;
  wire[1:0] htif_io_mem_acquire_bits_addr_beat;
  wire htif_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] htif_io_mem_acquire_bits_a_type;
  wire[16:0] htif_io_mem_acquire_bits_union;
  wire[127:0] htif_io_mem_acquire_bits_data;
  wire htif_io_mem_grant_ready;
  wire htif_io_scr_req_valid;
  wire htif_io_scr_req_bits_rw;
  wire[5:0] htif_io_scr_req_bits_addr;
  wire[63:0] htif_io_scr_req_bits_data;
  wire htif_io_scr_resp_ready;
  wire scrFile_io_smi_req_ready;
  wire scrFile_io_smi_resp_valid;
  wire[63:0] scrFile_io_smi_resp_bits;
  wire SMIArbiter_io_in_1_req_ready;
  wire SMIArbiter_io_in_1_resp_valid;
  wire[63:0] SMIArbiter_io_in_1_resp_bits;
  wire SMIArbiter_io_in_0_req_ready;
  wire SMIArbiter_io_in_0_resp_valid;
  wire[63:0] SMIArbiter_io_in_0_resp_bits;
  wire SMIArbiter_io_out_req_valid;
  wire SMIArbiter_io_out_req_bits_rw;
  wire[11:0] SMIArbiter_io_out_req_bits_addr;
  wire[63:0] SMIArbiter_io_out_req_bits_data;
  wire SMIArbiter_io_out_resp_ready;
  wire scrArb_io_in_1_req_ready;
  wire scrArb_io_in_1_resp_valid;
  wire[63:0] scrArb_io_in_1_resp_bits;
  wire scrArb_io_in_0_req_ready;
  wire scrArb_io_in_0_resp_valid;
  wire[63:0] scrArb_io_in_0_resp_bits;
  wire scrArb_io_out_req_valid;
  wire scrArb_io_out_req_bits_rw;
  wire[5:0] scrArb_io_out_req_bits_addr;
  wire[63:0] scrArb_io_out_req_bits_data;
  wire scrArb_io_out_resp_ready;
  wire deviceTree_io_aw_ready;
  wire deviceTree_io_w_ready;
  wire deviceTree_io_b_valid;
  wire deviceTree_io_ar_ready;
  wire deviceTree_io_r_valid;
  wire[1:0] deviceTree_io_r_bits_resp;
  wire[63:0] deviceTree_io_r_bits_data;
  wire deviceTree_io_r_bits_last;
  wire[3:0] deviceTree_io_r_bits_id;
  wire deviceTree_io_r_bits_user;
  wire outmemsys_io_tiles_cached_0_acquire_ready;
  wire outmemsys_io_tiles_cached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire outmemsys_io_tiles_cached_0_probe_valid;
  wire[25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire outmemsys_io_tiles_cached_0_release_ready;
  wire outmemsys_io_tiles_uncached_0_acquire_ready;
  wire outmemsys_io_tiles_uncached_0_grant_valid;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire outmemsys_io_htif_uncached_acquire_ready;
  wire outmemsys_io_htif_uncached_grant_valid;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_addr_beat;
  wire[1:0] outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  wire[2:0] outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  wire outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  wire[3:0] outmemsys_io_htif_uncached_grant_bits_g_type;
  wire[127:0] outmemsys_io_htif_uncached_grant_bits_data;
  wire outmemsys_io_mem_0_aw_valid;
  wire[31:0] outmemsys_io_mem_0_aw_bits_addr;
  wire[7:0] outmemsys_io_mem_0_aw_bits_len;
  wire[2:0] outmemsys_io_mem_0_aw_bits_size;
  wire[1:0] outmemsys_io_mem_0_aw_bits_burst;
  wire outmemsys_io_mem_0_aw_bits_lock;
  wire[3:0] outmemsys_io_mem_0_aw_bits_cache;
  wire[2:0] outmemsys_io_mem_0_aw_bits_prot;
  wire[3:0] outmemsys_io_mem_0_aw_bits_qos;
  wire[3:0] outmemsys_io_mem_0_aw_bits_region;
  wire[3:0] outmemsys_io_mem_0_aw_bits_id;
  wire outmemsys_io_mem_0_aw_bits_user;
  wire outmemsys_io_mem_0_w_valid;
  wire[63:0] outmemsys_io_mem_0_w_bits_data;
  wire outmemsys_io_mem_0_w_bits_last;
  wire[7:0] outmemsys_io_mem_0_w_bits_strb;
  wire outmemsys_io_mem_0_w_bits_user;
  wire outmemsys_io_mem_0_b_ready;
  wire outmemsys_io_mem_0_ar_valid;
  wire[31:0] outmemsys_io_mem_0_ar_bits_addr;
  wire[7:0] outmemsys_io_mem_0_ar_bits_len;
  wire[2:0] outmemsys_io_mem_0_ar_bits_size;
  wire[1:0] outmemsys_io_mem_0_ar_bits_burst;
  wire outmemsys_io_mem_0_ar_bits_lock;
  wire[3:0] outmemsys_io_mem_0_ar_bits_cache;
  wire[2:0] outmemsys_io_mem_0_ar_bits_prot;
  wire[3:0] outmemsys_io_mem_0_ar_bits_qos;
  wire[3:0] outmemsys_io_mem_0_ar_bits_region;
  wire[3:0] outmemsys_io_mem_0_ar_bits_id;
  wire outmemsys_io_mem_0_ar_bits_user;
  wire outmemsys_io_mem_0_r_ready;
  wire outmemsys_io_csr_0_req_valid;
  wire outmemsys_io_csr_0_req_bits_rw;
  wire[11:0] outmemsys_io_csr_0_req_bits_addr;
  wire[63:0] outmemsys_io_csr_0_req_bits_data;
  wire outmemsys_io_csr_0_resp_ready;
  wire outmemsys_io_scr_req_valid;
  wire outmemsys_io_scr_req_bits_rw;
  wire[5:0] outmemsys_io_scr_req_bits_addr;
  wire[63:0] outmemsys_io_scr_req_bits_data;
  wire outmemsys_io_scr_resp_ready;
  wire outmemsys_io_mmio_aw_valid;
  wire[31:0] outmemsys_io_mmio_aw_bits_addr;
  wire[7:0] outmemsys_io_mmio_aw_bits_len;
  wire[2:0] outmemsys_io_mmio_aw_bits_size;
  wire[1:0] outmemsys_io_mmio_aw_bits_burst;
  wire outmemsys_io_mmio_aw_bits_lock;
  wire[3:0] outmemsys_io_mmio_aw_bits_cache;
  wire[2:0] outmemsys_io_mmio_aw_bits_prot;
  wire[3:0] outmemsys_io_mmio_aw_bits_qos;
  wire[3:0] outmemsys_io_mmio_aw_bits_region;
  wire[3:0] outmemsys_io_mmio_aw_bits_id;
  wire outmemsys_io_mmio_aw_bits_user;
  wire outmemsys_io_mmio_w_valid;
  wire[63:0] outmemsys_io_mmio_w_bits_data;
  wire outmemsys_io_mmio_w_bits_last;
  wire[7:0] outmemsys_io_mmio_w_bits_strb;
  wire outmemsys_io_mmio_w_bits_user;
  wire outmemsys_io_mmio_b_ready;
  wire outmemsys_io_mmio_ar_valid;
  wire[31:0] outmemsys_io_mmio_ar_bits_addr;
  wire[7:0] outmemsys_io_mmio_ar_bits_len;
  wire[2:0] outmemsys_io_mmio_ar_bits_size;
  wire[1:0] outmemsys_io_mmio_ar_bits_burst;
  wire outmemsys_io_mmio_ar_bits_lock;
  wire[3:0] outmemsys_io_mmio_ar_bits_cache;
  wire[2:0] outmemsys_io_mmio_ar_bits_prot;
  wire[3:0] outmemsys_io_mmio_ar_bits_qos;
  wire[3:0] outmemsys_io_mmio_ar_bits_region;
  wire[3:0] outmemsys_io_mmio_ar_bits_id;
  wire outmemsys_io_mmio_ar_bits_user;
  wire outmemsys_io_mmio_r_ready;
  wire outmemsys_io_deviceTree_aw_valid;
  wire[31:0] outmemsys_io_deviceTree_aw_bits_addr;
  wire[7:0] outmemsys_io_deviceTree_aw_bits_len;
  wire[2:0] outmemsys_io_deviceTree_aw_bits_size;
  wire[1:0] outmemsys_io_deviceTree_aw_bits_burst;
  wire outmemsys_io_deviceTree_aw_bits_lock;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_cache;
  wire[2:0] outmemsys_io_deviceTree_aw_bits_prot;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_qos;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_region;
  wire[3:0] outmemsys_io_deviceTree_aw_bits_id;
  wire outmemsys_io_deviceTree_aw_bits_user;
  wire outmemsys_io_deviceTree_w_valid;
  wire[63:0] outmemsys_io_deviceTree_w_bits_data;
  wire outmemsys_io_deviceTree_w_bits_last;
  wire[7:0] outmemsys_io_deviceTree_w_bits_strb;
  wire outmemsys_io_deviceTree_w_bits_user;
  wire outmemsys_io_deviceTree_b_ready;
  wire outmemsys_io_deviceTree_ar_valid;
  wire[31:0] outmemsys_io_deviceTree_ar_bits_addr;
  wire[7:0] outmemsys_io_deviceTree_ar_bits_len;
  wire[2:0] outmemsys_io_deviceTree_ar_bits_size;
  wire[1:0] outmemsys_io_deviceTree_ar_bits_burst;
  wire outmemsys_io_deviceTree_ar_bits_lock;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_cache;
  wire[2:0] outmemsys_io_deviceTree_ar_bits_prot;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_qos;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_region;
  wire[3:0] outmemsys_io_deviceTree_ar_bits_id;
  wire outmemsys_io_deviceTree_ar_bits_user;
  wire outmemsys_io_deviceTree_r_ready;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_dma_0_resp_bits_status = {1{$random}};
//  assign io_dma_0_resp_bits_client_xact_id = {1{$random}};
//  assign io_dma_0_resp_valid = {1{$random}};
//  assign io_dma_0_req_ready = {1{$random}};
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_mmio_r_ready = outmemsys_io_mmio_r_ready;
  assign io_mmio_ar_bits_user = outmemsys_io_mmio_ar_bits_user;
  assign io_mmio_ar_bits_id = outmemsys_io_mmio_ar_bits_id;
  assign io_mmio_ar_bits_region = outmemsys_io_mmio_ar_bits_region;
  assign io_mmio_ar_bits_qos = outmemsys_io_mmio_ar_bits_qos;
  assign io_mmio_ar_bits_prot = outmemsys_io_mmio_ar_bits_prot;
  assign io_mmio_ar_bits_cache = outmemsys_io_mmio_ar_bits_cache;
  assign io_mmio_ar_bits_lock = outmemsys_io_mmio_ar_bits_lock;
  assign io_mmio_ar_bits_burst = outmemsys_io_mmio_ar_bits_burst;
  assign io_mmio_ar_bits_size = outmemsys_io_mmio_ar_bits_size;
  assign io_mmio_ar_bits_len = outmemsys_io_mmio_ar_bits_len;
  assign io_mmio_ar_bits_addr = outmemsys_io_mmio_ar_bits_addr;
  assign io_mmio_ar_valid = outmemsys_io_mmio_ar_valid;
  assign io_mmio_b_ready = outmemsys_io_mmio_b_ready;
  assign io_mmio_w_bits_user = outmemsys_io_mmio_w_bits_user;
  assign io_mmio_w_bits_strb = outmemsys_io_mmio_w_bits_strb;
  assign io_mmio_w_bits_last = outmemsys_io_mmio_w_bits_last;
  assign io_mmio_w_bits_data = outmemsys_io_mmio_w_bits_data;
  assign io_mmio_w_valid = outmemsys_io_mmio_w_valid;
  assign io_mmio_aw_bits_user = outmemsys_io_mmio_aw_bits_user;
  assign io_mmio_aw_bits_id = outmemsys_io_mmio_aw_bits_id;
  assign io_mmio_aw_bits_region = outmemsys_io_mmio_aw_bits_region;
  assign io_mmio_aw_bits_qos = outmemsys_io_mmio_aw_bits_qos;
  assign io_mmio_aw_bits_prot = outmemsys_io_mmio_aw_bits_prot;
  assign io_mmio_aw_bits_cache = outmemsys_io_mmio_aw_bits_cache;
  assign io_mmio_aw_bits_lock = outmemsys_io_mmio_aw_bits_lock;
  assign io_mmio_aw_bits_burst = outmemsys_io_mmio_aw_bits_burst;
  assign io_mmio_aw_bits_size = outmemsys_io_mmio_aw_bits_size;
  assign io_mmio_aw_bits_len = outmemsys_io_mmio_aw_bits_len;
  assign io_mmio_aw_bits_addr = outmemsys_io_mmio_aw_bits_addr;
  assign io_mmio_aw_valid = outmemsys_io_mmio_aw_valid;
  assign io_htif_0_csr_resp_ready = SMIArbiter_io_out_resp_ready;
  assign io_htif_0_csr_req_bits_data = SMIArbiter_io_out_req_bits_data;
  assign io_htif_0_csr_req_bits_addr = SMIArbiter_io_out_req_bits_addr;
  assign io_htif_0_csr_req_bits_rw = SMIArbiter_io_out_req_bits_rw;
  assign io_htif_0_csr_req_valid = SMIArbiter_io_out_req_valid;
  assign io_htif_0_id = htif_io_cpu_0_id;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_mem_0_r_ready = outmemsys_io_mem_0_r_ready;
  assign io_mem_0_ar_bits_user = outmemsys_io_mem_0_ar_bits_user;
  assign io_mem_0_ar_bits_id = outmemsys_io_mem_0_ar_bits_id;
  assign io_mem_0_ar_bits_region = outmemsys_io_mem_0_ar_bits_region;
  assign io_mem_0_ar_bits_qos = outmemsys_io_mem_0_ar_bits_qos;
  assign io_mem_0_ar_bits_prot = outmemsys_io_mem_0_ar_bits_prot;
  assign io_mem_0_ar_bits_cache = outmemsys_io_mem_0_ar_bits_cache;
  assign io_mem_0_ar_bits_lock = outmemsys_io_mem_0_ar_bits_lock;
  assign io_mem_0_ar_bits_burst = outmemsys_io_mem_0_ar_bits_burst;
  assign io_mem_0_ar_bits_size = outmemsys_io_mem_0_ar_bits_size;
  assign io_mem_0_ar_bits_len = outmemsys_io_mem_0_ar_bits_len;
  assign io_mem_0_ar_bits_addr = outmemsys_io_mem_0_ar_bits_addr;
  assign io_mem_0_ar_valid = outmemsys_io_mem_0_ar_valid;
  assign io_mem_0_b_ready = outmemsys_io_mem_0_b_ready;
  assign io_mem_0_w_bits_user = outmemsys_io_mem_0_w_bits_user;
  assign io_mem_0_w_bits_strb = outmemsys_io_mem_0_w_bits_strb;
  assign io_mem_0_w_bits_last = outmemsys_io_mem_0_w_bits_last;
  assign io_mem_0_w_bits_data = outmemsys_io_mem_0_w_bits_data;
  assign io_mem_0_w_valid = outmemsys_io_mem_0_w_valid;
  assign io_mem_0_aw_bits_user = outmemsys_io_mem_0_aw_bits_user;
  assign io_mem_0_aw_bits_id = outmemsys_io_mem_0_aw_bits_id;
  assign io_mem_0_aw_bits_region = outmemsys_io_mem_0_aw_bits_region;
  assign io_mem_0_aw_bits_qos = outmemsys_io_mem_0_aw_bits_qos;
  assign io_mem_0_aw_bits_prot = outmemsys_io_mem_0_aw_bits_prot;
  assign io_mem_0_aw_bits_cache = outmemsys_io_mem_0_aw_bits_cache;
  assign io_mem_0_aw_bits_lock = outmemsys_io_mem_0_aw_bits_lock;
  assign io_mem_0_aw_bits_burst = outmemsys_io_mem_0_aw_bits_burst;
  assign io_mem_0_aw_bits_size = outmemsys_io_mem_0_aw_bits_size;
  assign io_mem_0_aw_bits_len = outmemsys_io_mem_0_aw_bits_len;
  assign io_mem_0_aw_bits_addr = outmemsys_io_mem_0_aw_bits_addr;
  assign io_mem_0_aw_valid = outmemsys_io_mem_0_aw_valid;
  assign io_host_debug_stats_csr = htif_io_host_debug_stats_csr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  Htif htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_csr( htif_io_host_debug_stats_csr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       .io_cpu_0_id( htif_io_cpu_0_id ),
       .io_cpu_0_csr_req_ready( SMIArbiter_io_in_0_req_ready ),
       .io_cpu_0_csr_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_cpu_0_csr_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_cpu_0_csr_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_cpu_0_csr_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_cpu_0_csr_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_cpu_0_csr_resp_valid( SMIArbiter_io_in_0_resp_valid ),
       .io_cpu_0_csr_resp_bits( SMIArbiter_io_in_0_resp_bits ),
       .io_cpu_0_debug_stats_csr( io_htif_0_debug_stats_csr ),
       .io_mem_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_mem_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_mem_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_scr_req_ready( scrArb_io_in_0_req_ready ),
       .io_scr_req_valid( htif_io_scr_req_valid ),
       .io_scr_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( htif_io_scr_req_bits_data ),
       .io_scr_resp_ready( htif_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_0_resp_bits )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign htif.io_cpu_0_id = {1{$random}};
// synthesis translate_on
`endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_cached_0_acquire_ready( outmemsys_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( io_tiles_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( io_tiles_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( io_tiles_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( io_tiles_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( io_tiles_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( io_tiles_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( io_tiles_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( io_tiles_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( io_tiles_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( outmemsys_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( outmemsys_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( outmemsys_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( outmemsys_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( outmemsys_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( io_tiles_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( outmemsys_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( outmemsys_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( outmemsys_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( outmemsys_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( io_tiles_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( io_tiles_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( io_tiles_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( io_tiles_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_voluntary( io_tiles_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_r_type( io_tiles_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_data( io_tiles_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( outmemsys_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( io_tiles_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( io_tiles_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( io_tiles_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( io_tiles_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( io_tiles_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( io_tiles_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( io_tiles_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( io_tiles_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( io_tiles_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( outmemsys_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( outmemsys_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( outmemsys_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( outmemsys_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_uncached_acquire_ready( outmemsys_io_htif_uncached_acquire_ready ),
       .io_htif_uncached_acquire_valid( htif_io_mem_acquire_valid ),
       .io_htif_uncached_acquire_bits_addr_block( htif_io_mem_acquire_bits_addr_block ),
       .io_htif_uncached_acquire_bits_client_xact_id( htif_io_mem_acquire_bits_client_xact_id ),
       .io_htif_uncached_acquire_bits_addr_beat( htif_io_mem_acquire_bits_addr_beat ),
       .io_htif_uncached_acquire_bits_is_builtin_type( htif_io_mem_acquire_bits_is_builtin_type ),
       .io_htif_uncached_acquire_bits_a_type( htif_io_mem_acquire_bits_a_type ),
       .io_htif_uncached_acquire_bits_union( htif_io_mem_acquire_bits_union ),
       .io_htif_uncached_acquire_bits_data( htif_io_mem_acquire_bits_data ),
       .io_htif_uncached_grant_ready( htif_io_mem_grant_ready ),
       .io_htif_uncached_grant_valid( outmemsys_io_htif_uncached_grant_valid ),
       .io_htif_uncached_grant_bits_addr_beat( outmemsys_io_htif_uncached_grant_bits_addr_beat ),
       .io_htif_uncached_grant_bits_client_xact_id( outmemsys_io_htif_uncached_grant_bits_client_xact_id ),
       .io_htif_uncached_grant_bits_manager_xact_id( outmemsys_io_htif_uncached_grant_bits_manager_xact_id ),
       .io_htif_uncached_grant_bits_is_builtin_type( outmemsys_io_htif_uncached_grant_bits_is_builtin_type ),
       .io_htif_uncached_grant_bits_g_type( outmemsys_io_htif_uncached_grant_bits_g_type ),
       .io_htif_uncached_grant_bits_data( outmemsys_io_htif_uncached_grant_bits_data ),
       .io_incoherent_0( htif_io_cpu_0_reset ),
       .io_mem_0_aw_ready( io_mem_0_aw_ready ),
       .io_mem_0_aw_valid( outmemsys_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( outmemsys_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( outmemsys_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( outmemsys_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( outmemsys_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( outmemsys_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( outmemsys_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( outmemsys_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( outmemsys_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( outmemsys_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( outmemsys_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( outmemsys_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( io_mem_0_w_ready ),
       .io_mem_0_w_valid( outmemsys_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( outmemsys_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( outmemsys_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( outmemsys_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( outmemsys_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( outmemsys_io_mem_0_b_ready ),
       .io_mem_0_b_valid( io_mem_0_b_valid ),
       .io_mem_0_b_bits_resp( io_mem_0_b_bits_resp ),
       .io_mem_0_b_bits_id( io_mem_0_b_bits_id ),
       .io_mem_0_b_bits_user( io_mem_0_b_bits_user ),
       .io_mem_0_ar_ready( io_mem_0_ar_ready ),
       .io_mem_0_ar_valid( outmemsys_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( outmemsys_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( outmemsys_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( outmemsys_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( outmemsys_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( outmemsys_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( outmemsys_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( outmemsys_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( outmemsys_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( outmemsys_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( outmemsys_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( outmemsys_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( outmemsys_io_mem_0_r_ready ),
       .io_mem_0_r_valid( io_mem_0_r_valid ),
       .io_mem_0_r_bits_resp( io_mem_0_r_bits_resp ),
       .io_mem_0_r_bits_data( io_mem_0_r_bits_data ),
       .io_mem_0_r_bits_last( io_mem_0_r_bits_last ),
       .io_mem_0_r_bits_id( io_mem_0_r_bits_id ),
       .io_mem_0_r_bits_user( io_mem_0_r_bits_user ),
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
       .io_csr_0_req_ready( SMIArbiter_io_in_1_req_ready ),
       .io_csr_0_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_csr_0_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_csr_0_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_csr_0_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_csr_0_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_csr_0_resp_valid( SMIArbiter_io_in_1_resp_valid ),
       .io_csr_0_resp_bits( SMIArbiter_io_in_1_resp_bits ),
       .io_scr_req_ready( scrArb_io_in_1_req_ready ),
       .io_scr_req_valid( outmemsys_io_scr_req_valid ),
       .io_scr_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_scr_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_scr_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_scr_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_scr_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_scr_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_mmio_aw_ready( io_mmio_aw_ready ),
       .io_mmio_aw_valid( outmemsys_io_mmio_aw_valid ),
       .io_mmio_aw_bits_addr( outmemsys_io_mmio_aw_bits_addr ),
       .io_mmio_aw_bits_len( outmemsys_io_mmio_aw_bits_len ),
       .io_mmio_aw_bits_size( outmemsys_io_mmio_aw_bits_size ),
       .io_mmio_aw_bits_burst( outmemsys_io_mmio_aw_bits_burst ),
       .io_mmio_aw_bits_lock( outmemsys_io_mmio_aw_bits_lock ),
       .io_mmio_aw_bits_cache( outmemsys_io_mmio_aw_bits_cache ),
       .io_mmio_aw_bits_prot( outmemsys_io_mmio_aw_bits_prot ),
       .io_mmio_aw_bits_qos( outmemsys_io_mmio_aw_bits_qos ),
       .io_mmio_aw_bits_region( outmemsys_io_mmio_aw_bits_region ),
       .io_mmio_aw_bits_id( outmemsys_io_mmio_aw_bits_id ),
       .io_mmio_aw_bits_user( outmemsys_io_mmio_aw_bits_user ),
       .io_mmio_w_ready( io_mmio_w_ready ),
       .io_mmio_w_valid( outmemsys_io_mmio_w_valid ),
       .io_mmio_w_bits_data( outmemsys_io_mmio_w_bits_data ),
       .io_mmio_w_bits_last( outmemsys_io_mmio_w_bits_last ),
       .io_mmio_w_bits_strb( outmemsys_io_mmio_w_bits_strb ),
       .io_mmio_w_bits_user( outmemsys_io_mmio_w_bits_user ),
       .io_mmio_b_ready( outmemsys_io_mmio_b_ready ),
       .io_mmio_b_valid( io_mmio_b_valid ),
       .io_mmio_b_bits_resp( io_mmio_b_bits_resp ),
       .io_mmio_b_bits_id( io_mmio_b_bits_id ),
       .io_mmio_b_bits_user( io_mmio_b_bits_user ),
       .io_mmio_ar_ready( io_mmio_ar_ready ),
       .io_mmio_ar_valid( outmemsys_io_mmio_ar_valid ),
       .io_mmio_ar_bits_addr( outmemsys_io_mmio_ar_bits_addr ),
       .io_mmio_ar_bits_len( outmemsys_io_mmio_ar_bits_len ),
       .io_mmio_ar_bits_size( outmemsys_io_mmio_ar_bits_size ),
       .io_mmio_ar_bits_burst( outmemsys_io_mmio_ar_bits_burst ),
       .io_mmio_ar_bits_lock( outmemsys_io_mmio_ar_bits_lock ),
       .io_mmio_ar_bits_cache( outmemsys_io_mmio_ar_bits_cache ),
       .io_mmio_ar_bits_prot( outmemsys_io_mmio_ar_bits_prot ),
       .io_mmio_ar_bits_qos( outmemsys_io_mmio_ar_bits_qos ),
       .io_mmio_ar_bits_region( outmemsys_io_mmio_ar_bits_region ),
       .io_mmio_ar_bits_id( outmemsys_io_mmio_ar_bits_id ),
       .io_mmio_ar_bits_user( outmemsys_io_mmio_ar_bits_user ),
       .io_mmio_r_ready( outmemsys_io_mmio_r_ready ),
       .io_mmio_r_valid( io_mmio_r_valid ),
       .io_mmio_r_bits_resp( io_mmio_r_bits_resp ),
       .io_mmio_r_bits_data( io_mmio_r_bits_data ),
       .io_mmio_r_bits_last( io_mmio_r_bits_last ),
       .io_mmio_r_bits_id( io_mmio_r_bits_id ),
       .io_mmio_r_bits_user( io_mmio_r_bits_user ),
       .io_deviceTree_aw_ready( deviceTree_io_aw_ready ),
       .io_deviceTree_aw_valid( outmemsys_io_deviceTree_aw_valid ),
       .io_deviceTree_aw_bits_addr( outmemsys_io_deviceTree_aw_bits_addr ),
       .io_deviceTree_aw_bits_len( outmemsys_io_deviceTree_aw_bits_len ),
       .io_deviceTree_aw_bits_size( outmemsys_io_deviceTree_aw_bits_size ),
       .io_deviceTree_aw_bits_burst( outmemsys_io_deviceTree_aw_bits_burst ),
       .io_deviceTree_aw_bits_lock( outmemsys_io_deviceTree_aw_bits_lock ),
       .io_deviceTree_aw_bits_cache( outmemsys_io_deviceTree_aw_bits_cache ),
       .io_deviceTree_aw_bits_prot( outmemsys_io_deviceTree_aw_bits_prot ),
       .io_deviceTree_aw_bits_qos( outmemsys_io_deviceTree_aw_bits_qos ),
       .io_deviceTree_aw_bits_region( outmemsys_io_deviceTree_aw_bits_region ),
       .io_deviceTree_aw_bits_id( outmemsys_io_deviceTree_aw_bits_id ),
       .io_deviceTree_aw_bits_user( outmemsys_io_deviceTree_aw_bits_user ),
       .io_deviceTree_w_ready( deviceTree_io_w_ready ),
       .io_deviceTree_w_valid( outmemsys_io_deviceTree_w_valid ),
       .io_deviceTree_w_bits_data( outmemsys_io_deviceTree_w_bits_data ),
       .io_deviceTree_w_bits_last( outmemsys_io_deviceTree_w_bits_last ),
       .io_deviceTree_w_bits_strb( outmemsys_io_deviceTree_w_bits_strb ),
       .io_deviceTree_w_bits_user( outmemsys_io_deviceTree_w_bits_user ),
       .io_deviceTree_b_ready( outmemsys_io_deviceTree_b_ready ),
       .io_deviceTree_b_valid( deviceTree_io_b_valid ),
       //.io_deviceTree_b_bits_resp(  )
       //.io_deviceTree_b_bits_id(  )
       //.io_deviceTree_b_bits_user(  )
       .io_deviceTree_ar_ready( deviceTree_io_ar_ready ),
       .io_deviceTree_ar_valid( outmemsys_io_deviceTree_ar_valid ),
       .io_deviceTree_ar_bits_addr( outmemsys_io_deviceTree_ar_bits_addr ),
       .io_deviceTree_ar_bits_len( outmemsys_io_deviceTree_ar_bits_len ),
       .io_deviceTree_ar_bits_size( outmemsys_io_deviceTree_ar_bits_size ),
       .io_deviceTree_ar_bits_burst( outmemsys_io_deviceTree_ar_bits_burst ),
       .io_deviceTree_ar_bits_lock( outmemsys_io_deviceTree_ar_bits_lock ),
       .io_deviceTree_ar_bits_cache( outmemsys_io_deviceTree_ar_bits_cache ),
       .io_deviceTree_ar_bits_prot( outmemsys_io_deviceTree_ar_bits_prot ),
       .io_deviceTree_ar_bits_qos( outmemsys_io_deviceTree_ar_bits_qos ),
       .io_deviceTree_ar_bits_region( outmemsys_io_deviceTree_ar_bits_region ),
       .io_deviceTree_ar_bits_id( outmemsys_io_deviceTree_ar_bits_id ),
       .io_deviceTree_ar_bits_user( outmemsys_io_deviceTree_ar_bits_user ),
       .io_deviceTree_r_ready( outmemsys_io_deviceTree_r_ready ),
       .io_deviceTree_r_valid( deviceTree_io_r_valid ),
       .io_deviceTree_r_bits_resp( deviceTree_io_r_bits_resp ),
       .io_deviceTree_r_bits_data( deviceTree_io_r_bits_data ),
       .io_deviceTree_r_bits_last( deviceTree_io_r_bits_last ),
       .io_deviceTree_r_bits_id( deviceTree_io_r_bits_id ),
       .io_deviceTree_r_bits_user( deviceTree_io_r_bits_user )
       //.io_dma_req_ready(  )
       //.io_dma_req_valid(  )
       //.io_dma_req_bits_client_xact_id(  )
       //.io_dma_req_bits_cmd(  )
       //.io_dma_req_bits_source(  )
       //.io_dma_req_bits_dest(  )
       //.io_dma_req_bits_length(  )
       //.io_dma_resp_ready(  )
       //.io_dma_resp_valid(  )
       //.io_dma_resp_bits_client_xact_id(  )
       //.io_dma_resp_bits_status(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign outmemsys.io_deviceTree_b_bits_resp = {1{$random}};
    assign outmemsys.io_deviceTree_b_bits_id = {1{$random}};
    assign outmemsys.io_deviceTree_b_bits_user = {1{$random}};
// synthesis translate_on
`endif
  SMIArbiter_0 SMIArbiter(.clk(clk), .reset(reset),
       .io_in_1_req_ready( SMIArbiter_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_csr_0_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_csr_0_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_csr_0_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_csr_0_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_csr_0_resp_ready ),
       .io_in_1_resp_valid( SMIArbiter_io_in_1_resp_valid ),
       .io_in_1_resp_bits( SMIArbiter_io_in_1_resp_bits ),
       .io_in_0_req_ready( SMIArbiter_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_cpu_0_csr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_cpu_0_csr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_cpu_0_csr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_cpu_0_csr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_cpu_0_csr_resp_ready ),
       .io_in_0_resp_valid( SMIArbiter_io_in_0_resp_valid ),
       .io_in_0_resp_bits( SMIArbiter_io_in_0_resp_bits ),
       .io_out_req_ready( io_htif_0_csr_req_ready ),
       .io_out_req_valid( SMIArbiter_io_out_req_valid ),
       .io_out_req_bits_rw( SMIArbiter_io_out_req_bits_rw ),
       .io_out_req_bits_addr( SMIArbiter_io_out_req_bits_addr ),
       .io_out_req_bits_data( SMIArbiter_io_out_req_bits_data ),
       .io_out_resp_ready( SMIArbiter_io_out_resp_ready ),
       .io_out_resp_valid( io_htif_0_csr_resp_valid ),
       .io_out_resp_bits( io_htif_0_csr_resp_bits )
  );
  SCRFile scrFile(.clk(clk), .reset(reset),
       .io_smi_req_ready( scrFile_io_smi_req_ready ),
       .io_smi_req_valid( scrArb_io_out_req_valid ),
       .io_smi_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_smi_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_smi_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_smi_resp_ready( scrArb_io_out_resp_ready ),
       .io_smi_resp_valid( scrFile_io_smi_resp_valid ),
       .io_smi_resp_bits( scrFile_io_smi_resp_bits )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign scrFile.io_scr_rdata_63 = {2{$random}};
    assign scrFile.io_scr_rdata_62 = {2{$random}};
    assign scrFile.io_scr_rdata_61 = {2{$random}};
    assign scrFile.io_scr_rdata_60 = {2{$random}};
    assign scrFile.io_scr_rdata_59 = {2{$random}};
    assign scrFile.io_scr_rdata_58 = {2{$random}};
    assign scrFile.io_scr_rdata_57 = {2{$random}};
    assign scrFile.io_scr_rdata_56 = {2{$random}};
    assign scrFile.io_scr_rdata_55 = {2{$random}};
    assign scrFile.io_scr_rdata_54 = {2{$random}};
    assign scrFile.io_scr_rdata_53 = {2{$random}};
    assign scrFile.io_scr_rdata_52 = {2{$random}};
    assign scrFile.io_scr_rdata_51 = {2{$random}};
    assign scrFile.io_scr_rdata_50 = {2{$random}};
    assign scrFile.io_scr_rdata_49 = {2{$random}};
    assign scrFile.io_scr_rdata_48 = {2{$random}};
    assign scrFile.io_scr_rdata_47 = {2{$random}};
    assign scrFile.io_scr_rdata_46 = {2{$random}};
    assign scrFile.io_scr_rdata_45 = {2{$random}};
    assign scrFile.io_scr_rdata_44 = {2{$random}};
    assign scrFile.io_scr_rdata_43 = {2{$random}};
    assign scrFile.io_scr_rdata_42 = {2{$random}};
    assign scrFile.io_scr_rdata_41 = {2{$random}};
    assign scrFile.io_scr_rdata_40 = {2{$random}};
    assign scrFile.io_scr_rdata_39 = {2{$random}};
    assign scrFile.io_scr_rdata_38 = {2{$random}};
    assign scrFile.io_scr_rdata_37 = {2{$random}};
    assign scrFile.io_scr_rdata_36 = {2{$random}};
    assign scrFile.io_scr_rdata_35 = {2{$random}};
    assign scrFile.io_scr_rdata_34 = {2{$random}};
    assign scrFile.io_scr_rdata_33 = {2{$random}};
    assign scrFile.io_scr_rdata_32 = {2{$random}};
    assign scrFile.io_scr_rdata_31 = {2{$random}};
    assign scrFile.io_scr_rdata_30 = {2{$random}};
    assign scrFile.io_scr_rdata_29 = {2{$random}};
    assign scrFile.io_scr_rdata_28 = {2{$random}};
    assign scrFile.io_scr_rdata_27 = {2{$random}};
    assign scrFile.io_scr_rdata_26 = {2{$random}};
    assign scrFile.io_scr_rdata_25 = {2{$random}};
    assign scrFile.io_scr_rdata_24 = {2{$random}};
    assign scrFile.io_scr_rdata_23 = {2{$random}};
    assign scrFile.io_scr_rdata_22 = {2{$random}};
    assign scrFile.io_scr_rdata_21 = {2{$random}};
    assign scrFile.io_scr_rdata_20 = {2{$random}};
    assign scrFile.io_scr_rdata_19 = {2{$random}};
    assign scrFile.io_scr_rdata_18 = {2{$random}};
    assign scrFile.io_scr_rdata_17 = {2{$random}};
    assign scrFile.io_scr_rdata_16 = {2{$random}};
    assign scrFile.io_scr_rdata_15 = {2{$random}};
    assign scrFile.io_scr_rdata_14 = {2{$random}};
    assign scrFile.io_scr_rdata_13 = {2{$random}};
    assign scrFile.io_scr_rdata_12 = {2{$random}};
    assign scrFile.io_scr_rdata_11 = {2{$random}};
    assign scrFile.io_scr_rdata_10 = {2{$random}};
    assign scrFile.io_scr_rdata_9 = {2{$random}};
    assign scrFile.io_scr_rdata_8 = {2{$random}};
    assign scrFile.io_scr_rdata_7 = {2{$random}};
    assign scrFile.io_scr_rdata_6 = {2{$random}};
    assign scrFile.io_scr_rdata_5 = {2{$random}};
    assign scrFile.io_scr_rdata_4 = {2{$random}};
    assign scrFile.io_scr_rdata_3 = {2{$random}};
    assign scrFile.io_scr_rdata_2 = {2{$random}};
// synthesis translate_on
`endif
  SMIArbiter_1 scrArb(.clk(clk), .reset(reset),
       .io_in_1_req_ready( scrArb_io_in_1_req_ready ),
       .io_in_1_req_valid( outmemsys_io_scr_req_valid ),
       .io_in_1_req_bits_rw( outmemsys_io_scr_req_bits_rw ),
       .io_in_1_req_bits_addr( outmemsys_io_scr_req_bits_addr ),
       .io_in_1_req_bits_data( outmemsys_io_scr_req_bits_data ),
       .io_in_1_resp_ready( outmemsys_io_scr_resp_ready ),
       .io_in_1_resp_valid( scrArb_io_in_1_resp_valid ),
       .io_in_1_resp_bits( scrArb_io_in_1_resp_bits ),
       .io_in_0_req_ready( scrArb_io_in_0_req_ready ),
       .io_in_0_req_valid( htif_io_scr_req_valid ),
       .io_in_0_req_bits_rw( htif_io_scr_req_bits_rw ),
       .io_in_0_req_bits_addr( htif_io_scr_req_bits_addr ),
       .io_in_0_req_bits_data( htif_io_scr_req_bits_data ),
       .io_in_0_resp_ready( htif_io_scr_resp_ready ),
       .io_in_0_resp_valid( scrArb_io_in_0_resp_valid ),
       .io_in_0_resp_bits( scrArb_io_in_0_resp_bits ),
       .io_out_req_ready( scrFile_io_smi_req_ready ),
       .io_out_req_valid( scrArb_io_out_req_valid ),
       .io_out_req_bits_rw( scrArb_io_out_req_bits_rw ),
       .io_out_req_bits_addr( scrArb_io_out_req_bits_addr ),
       .io_out_req_bits_data( scrArb_io_out_req_bits_data ),
       .io_out_resp_ready( scrArb_io_out_resp_ready ),
       .io_out_resp_valid( scrFile_io_smi_resp_valid ),
       .io_out_resp_bits( scrFile_io_smi_resp_bits )
  );
  NastiROM deviceTree(.clk(clk), .reset(reset),
       .io_aw_ready( deviceTree_io_aw_ready ),
       .io_aw_valid( outmemsys_io_deviceTree_aw_valid ),
       .io_aw_bits_addr( outmemsys_io_deviceTree_aw_bits_addr ),
       .io_aw_bits_len( outmemsys_io_deviceTree_aw_bits_len ),
       .io_aw_bits_size( outmemsys_io_deviceTree_aw_bits_size ),
       .io_aw_bits_burst( outmemsys_io_deviceTree_aw_bits_burst ),
       .io_aw_bits_lock( outmemsys_io_deviceTree_aw_bits_lock ),
       .io_aw_bits_cache( outmemsys_io_deviceTree_aw_bits_cache ),
       .io_aw_bits_prot( outmemsys_io_deviceTree_aw_bits_prot ),
       .io_aw_bits_qos( outmemsys_io_deviceTree_aw_bits_qos ),
       .io_aw_bits_region( outmemsys_io_deviceTree_aw_bits_region ),
       .io_aw_bits_id( outmemsys_io_deviceTree_aw_bits_id ),
       .io_aw_bits_user( outmemsys_io_deviceTree_aw_bits_user ),
       .io_w_ready( deviceTree_io_w_ready ),
       .io_w_valid( outmemsys_io_deviceTree_w_valid ),
       .io_w_bits_data( outmemsys_io_deviceTree_w_bits_data ),
       .io_w_bits_last( outmemsys_io_deviceTree_w_bits_last ),
       .io_w_bits_strb( outmemsys_io_deviceTree_w_bits_strb ),
       .io_w_bits_user( outmemsys_io_deviceTree_w_bits_user ),
       .io_b_ready( outmemsys_io_deviceTree_b_ready ),
       .io_b_valid( deviceTree_io_b_valid ),
       //.io_b_bits_resp(  )
       //.io_b_bits_id(  )
       //.io_b_bits_user(  )
       .io_ar_ready( deviceTree_io_ar_ready ),
       .io_ar_valid( outmemsys_io_deviceTree_ar_valid ),
       .io_ar_bits_addr( outmemsys_io_deviceTree_ar_bits_addr ),
       .io_ar_bits_len( outmemsys_io_deviceTree_ar_bits_len ),
       .io_ar_bits_size( outmemsys_io_deviceTree_ar_bits_size ),
       .io_ar_bits_burst( outmemsys_io_deviceTree_ar_bits_burst ),
       .io_ar_bits_lock( outmemsys_io_deviceTree_ar_bits_lock ),
       .io_ar_bits_cache( outmemsys_io_deviceTree_ar_bits_cache ),
       .io_ar_bits_prot( outmemsys_io_deviceTree_ar_bits_prot ),
       .io_ar_bits_qos( outmemsys_io_deviceTree_ar_bits_qos ),
       .io_ar_bits_region( outmemsys_io_deviceTree_ar_bits_region ),
       .io_ar_bits_id( outmemsys_io_deviceTree_ar_bits_id ),
       .io_ar_bits_user( outmemsys_io_deviceTree_ar_bits_user ),
       .io_r_ready( outmemsys_io_deviceTree_r_ready ),
       .io_r_valid( deviceTree_io_r_valid ),
       .io_r_bits_resp( deviceTree_io_r_bits_resp ),
       .io_r_bits_data( deviceTree_io_r_bits_data ),
       .io_r_bits_last( deviceTree_io_r_bits_last ),
       .io_r_bits_id( deviceTree_io_r_bits_id ),
       .io_r_bits_user( deviceTree_io_r_bits_user )
  );
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    input [11:0] io_rw_addr,
    input [2:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output io_csr_stall,
    output io_csr_xcpt,
    output io_eret,
    output io_status_sd,
    output[30:0] io_status_zero2,
    output io_status_sd_rv32,
    output[8:0] io_status_zero1,
    output[4:0] io_status_vm,
    output io_status_mprv,
    output[1:0] io_status_xs,
    output[1:0] io_status_fs,
    output[1:0] io_status_prv3,
    output io_status_ie3,
    output[1:0] io_status_prv2,
    output io_status_ie2,
    output[1:0] io_status_prv1,
    output io_status_ie1,
    output[1:0] io_status_prv,
    output io_status_ie,
    output[31:0] io_ptbr,
    output[39:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input [39:0] io_pc,
    output io_fatc,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_autl_acquire_ready
    input  io_rocc_autl_acquire_valid,
    input [25:0] io_rocc_autl_acquire_bits_addr_block,
    input [1:0] io_rocc_autl_acquire_bits_client_xact_id,
    input [1:0] io_rocc_autl_acquire_bits_addr_beat,
    input  io_rocc_autl_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_autl_acquire_bits_a_type,
    input [16:0] io_rocc_autl_acquire_bits_union,
    input [127:0] io_rocc_autl_acquire_bits_data,
    input  io_rocc_autl_grant_ready,
    //output io_rocc_autl_grant_valid
    //output[1:0] io_rocc_autl_grant_bits_addr_beat
    //output[1:0] io_rocc_autl_grant_bits_client_xact_id
    //output[2:0] io_rocc_autl_grant_bits_manager_xact_id
    //output io_rocc_autl_grant_bits_is_builtin_type
    //output[3:0] io_rocc_autl_grant_bits_g_type
    //output[127:0] io_rocc_autl_grant_bits_data
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    //output io_rocc_fpu_req_ready
    input  io_rocc_fpu_req_valid,
    input [4:0] io_rocc_fpu_req_bits_cmd,
    input  io_rocc_fpu_req_bits_ldst,
    input  io_rocc_fpu_req_bits_wen,
    input  io_rocc_fpu_req_bits_ren1,
    input  io_rocc_fpu_req_bits_ren2,
    input  io_rocc_fpu_req_bits_ren3,
    input  io_rocc_fpu_req_bits_swap12,
    input  io_rocc_fpu_req_bits_swap23,
    input  io_rocc_fpu_req_bits_single,
    input  io_rocc_fpu_req_bits_fromint,
    input  io_rocc_fpu_req_bits_toint,
    input  io_rocc_fpu_req_bits_fastpipe,
    input  io_rocc_fpu_req_bits_fma,
    input  io_rocc_fpu_req_bits_div,
    input  io_rocc_fpu_req_bits_sqrt,
    input  io_rocc_fpu_req_bits_round,
    input  io_rocc_fpu_req_bits_wflags,
    input [2:0] io_rocc_fpu_req_bits_rm,
    input [1:0] io_rocc_fpu_req_bits_typ,
    input [64:0] io_rocc_fpu_req_bits_in1,
    input [64:0] io_rocc_fpu_req_bits_in2,
    input [64:0] io_rocc_fpu_req_bits_in3,
    input  io_rocc_fpu_resp_ready,
    //output io_rocc_fpu_resp_valid
    //output[64:0] io_rocc_fpu_resp_bits_data
    //output[4:0] io_rocc_fpu_resp_bits_exc
    //output io_rocc_exception
    //output io_rocc_dma_req_ready
    input  io_rocc_dma_req_valid,
    input [1:0] io_rocc_dma_req_bits_client_xact_id,
    input [1:0] io_rocc_dma_req_bits_cmd,
    input [31:0] io_rocc_dma_req_bits_source,
    input [31:0] io_rocc_dma_req_bits_dest,
    input [31:0] io_rocc_dma_req_bits_length,
    input  io_rocc_dma_resp_ready,
    //output io_rocc_dma_resp_valid
    //output[1:0] io_rocc_dma_resp_bits_client_xact_id
    //output[1:0] io_rocc_dma_resp_bits_status
    output io_interrupt,
    output[63:0] io_interrupt_cause
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire csr_xcpt;
  wire insn_break;
  wire system_insn;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire insn_call;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire priv_sufficient;
  reg [1:0] reg_mstatus_prv;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  reg [1:0] reg_mstatus_prv1;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire[1:0] T30;
  reg [1:0] reg_mstatus_prv2;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T35;
  wire[63:0] wdata;
  wire[63:0] T36;
  wire[63:0] T37;
  reg [63:0] host_csr_bits_data;
  wire[63:0] T38;
  wire[63:0] T39;
  wire T40;
  wire host_csr_req_fire;
  wire T41;
  wire cpu_ren;
  wire T42;
  wire T43;
  reg  host_csr_req_valid;
  wire T44;
  wire T45;
  wire[63:0] T46;
  wire T47;
  wire[63:0] T48;
  wire[63:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire[11:0] addr;
  reg [11:0] host_csr_bits_addr;
  wire[11:0] T60;
  wire wen;
  wire T61;
  reg  host_csr_bits_rw;
  wire T62;
  wire T63;
  wire T64;
  wire read_only;
  wire[1:0] T65;
  wire cpu_wen;
  wire T66;
  wire T67;
  wire[1:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire[1:0] T881;
  wire T75;
  wire T76;
  wire T77;
  wire insn_ret;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire insn_redirect_trap;
  wire maybe_insn_redirect_trap;
  wire T86;
  wire[1:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire[1:0] csr_addr_priv;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire fp_csr;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire addr_valid;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire[1:0] T882;
  wire[2:0] T883;
  wire[1:0] T215;
  wire[1:0] T216;
  wire[1:0] T884;
  wire[63:0] T217;
  wire[63:0] T218;
  wire[63:0] T219;
  wire[63:0] T220;
  wire[63:0] T221;
  wire T222;
  wire T223;
  wire T224;
  reg  reg_mstatus_ie;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  reg  reg_mstatus_ie1;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  reg  reg_mstatus_ie2;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  reg  reg_mip_ssip;
  wire T885;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  reg  reg_mie_ssip;
  wire T886;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  reg  reg_mip_msip;
  wire T887;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  reg  reg_mie_msip;
  wire T888;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  reg  reg_mip_stip;
  wire T889;
  wire T277;
  wire T278;
  reg  reg_mie_stip;
  wire T890;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  reg  reg_mip_mtip;
  wire T891;
  wire T289;
  wire T290;
  wire T291;
  reg [63:0] read_time;
  wire[63:0] T292;
  wire T293;
  reg [63:0] reg_mtimecmp;
  wire[63:0] T294;
  wire T295;
  reg  reg_mie_mtip;
  wire T892;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  reg [63:0] reg_fromhost;
  wire[63:0] T893;
  wire[63:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  reg [2:0] reg_frm;
  wire[2:0] T894;
  wire[63:0] T311;
  wire[63:0] T312;
  wire[63:0] T895;
  wire T313;
  wire[63:0] T896;
  wire[58:0] T314;
  wire T315;
  wire[63:0] T316;
  reg [5:0] R317;
  wire[5:0] T897;
  wire[5:0] T318;
  wire[6:0] T319;
  wire[6:0] T898;
  reg [57:0] R320;
  wire[57:0] T899;
  wire[57:0] T321;
  wire[57:0] T322;
  wire T323;
  wire insn_sfence_vm;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire[39:0] T331;
  wire[39:0] T332;
  wire[39:0] T333;
  reg [39:0] reg_sepc;
  wire[39:0] T900;
  wire[63:0] T334;
  wire[63:0] T901;
  wire[39:0] T335;
  wire[63:0] T336;
  wire[63:0] T337;
  wire[63:0] T338;
  wire T339;
  reg [39:0] reg_mepc;
  wire[39:0] T902;
  wire[63:0] T340;
  wire[63:0] T903;
  wire[39:0] T341;
  wire[39:0] T342;
  wire[39:0] T343;
  wire[39:0] T344;
  wire[63:0] T345;
  wire[63:0] T346;
  wire[63:0] T347;
  wire T348;
  wire T349;
  wire[39:0] T350;
  reg [38:0] reg_stvec;
  wire[38:0] T904;
  wire[63:0] T351;
  wire[63:0] T905;
  wire[63:0] T352;
  wire[63:0] T353;
  wire[63:0] T354;
  wire T355;
  wire T356;
  wire[39:0] T906;
  wire[8:0] T357;
  wire[8:0] T907;
  wire[7:0] T358;
  wire T359;
  reg [31:0] reg_sptbr;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[19:0] T362;
  wire T363;
  reg  reg_mstatus_ie3;
  wire T364;
  reg [1:0] reg_mstatus_prv3;
  wire[1:0] T365;
  wire[1:0] T366;
  wire[1:0] T908;
  wire T367;
  reg [1:0] reg_mstatus_fs;
  wire[1:0] T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[1:0] T909;
  wire T374;
  reg [1:0] reg_mstatus_xs;
  wire[1:0] T375;
  reg  reg_mstatus_mprv;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  reg [4:0] reg_mstatus_vm;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire T385;
  wire T386;
  wire[4:0] T387;
  wire T388;
  wire T389;
  reg [8:0] reg_mstatus_zero1;
  wire[8:0] T390;
  reg  reg_mstatus_sd_rv32;
  wire T391;
  reg [30:0] reg_mstatus_zero2;
  wire[30:0] T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg  reg_wfi;
  wire T910;
  wire T397;
  wire T398;
  wire insn_wfi;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire some_interrupt_pending;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[63:0] T420;
  wire[63:0] T421;
  wire[63:0] T422;
  wire[24:0] T423;
  wire[24:0] T911;
  wire T424;
  wire[63:0] T425;
  wire[63:0] T426;
  wire[63:0] T427;
  wire[23:0] T428;
  wire[23:0] T912;
  wire T429;
  wire[63:0] T430;
  wire[63:0] T431;
  wire[63:0] T913;
  wire[31:0] T432;
  wire[63:0] T433;
  wire[63:0] T434;
  wire[63:0] T435;
  reg [39:0] reg_sbadaddr;
  wire[39:0] T436;
  reg [39:0] reg_mbadaddr;
  wire[39:0] T437;
  wire[39:0] T438;
  wire[39:0] T439;
  wire[39:0] T440;
  wire[38:0] T441;
  wire T442;
  wire T443;
  wire[24:0] T444;
  wire T445;
  wire T446;
  wire[38:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire[39:0] T456;
  wire T457;
  wire[23:0] T458;
  wire[23:0] T914;
  wire T459;
  wire[63:0] T460;
  wire[63:0] T461;
  reg [63:0] reg_scause;
  wire[63:0] T462;
  reg [63:0] reg_mcause;
  wire[63:0] T463;
  wire[63:0] T464;
  wire[63:0] T465;
  wire[63:0] T466;
  wire[63:0] T467;
  wire T468;
  wire T469;
  wire[63:0] T915;
  wire[3:0] T470;
  wire[3:0] T916;
  wire T471;
  wire[63:0] T472;
  wire T473;
  wire[63:0] T474;
  wire[63:0] T475;
  reg [63:0] reg_sscratch;
  wire[63:0] T476;
  wire T477;
  wire[63:0] T478;
  wire[63:0] T917;
  wire[7:0] T479;
  wire[7:0] T480;
  wire[7:0] T481;
  wire[3:0] T482;
  wire[1:0] T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[1:0] T490;
  wire T491;
  wire T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire[63:0] T496;
  wire[63:0] T918;
  wire[7:0] T497;
  wire[7:0] T498;
  wire[7:0] T499;
  wire[3:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire T505;
  wire T506;
  wire[3:0] T507;
  wire[1:0] T508;
  wire T509;
  wire T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire[63:0] T514;
  wire[63:0] T515;
  wire[63:0] T516;
  wire[63:0] T517;
  wire[13:0] T518;
  wire[3:0] T519;
  wire[2:0] T520;
  wire T521;
  wire T522;
  wire[63:0] read_mstatus;
  wire[63:0] T523;
  wire[11:0] T524;
  wire[5:0] T525;
  wire[2:0] T526;
  wire[2:0] T527;
  wire[5:0] T528;
  wire[2:0] T529;
  wire[2:0] T530;
  wire[51:0] T531;
  wire[9:0] T532;
  wire[3:0] T533;
  wire[5:0] T534;
  wire[41:0] T535;
  wire[9:0] T536;
  wire[31:0] T537;
  wire[1:0] T538;
  wire T539;
  wire T540;
  wire[9:0] T541;
  wire[7:0] T542;
  wire T543;
  wire T544;
  wire[6:0] T545;
  wire[1:0] T546;
  wire[1:0] T547;
  wire[49:0] T548;
  wire[16:0] T549;
  wire[2:0] T550;
  wire[1:0] T551;
  wire[1:0] T552;
  wire T553;
  wire T554;
  wire[13:0] T555;
  wire[32:0] T556;
  wire[31:0] T557;
  wire T558;
  wire T559;
  wire[30:0] T560;
  wire T561;
  wire T562;
  wire[63:0] T563;
  wire[63:0] T564;
  wire[63:0] T565;
  reg [5:0] R566;
  wire[5:0] T919;
  wire[5:0] T567;
  wire[5:0] T568;
  wire[6:0] T569;
  wire[6:0] T920;
  wire T570;
  reg [57:0] R571;
  wire[57:0] T921;
  wire[57:0] T572;
  wire[57:0] T573;
  wire T574;
  wire T575;
  wire[63:0] T576;
  wire[63:0] T577;
  wire[63:0] T578;
  reg [5:0] R579;
  wire[5:0] T922;
  wire[5:0] T580;
  wire[5:0] T581;
  wire[6:0] T582;
  wire[6:0] T923;
  wire T583;
  reg [57:0] R584;
  wire[57:0] T924;
  wire[57:0] T585;
  wire[57:0] T586;
  wire T587;
  wire T588;
  wire[63:0] T589;
  wire[63:0] T590;
  wire[63:0] T591;
  reg [5:0] R592;
  wire[5:0] T925;
  wire[5:0] T593;
  wire[5:0] T594;
  wire[6:0] T595;
  wire[6:0] T926;
  wire T596;
  reg [57:0] R597;
  wire[57:0] T927;
  wire[57:0] T598;
  wire[57:0] T599;
  wire T600;
  wire T601;
  wire[63:0] T602;
  wire[63:0] T603;
  wire[63:0] T604;
  reg [5:0] R605;
  wire[5:0] T928;
  wire[5:0] T606;
  wire[5:0] T607;
  wire[6:0] T608;
  wire[6:0] T929;
  wire T609;
  reg [57:0] R610;
  wire[57:0] T930;
  wire[57:0] T611;
  wire[57:0] T612;
  wire T613;
  wire T614;
  wire[63:0] T615;
  wire[63:0] T616;
  wire[63:0] T617;
  reg [5:0] R618;
  wire[5:0] T931;
  wire[5:0] T619;
  wire[5:0] T620;
  wire[6:0] T621;
  wire[6:0] T932;
  wire T622;
  reg [57:0] R623;
  wire[57:0] T933;
  wire[57:0] T624;
  wire[57:0] T625;
  wire T626;
  wire T627;
  wire[63:0] T628;
  wire[63:0] T629;
  wire[63:0] T630;
  reg [5:0] R631;
  wire[5:0] T934;
  wire[5:0] T632;
  wire[5:0] T633;
  wire[6:0] T634;
  wire[6:0] T935;
  wire T635;
  reg [57:0] R636;
  wire[57:0] T936;
  wire[57:0] T637;
  wire[57:0] T638;
  wire T639;
  wire T640;
  wire[63:0] T641;
  wire[63:0] T642;
  wire[63:0] T643;
  reg [5:0] R644;
  wire[5:0] T937;
  wire[5:0] T645;
  wire[5:0] T646;
  wire[6:0] T647;
  wire[6:0] T938;
  wire T648;
  reg [57:0] R649;
  wire[57:0] T939;
  wire[57:0] T650;
  wire[57:0] T651;
  wire T652;
  wire T653;
  wire[63:0] T654;
  wire[63:0] T655;
  wire[63:0] T656;
  reg [5:0] R657;
  wire[5:0] T940;
  wire[5:0] T658;
  wire[5:0] T659;
  wire[6:0] T660;
  wire[6:0] T941;
  wire T661;
  reg [57:0] R662;
  wire[57:0] T942;
  wire[57:0] T663;
  wire[57:0] T664;
  wire T665;
  wire T666;
  wire[63:0] T667;
  wire[63:0] T668;
  wire[63:0] T669;
  reg [5:0] R670;
  wire[5:0] T943;
  wire[5:0] T671;
  wire[5:0] T672;
  wire[6:0] T673;
  wire[6:0] T944;
  wire T674;
  reg [57:0] R675;
  wire[57:0] T945;
  wire[57:0] T676;
  wire[57:0] T677;
  wire T678;
  wire T679;
  wire[63:0] T680;
  wire[63:0] T681;
  wire[63:0] T682;
  reg [5:0] R683;
  wire[5:0] T946;
  wire[5:0] T684;
  wire[5:0] T685;
  wire[6:0] T686;
  wire[6:0] T947;
  wire T687;
  reg [57:0] R688;
  wire[57:0] T948;
  wire[57:0] T689;
  wire[57:0] T690;
  wire T691;
  wire T692;
  wire[63:0] T693;
  wire[63:0] T694;
  wire[63:0] T695;
  reg [5:0] R696;
  wire[5:0] T949;
  wire[5:0] T697;
  wire[5:0] T698;
  wire[6:0] T699;
  wire[6:0] T950;
  wire T700;
  reg [57:0] R701;
  wire[57:0] T951;
  wire[57:0] T702;
  wire[57:0] T703;
  wire T704;
  wire T705;
  wire[63:0] T706;
  wire[63:0] T707;
  wire[63:0] T708;
  reg [5:0] R709;
  wire[5:0] T952;
  wire[5:0] T710;
  wire[5:0] T711;
  wire[6:0] T712;
  wire[6:0] T953;
  wire T713;
  reg [57:0] R714;
  wire[57:0] T954;
  wire[57:0] T715;
  wire[57:0] T716;
  wire T717;
  wire T718;
  wire[63:0] T719;
  wire[63:0] T720;
  wire[63:0] T721;
  reg [5:0] R722;
  wire[5:0] T955;
  wire[5:0] T723;
  wire[5:0] T724;
  wire[6:0] T725;
  wire[6:0] T956;
  wire T726;
  reg [57:0] R727;
  wire[57:0] T957;
  wire[57:0] T728;
  wire[57:0] T729;
  wire T730;
  wire T731;
  wire[63:0] T732;
  wire[63:0] T733;
  wire[63:0] T734;
  reg [5:0] R735;
  wire[5:0] T958;
  wire[5:0] T736;
  wire[5:0] T737;
  wire[6:0] T738;
  wire[6:0] T959;
  wire T739;
  reg [57:0] R740;
  wire[57:0] T960;
  wire[57:0] T741;
  wire[57:0] T742;
  wire T743;
  wire T744;
  wire[63:0] T745;
  wire[63:0] T746;
  wire[63:0] T747;
  reg [5:0] R748;
  wire[5:0] T961;
  wire[5:0] T749;
  wire[5:0] T750;
  wire[6:0] T751;
  wire[6:0] T962;
  wire T752;
  reg [57:0] R753;
  wire[57:0] T963;
  wire[57:0] T754;
  wire[57:0] T755;
  wire T756;
  wire T757;
  wire[63:0] T758;
  wire[63:0] T759;
  wire[63:0] T760;
  reg [5:0] R761;
  wire[5:0] T964;
  wire[5:0] T762;
  wire[5:0] T763;
  wire[6:0] T764;
  wire[6:0] T965;
  wire T765;
  reg [57:0] R766;
  wire[57:0] T966;
  wire[57:0] T767;
  wire[57:0] T768;
  wire T769;
  wire T770;
  wire[63:0] T771;
  wire[63:0] T772;
  wire[63:0] T773;
  reg [5:0] R774;
  wire[5:0] T967;
  wire[5:0] T775;
  wire[5:0] T776;
  wire[5:0] T777;
  wire[6:0] T778;
  wire[6:0] T968;
  wire T779;
  wire[5:0] T780;
  wire T781;
  reg [57:0] R782;
  wire[57:0] T969;
  wire[57:0] T783;
  wire[57:0] T784;
  wire[57:0] T785;
  wire T786;
  wire T787;
  wire[57:0] T788;
  wire[63:0] T789;
  wire[63:0] T790;
  wire[63:0] T791;
  wire[63:0] T792;
  wire[63:0] T793;
  wire[63:0] T794;
  reg [63:0] reg_tohost;
  wire[63:0] T970;
  wire[63:0] T795;
  wire[63:0] T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[63:0] T804;
  wire[63:0] T971;
  wire T805;
  reg  reg_stats;
  wire T972;
  wire T806;
  wire T807;
  wire T808;
  wire[63:0] T809;
  wire[63:0] T973;
  wire T810;
  wire[63:0] T811;
  wire[63:0] T812;
  wire[63:0] T813;
  wire[63:0] T814;
  wire[63:0] T815;
  wire[63:0] T816;
  wire[63:0] T817;
  wire[23:0] T818;
  wire[23:0] T974;
  wire T819;
  wire[63:0] T820;
  wire[63:0] T821;
  wire[63:0] T822;
  wire[23:0] T823;
  wire[23:0] T975;
  wire T824;
  wire[63:0] T825;
  wire[63:0] T826;
  reg [63:0] reg_mscratch;
  wire[63:0] T827;
  wire T828;
  wire[63:0] T829;
  wire[63:0] T976;
  wire[7:0] T830;
  wire[7:0] T831;
  wire[7:0] T832;
  wire[3:0] T833;
  wire[1:0] T834;
  reg  reg_mie_usip;
  wire T977;
  wire[1:0] T835;
  reg  reg_mie_hsip;
  wire T978;
  wire[3:0] T836;
  wire[1:0] T837;
  reg  reg_mie_utip;
  wire T979;
  wire[1:0] T838;
  reg  reg_mie_htip;
  wire T980;
  wire[63:0] T839;
  wire[63:0] T981;
  wire[7:0] T840;
  wire[7:0] T841;
  wire[7:0] T842;
  wire[3:0] T843;
  wire[1:0] T844;
  reg  reg_mip_usip;
  wire T982;
  wire[1:0] T845;
  reg  reg_mip_hsip;
  wire T983;
  wire[3:0] T846;
  wire[1:0] T847;
  reg  reg_mip_utip;
  wire T984;
  wire[1:0] T848;
  reg  reg_mip_htip;
  wire T985;
  wire[63:0] T849;
  wire[63:0] T850;
  wire[63:0] T986;
  wire[30:0] T851;
  wire[63:0] T852;
  wire[63:0] T987;
  wire[8:0] T853;
  wire[63:0] T854;
  wire[63:0] T855;
  wire[63:0] T856;
  wire[63:0] T857;
  wire[63:0] T858;
  wire[63:0] T988;
  wire[63:0] T859;
  wire[63:0] T860;
  wire[63:0] T861;
  wire[63:0] T862;
  wire[63:0] T863;
  wire[63:0] T864;
  wire[63:0] T865;
  wire[63:0] T866;
  wire[63:0] T867;
  wire[63:0] T868;
  wire[63:0] T869;
  wire[63:0] T870;
  wire[63:0] T871;
  wire[63:0] T872;
  wire[63:0] T873;
  wire[63:0] T874;
  reg  host_csr_rep_valid;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    reg_mstatus_prv = {1{$random}};
    reg_mstatus_prv1 = {1{$random}};
    reg_mstatus_prv2 = {1{$random}};
    host_csr_bits_data = {2{$random}};
    host_csr_req_valid = {1{$random}};
    host_csr_bits_addr = {1{$random}};
    host_csr_bits_rw = {1{$random}};
    reg_mstatus_ie = {1{$random}};
    reg_mstatus_ie1 = {1{$random}};
    reg_mstatus_ie2 = {1{$random}};
    reg_mip_ssip = {1{$random}};
    reg_mie_ssip = {1{$random}};
    reg_mip_msip = {1{$random}};
    reg_mie_msip = {1{$random}};
    reg_mip_stip = {1{$random}};
    reg_mie_stip = {1{$random}};
    reg_mip_mtip = {1{$random}};
    read_time = {2{$random}};
    reg_mtimecmp = {2{$random}};
    reg_mie_mtip = {1{$random}};
    reg_fromhost = {2{$random}};
    reg_frm = {1{$random}};
    R317 = {1{$random}};
    R320 = {2{$random}};
    reg_sepc = {2{$random}};
    reg_mepc = {2{$random}};
    reg_stvec = {2{$random}};
    reg_sptbr = {1{$random}};
    reg_mstatus_ie3 = {1{$random}};
    reg_mstatus_prv3 = {1{$random}};
    reg_mstatus_fs = {1{$random}};
    reg_mstatus_xs = {1{$random}};
    reg_mstatus_mprv = {1{$random}};
    reg_mstatus_vm = {1{$random}};
    reg_mstatus_zero1 = {1{$random}};
    reg_mstatus_sd_rv32 = {1{$random}};
    reg_mstatus_zero2 = {1{$random}};
    reg_wfi = {1{$random}};
    reg_sbadaddr = {2{$random}};
    reg_mbadaddr = {2{$random}};
    reg_scause = {2{$random}};
    reg_mcause = {2{$random}};
    reg_sscratch = {2{$random}};
    R566 = {1{$random}};
    R571 = {2{$random}};
    R579 = {1{$random}};
    R584 = {2{$random}};
    R592 = {1{$random}};
    R597 = {2{$random}};
    R605 = {1{$random}};
    R610 = {2{$random}};
    R618 = {1{$random}};
    R623 = {2{$random}};
    R631 = {1{$random}};
    R636 = {2{$random}};
    R644 = {1{$random}};
    R649 = {2{$random}};
    R657 = {1{$random}};
    R662 = {2{$random}};
    R670 = {1{$random}};
    R675 = {2{$random}};
    R683 = {1{$random}};
    R688 = {2{$random}};
    R696 = {1{$random}};
    R701 = {2{$random}};
    R709 = {1{$random}};
    R714 = {2{$random}};
    R722 = {1{$random}};
    R727 = {2{$random}};
    R735 = {1{$random}};
    R740 = {2{$random}};
    R748 = {1{$random}};
    R753 = {2{$random}};
    R761 = {1{$random}};
    R766 = {2{$random}};
    R774 = {1{$random}};
    R782 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_mscratch = {2{$random}};
    reg_mie_usip = {1{$random}};
    reg_mie_hsip = {1{$random}};
    reg_mie_utip = {1{$random}};
    reg_mie_htip = {1{$random}};
    reg_mip_usip = {1{$random}};
    reg_mip_hsip = {1{$random}};
    reg_mip_utip = {1{$random}};
    reg_mip_htip = {1{$random}};
    host_csr_rep_valid = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_dma_resp_bits_status = {1{$random}};
//  assign io_rocc_dma_resp_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dma_resp_valid = {1{$random}};
//  assign io_rocc_dma_req_ready = {1{$random}};
//  assign io_rocc_exception = {1{$random}};
//  assign io_rocc_fpu_resp_bits_exc = {1{$random}};
//  assign io_rocc_fpu_resp_bits_data = {3{$random}};
//  assign io_rocc_fpu_resp_valid = {1{$random}};
//  assign io_rocc_fpu_req_ready = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_autl_grant_bits_data = {4{$random}};
//  assign io_rocc_autl_grant_bits_g_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_autl_grant_valid = {1{$random}};
//  assign io_rocc_autl_acquire_ready = {1{$random}};
//  assign io_rocc_s = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_rocc_cmd_bits_rs2 = {2{$random}};
//  assign io_rocc_cmd_bits_rs1 = {2{$random}};
//  assign io_rocc_cmd_bits_inst_opcode = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_xd = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs1 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_rs2 = {1{$random}};
//  assign io_rocc_cmd_bits_inst_funct = {1{$random}};
//  assign io_rocc_cmd_valid = {1{$random}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T3 <= 3'h1;
  assign T3 = T883 + T4;
  assign T4 = {1'h0, T5};
  assign T5 = T882 + T6;
  assign T6 = {1'h0, csr_xcpt};
  assign csr_xcpt = T11 | insn_break;
  assign insn_break = T7 & system_insn;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T7 = T9 & T8;
  assign T8 = io_rw_addr[1'h0:1'h0];
  assign T9 = T10 ^ 1'h1;
  assign T10 = io_rw_addr[4'h8:4'h8];
  assign T11 = T17 | insn_call;
  assign insn_call = T12 & system_insn;
  assign T12 = T15 & T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = io_rw_addr[1'h0:1'h0];
  assign T15 = T16 ^ 1'h1;
  assign T16 = io_rw_addr[4'h8:4'h8];
  assign T17 = T94 | T18;
  assign T18 = system_insn & T19;
  assign T19 = priv_sufficient ^ 1'h1;
  assign priv_sufficient = csr_addr_priv <= reg_mstatus_prv;
  assign T20 = reset ? 2'h3 : T21;
  assign T21 = T88 ? T87 : T22;
  assign T22 = insn_redirect_trap ? 2'h1 : T23;
  assign T23 = insn_ret ? reg_mstatus_prv1 : T24;
  assign T24 = T25 ? 2'h3 : reg_mstatus_prv;
  assign T25 = io_exception | csr_xcpt;
  assign T26 = reset ? 2'h3 : T27;
  assign T27 = T76 ? T881 : T28;
  assign T28 = T69 ? T68 : T29;
  assign T29 = insn_ret ? reg_mstatus_prv2 : T30;
  assign T30 = T25 ? reg_mstatus_prv : reg_mstatus_prv1;
  assign T31 = reset ? 2'h0 : T32;
  assign T32 = T52 ? T35 : T33;
  assign T33 = insn_ret ? 2'h0 : T34;
  assign T34 = T25 ? reg_mstatus_prv1 : reg_mstatus_prv2;
  assign T35 = wdata[4'h8:3'h7];
  assign wdata = T51 ? io_rw_wdata : T36;
  assign T36 = T50 ? T48 : T37;
  assign T37 = T47 ? T46 : host_csr_bits_data;
  assign T38 = host_csr_req_fire ? io_rw_rdata : T39;
  assign T39 = T40 ? io_host_csr_req_bits_data : host_csr_bits_data;
  assign T40 = io_host_csr_req_ready & io_host_csr_req_valid;
  assign host_csr_req_fire = host_csr_req_valid & T41;
  assign T41 = cpu_ren ^ 1'h1;
  assign cpu_ren = T43 & T42;
  assign T42 = system_insn ^ 1'h1;
  assign T43 = io_rw_cmd != 3'h0;
  assign T44 = host_csr_req_fire ? 1'h0 : T45;
  assign T45 = T40 ? 1'h1 : host_csr_req_valid;
  assign T46 = io_rw_rdata | io_rw_wdata;
  assign T47 = io_rw_cmd == 3'h2;
  assign T48 = io_rw_rdata & T49;
  assign T49 = ~ io_rw_wdata;
  assign T50 = io_rw_cmd == 3'h3;
  assign T51 = io_rw_cmd == 3'h1;
  assign T52 = T58 & T53;
  assign T53 = T55 | T54;
  assign T54 = 2'h1 == T35;
  assign T55 = T57 | T56;
  assign T56 = 2'h0 == T35;
  assign T57 = 2'h3 == T35;
  assign T58 = wen & T59;
  assign T59 = addr == 12'h300;
  assign addr = cpu_ren ? io_rw_addr : host_csr_bits_addr;
  assign T60 = T40 ? io_host_csr_req_bits_addr : host_csr_bits_addr;
  assign wen = T63 | T61;
  assign T61 = host_csr_req_fire & host_csr_bits_rw;
  assign T62 = T40 ? io_host_csr_req_bits_rw : host_csr_bits_rw;
  assign T63 = cpu_wen & T64;
  assign T64 = read_only ^ 1'h1;
  assign read_only = T65 == 2'h3;
  assign T65 = io_rw_addr[4'hb:4'ha];
  assign cpu_wen = T66 & priv_sufficient;
  assign T66 = cpu_ren & T67;
  assign T67 = io_rw_cmd != 3'h5;
  assign T68 = wdata[3'h5:3'h4];
  assign T69 = T58 & T70;
  assign T70 = T72 | T71;
  assign T71 = 2'h1 == T68;
  assign T72 = T74 | T73;
  assign T73 = 2'h0 == T68;
  assign T74 = 2'h3 == T68;
  assign T881 = {1'h0, T75};
  assign T75 = wdata[3'h4:3'h4];
  assign T76 = wen & T77;
  assign T77 = addr == 12'h100;
  assign insn_ret = T78 & priv_sufficient;
  assign T78 = T79 & system_insn;
  assign T79 = T82 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = io_rw_addr[1'h0:1'h0];
  assign T82 = T85 & T83;
  assign T83 = T84 ^ 1'h1;
  assign T84 = io_rw_addr[1'h1:1'h1];
  assign T85 = io_rw_addr[4'h8:4'h8];
  assign insn_redirect_trap = maybe_insn_redirect_trap & priv_sufficient;
  assign maybe_insn_redirect_trap = T86 & system_insn;
  assign T86 = io_rw_addr[2'h2:2'h2];
  assign T87 = wdata[2'h2:1'h1];
  assign T88 = T58 & T89;
  assign T89 = T91 | T90;
  assign T90 = 2'h1 == T87;
  assign T91 = T93 | T92;
  assign T92 = 2'h0 == T87;
  assign T93 = 2'h3 == T87;
  assign csr_addr_priv = io_rw_addr[4'h9:4'h8];
  assign T94 = T214 | T95;
  assign T95 = cpu_ren & T96;
  assign T96 = T104 | T97;
  assign T97 = fp_csr & T98;
  assign T98 = T99 ^ 1'h1;
  assign T99 = io_status_fs != 2'h0;
  assign fp_csr = T101 | T100;
  assign T100 = addr == 12'h3;
  assign T101 = T103 | T102;
  assign T102 = addr == 12'h2;
  assign T103 = addr == 12'h1;
  assign T104 = T213 | T105;
  assign T105 = addr_valid ^ 1'h1;
  assign addr_valid = T107 | T106;
  assign T106 = addr == 12'h101;
  assign T107 = T109 | T108;
  assign T108 = addr == 12'h141;
  assign T109 = T111 | T110;
  assign T110 = addr == 12'h181;
  assign T111 = T113 | T112;
  assign T112 = addr == 12'h180;
  assign T113 = T115 | T114;
  assign T114 = addr == 12'hd43;
  assign T115 = T117 | T116;
  assign T116 = addr == 12'hd42;
  assign T117 = T119 | T118;
  assign T118 = addr == 12'h140;
  assign T119 = T121 | T120;
  assign T120 = addr == 12'h104;
  assign T121 = T123 | T122;
  assign T122 = addr == 12'h144;
  assign T123 = T124 | T77;
  assign T124 = T126 | T125;
  assign T125 = addr == 12'hccf;
  assign T126 = T128 | T127;
  assign T127 = addr == 12'hcce;
  assign T128 = T130 | T129;
  assign T129 = addr == 12'hccd;
  assign T130 = T132 | T131;
  assign T131 = addr == 12'hccc;
  assign T132 = T134 | T133;
  assign T133 = addr == 12'hccb;
  assign T134 = T136 | T135;
  assign T135 = addr == 12'hcca;
  assign T136 = T138 | T137;
  assign T137 = addr == 12'hcc9;
  assign T138 = T140 | T139;
  assign T139 = addr == 12'hcc8;
  assign T140 = T142 | T141;
  assign T141 = addr == 12'hcc7;
  assign T142 = T144 | T143;
  assign T143 = addr == 12'hcc6;
  assign T144 = T146 | T145;
  assign T145 = addr == 12'hcc5;
  assign T146 = T148 | T147;
  assign T147 = addr == 12'hcc4;
  assign T148 = T150 | T149;
  assign T149 = addr == 12'hcc3;
  assign T150 = T152 | T151;
  assign T151 = addr == 12'hcc2;
  assign T152 = T154 | T153;
  assign T153 = addr == 12'hcc1;
  assign T154 = T156 | T155;
  assign T155 = addr == 12'hcc0;
  assign T156 = T158 | T157;
  assign T157 = addr == 12'h902;
  assign T158 = T160 | T159;
  assign T159 = addr == 12'hc02;
  assign T160 = T162 | T161;
  assign T161 = addr == 12'h781;
  assign T162 = T164 | T163;
  assign T163 = addr == 12'h780;
  assign T164 = T166 | T165;
  assign T165 = addr == 12'hc0;
  assign T166 = T168 | T167;
  assign T167 = addr == 12'hf10;
  assign T168 = T170 | T169;
  assign T169 = addr == 12'h321;
  assign T170 = T172 | T171;
  assign T171 = addr == 12'h342;
  assign T172 = T174 | T173;
  assign T173 = addr == 12'h343;
  assign T174 = T176 | T175;
  assign T175 = addr == 12'h341;
  assign T176 = T178 | T177;
  assign T177 = addr == 12'h340;
  assign T178 = T180 | T179;
  assign T179 = addr == 12'h304;
  assign T180 = T182 | T181;
  assign T181 = addr == 12'h344;
  assign T182 = T184 | T183;
  assign T183 = addr == 12'h783;
  assign T184 = T186 | T185;
  assign T185 = addr == 12'h784;
  assign T186 = T188 | T187;
  assign T187 = addr == 12'h301;
  assign T188 = T190 | T189;
  assign T189 = addr == 12'h782;
  assign T190 = T192 | T191;
  assign T191 = addr == 12'h302;
  assign T192 = T193 | T59;
  assign T193 = T195 | T194;
  assign T194 = addr == 12'hf01;
  assign T195 = T197 | T196;
  assign T196 = addr == 12'hf00;
  assign T197 = T199 | T198;
  assign T198 = addr == 12'h701;
  assign T199 = T201 | T200;
  assign T200 = addr == 12'ha01;
  assign T201 = T203 | T202;
  assign T202 = addr == 12'hd01;
  assign T203 = T205 | T204;
  assign T204 = addr == 12'h901;
  assign T205 = T207 | T206;
  assign T206 = addr == 12'hc01;
  assign T207 = T209 | T208;
  assign T208 = addr == 12'h900;
  assign T209 = T211 | T210;
  assign T210 = addr == 12'hc00;
  assign T211 = T212 | T100;
  assign T212 = T103 | T102;
  assign T213 = priv_sufficient ^ 1'h1;
  assign T214 = cpu_wen & read_only;
  assign T882 = {1'h0, io_exception};
  assign T883 = {1'h0, T215};
  assign T215 = T884 + T216;
  assign T216 = {1'h0, insn_redirect_trap};
  assign T884 = {1'h0, insn_ret};
  assign io_interrupt_cause = T217;
  assign T217 = T298 ? 64'h8000000000000002 : T218;
  assign T218 = T283 ? 64'h8000000000000001 : T219;
  assign T219 = T271 ? 64'h8000000000000001 : T220;
  assign T220 = T259 ? 64'h8000000000000000 : T221;
  assign T221 = T222 ? 64'h8000000000000000 : 64'h0;
  assign T222 = T246 & T223;
  assign T223 = T245 | T224;
  assign T224 = T244 & reg_mstatus_ie;
  assign T225 = reset ? 1'h0 : T226;
  assign T226 = T76 ? T243 : T227;
  assign T227 = T58 ? T242 : T228;
  assign T228 = insn_ret ? reg_mstatus_ie1 : T229;
  assign T229 = T25 ? 1'h0 : reg_mstatus_ie;
  assign T230 = reset ? 1'h0 : T231;
  assign T231 = T76 ? T241 : T232;
  assign T232 = T58 ? T240 : T233;
  assign T233 = insn_ret ? reg_mstatus_ie2 : T234;
  assign T234 = T25 ? reg_mstatus_ie : reg_mstatus_ie1;
  assign T235 = reset ? 1'h0 : T236;
  assign T236 = T58 ? T239 : T237;
  assign T237 = insn_ret ? 1'h1 : T238;
  assign T238 = T25 ? reg_mstatus_ie1 : reg_mstatus_ie2;
  assign T239 = wdata[3'h6:3'h6];
  assign T240 = wdata[2'h3:2'h3];
  assign T241 = wdata[2'h3:2'h3];
  assign T242 = wdata[1'h0:1'h0];
  assign T243 = wdata[1'h0:1'h0];
  assign T244 = reg_mstatus_prv == 2'h1;
  assign T245 = reg_mstatus_prv < 2'h1;
  assign T246 = reg_mie_ssip & reg_mip_ssip;
  assign T885 = reset ? 1'h0 : T247;
  assign T247 = T252 ? T251 : T248;
  assign T248 = T250 ? T249 : reg_mip_ssip;
  assign T249 = wdata[1'h1:1'h1];
  assign T250 = wen & T181;
  assign T251 = wdata[1'h1:1'h1];
  assign T252 = wen & T122;
  assign T886 = reset ? 1'h0 : T253;
  assign T253 = T258 ? T257 : T254;
  assign T254 = T256 ? T255 : reg_mie_ssip;
  assign T255 = wdata[1'h1:1'h1];
  assign T256 = wen & T179;
  assign T257 = wdata[1'h1:1'h1];
  assign T258 = wen & T120;
  assign T259 = T264 & T260;
  assign T260 = T263 | T261;
  assign T261 = T262 & reg_mstatus_ie;
  assign T262 = reg_mstatus_prv == 2'h3;
  assign T263 = reg_mstatus_prv < 2'h3;
  assign T264 = reg_mie_msip & reg_mip_msip;
  assign T887 = reset ? 1'h0 : T265;
  assign T265 = T268 ? 1'h1 : T266;
  assign T266 = T250 ? T267 : reg_mip_msip;
  assign T267 = wdata[2'h3:2'h3];
  assign T268 = wen & T183;
  assign T888 = reset ? 1'h0 : T269;
  assign T269 = T256 ? T270 : reg_mie_msip;
  assign T270 = wdata[2'h3:2'h3];
  assign T271 = T276 & T272;
  assign T272 = T275 | T273;
  assign T273 = T274 & reg_mstatus_ie;
  assign T274 = reg_mstatus_prv == 2'h1;
  assign T275 = reg_mstatus_prv < 2'h1;
  assign T276 = reg_mie_stip & reg_mip_stip;
  assign T889 = reset ? 1'h0 : T277;
  assign T277 = T250 ? T278 : reg_mip_stip;
  assign T278 = wdata[3'h5:3'h5];
  assign T890 = reset ? 1'h0 : T279;
  assign T279 = T258 ? T282 : T280;
  assign T280 = T256 ? T281 : reg_mie_stip;
  assign T281 = wdata[3'h5:3'h5];
  assign T282 = wdata[3'h5:3'h5];
  assign T283 = T288 & T284;
  assign T284 = T287 | T285;
  assign T285 = T286 & reg_mstatus_ie;
  assign T286 = reg_mstatus_prv == 2'h3;
  assign T287 = reg_mstatus_prv < 2'h3;
  assign T288 = reg_mie_mtip & reg_mip_mtip;
  assign T891 = reset ? 1'h0 : T289;
  assign T289 = T295 ? 1'h0 : T290;
  assign T290 = T291 ? 1'h1 : reg_mip_mtip;
  assign T291 = reg_mtimecmp <= read_time;
  assign T292 = T293 ? wdata : read_time;
  assign T293 = wen & T198;
  assign T294 = T295 ? wdata : reg_mtimecmp;
  assign T295 = wen & T169;
  assign T892 = reset ? 1'h0 : T296;
  assign T296 = T256 ? T297 : reg_mie_mtip;
  assign T297 = wdata[3'h7:3'h7];
  assign T298 = T303 & T299;
  assign T299 = T302 | T300;
  assign T300 = T301 & reg_mstatus_ie;
  assign T301 = reg_mstatus_prv == 2'h3;
  assign T302 = reg_mstatus_prv < 2'h3;
  assign T303 = reg_fromhost != 64'h0;
  assign T893 = reset ? 64'h0 : T304;
  assign T304 = T305 ? wdata : reg_fromhost;
  assign T305 = T309 & T306;
  assign T306 = T308 | T307;
  assign T307 = host_csr_req_fire ^ 1'h1;
  assign T308 = reg_fromhost == 64'h0;
  assign T309 = wen & T161;
  assign io_interrupt = T310;
  assign T310 = io_interrupt_cause[6'h3f:6'h3f];
  assign io_fcsr_rm = reg_frm;
  assign T894 = T311[2'h2:1'h0];
  assign T311 = T315 ? T896 : T312;
  assign T312 = T313 ? wdata : T895;
  assign T895 = {61'h0, reg_frm};
  assign T313 = wen & T102;
  assign T896 = {5'h0, T314};
  assign T314 = wdata >> 3'h5;
  assign T315 = wen & T100;
  assign io_time = T316;
  assign T316 = {R320, R317};
  assign T897 = reset ? 6'h0 : T318;
  assign T318 = T319[3'h5:1'h0];
  assign T319 = T898 + 7'h1;
  assign T898 = {1'h0, R317};
  assign T899 = reset ? 58'h0 : T321;
  assign T321 = T323 ? T322 : R320;
  assign T322 = R320 + 58'h1;
  assign T323 = T319[3'h6:3'h6];
  assign io_fatc = insn_sfence_vm;
  assign insn_sfence_vm = T324 & priv_sufficient;
  assign T324 = T325 & system_insn;
  assign T325 = T327 & T326;
  assign T326 = io_rw_addr[1'h0:1'h0];
  assign T327 = T330 & T328;
  assign T328 = T329 ^ 1'h1;
  assign T329 = io_rw_addr[1'h1:1'h1];
  assign T330 = io_rw_addr[4'h8:4'h8];
  assign io_evec = T331;
  assign T331 = T359 ? T906 : T332;
  assign T332 = maybe_insn_redirect_trap ? T350 : T333;
  assign T333 = T349 ? reg_mepc : reg_sepc;
  assign T900 = T334[6'h27:1'h0];
  assign T334 = T339 ? T336 : T901;
  assign T901 = {24'h0, T335};
  assign T335 = insn_redirect_trap ? reg_mepc : reg_sepc;
  assign T336 = ~ T337;
  assign T337 = T338 | 64'h3;
  assign T338 = ~ wdata;
  assign T339 = wen & T108;
  assign T902 = T340[6'h27:1'h0];
  assign T340 = T348 ? T345 : T903;
  assign T903 = {24'h0, T341};
  assign T341 = T25 ? T342 : reg_mepc;
  assign T342 = ~ T343;
  assign T343 = T344 | 40'h3;
  assign T344 = ~ io_pc;
  assign T345 = ~ T346;
  assign T346 = T347 | 64'h3;
  assign T347 = ~ wdata;
  assign T348 = wen & T175;
  assign T349 = reg_mstatus_prv[1'h1:1'h1];
  assign T350 = {T356, reg_stvec};
  assign T904 = T351[6'h26:1'h0];
  assign T351 = T355 ? T352 : T905;
  assign T905 = {25'h0, reg_stvec};
  assign T352 = ~ T353;
  assign T353 = T354 | 64'h3;
  assign T354 = ~ wdata;
  assign T355 = wen & T106;
  assign T356 = reg_stvec[6'h26:6'h26];
  assign T906 = {31'h0, T357};
  assign T357 = T907 + 9'h100;
  assign T907 = {1'h0, T358};
  assign T358 = reg_mstatus_prv << 3'h6;
  assign T359 = io_exception | csr_xcpt;
  assign io_ptbr = reg_sptbr;
  assign T360 = T363 ? T361 : reg_sptbr;
  assign T361 = {T362, 12'h0};
  assign T362 = wdata[5'h1f:4'hc];
  assign T363 = wen & T112;
  assign io_status_ie = reg_mstatus_ie;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_ie1 = reg_mstatus_ie1;
  assign io_status_prv1 = reg_mstatus_prv1;
  assign io_status_ie2 = reg_mstatus_ie2;
  assign io_status_prv2 = reg_mstatus_prv2;
  assign io_status_ie3 = reg_mstatus_ie3;
  assign T364 = reset ? 1'h0 : reg_mstatus_ie3;
  assign io_status_prv3 = reg_mstatus_prv3;
  assign T365 = reset ? 2'h0 : reg_mstatus_prv3;
  assign io_status_fs = T366;
  assign T366 = 2'h0 - T908;
  assign T908 = {1'h0, T367};
  assign T367 = reg_mstatus_fs != 2'h0;
  assign T368 = reset ? 2'h0 : T369;
  assign T369 = T76 ? T372 : T370;
  assign T370 = T58 ? T371 : reg_mstatus_fs;
  assign T371 = wdata[4'hd:4'hc];
  assign T372 = wdata[4'hd:4'hc];
  assign io_status_xs = T373;
  assign T373 = 2'h0 - T909;
  assign T909 = {1'h0, T374};
  assign T374 = reg_mstatus_xs != 2'h0;
  assign T375 = reset ? 2'h0 : reg_mstatus_xs;
  assign io_status_mprv = reg_mstatus_mprv;
  assign T376 = reset ? 1'h0 : T377;
  assign T377 = T76 ? T381 : T378;
  assign T378 = T58 ? T380 : T379;
  assign T379 = T25 ? 1'h0 : reg_mstatus_mprv;
  assign T380 = wdata[5'h10:5'h10];
  assign T381 = wdata[5'h10:5'h10];
  assign io_status_vm = reg_mstatus_vm;
  assign T382 = reset ? 5'h0 : T383;
  assign T383 = T388 ? 5'h9 : T384;
  assign T384 = T385 ? 5'h0 : reg_mstatus_vm;
  assign T385 = T58 & T386;
  assign T386 = T387 == 5'h0;
  assign T387 = wdata[5'h15:5'h11];
  assign T388 = T58 & T389;
  assign T389 = T387 == 5'h9;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign T390 = reset ? 9'h0 : reg_mstatus_zero1;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign T391 = reset ? 1'h0 : reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign T392 = reset ? 31'h0 : reg_mstatus_zero2;
  assign io_status_sd = T393;
  assign T393 = T395 | T394;
  assign T394 = io_status_xs == 2'h3;
  assign T395 = io_status_fs == 2'h3;
  assign io_eret = T396;
  assign T396 = insn_ret | insn_redirect_trap;
  assign io_csr_xcpt = csr_xcpt;
  assign io_csr_stall = reg_wfi;
  assign T910 = reset ? 1'h0 : T397;
  assign T397 = some_interrupt_pending ? 1'h0 : T398;
  assign T398 = insn_wfi ? 1'h1 : reg_wfi;
  assign insn_wfi = T399 & priv_sufficient;
  assign T399 = T400 & system_insn;
  assign T400 = T403 & T401;
  assign T401 = T402 ^ 1'h1;
  assign T402 = io_rw_addr[1'h0:1'h0];
  assign T403 = T405 & T404;
  assign T404 = io_rw_addr[1'h1:1'h1];
  assign T405 = io_rw_addr[4'h8:4'h8];
  assign some_interrupt_pending = T406;
  assign T406 = T418 ? 1'h1 : T407;
  assign T407 = T416 ? 1'h1 : T408;
  assign T408 = T414 ? 1'h1 : T409;
  assign T409 = T412 ? 1'h1 : T410;
  assign T410 = T246 & T411;
  assign T411 = reg_mstatus_prv <= 2'h1;
  assign T412 = T264 & T413;
  assign T413 = reg_mstatus_prv <= 2'h3;
  assign T414 = T276 & T415;
  assign T415 = reg_mstatus_prv <= 2'h1;
  assign T416 = T288 & T417;
  assign T417 = reg_mstatus_prv <= 2'h3;
  assign T418 = T303 & T419;
  assign T419 = reg_mstatus_prv <= 2'h3;
  assign io_rw_rdata = T420;
  assign T420 = T425 | T421;
  assign T421 = T106 ? T422 : 64'h0;
  assign T422 = {T423, reg_stvec};
  assign T423 = 25'h0 - T911;
  assign T911 = {24'h0, T424};
  assign T424 = reg_stvec[6'h26:6'h26];
  assign T425 = T430 | T426;
  assign T426 = T108 ? T427 : 64'h0;
  assign T427 = {T428, reg_sepc};
  assign T428 = 24'h0 - T912;
  assign T912 = {23'h0, T429};
  assign T429 = reg_sepc[6'h27:6'h27];
  assign T430 = T431 | 64'h0;
  assign T431 = T433 | T913;
  assign T913 = {32'h0, T432};
  assign T432 = T112 ? reg_sptbr : 32'h0;
  assign T433 = T460 | T434;
  assign T434 = T114 ? T435 : 64'h0;
  assign T435 = {T458, reg_sbadaddr};
  assign T436 = insn_redirect_trap ? reg_mbadaddr : reg_sbadaddr;
  assign T437 = T457 ? T456 : T438;
  assign T438 = T448 ? T440 : T439;
  assign T439 = T25 ? io_pc : reg_mbadaddr;
  assign T440 = {T442, T441};
  assign T441 = io_rw_wdata[6'h26:1'h0];
  assign T442 = T446 ? T445 : T443;
  assign T443 = T444 != 25'h0;
  assign T444 = io_rw_wdata[6'h3f:6'h27];
  assign T445 = T444 == 25'h1ffffff;
  assign T446 = $signed(T447) < $signed(1'h0);
  assign T447 = T441;
  assign T448 = T25 & T449;
  assign T449 = T451 | T450;
  assign T450 = io_cause == 64'h6;
  assign T451 = T453 | T452;
  assign T452 = io_cause == 64'h7;
  assign T453 = T455 | T454;
  assign T454 = io_cause == 64'h4;
  assign T455 = io_cause == 64'h5;
  assign T456 = wdata[6'h27:1'h0];
  assign T457 = wen & T173;
  assign T458 = 24'h0 - T914;
  assign T914 = {23'h0, T459};
  assign T459 = reg_sbadaddr[6'h27:6'h27];
  assign T460 = T474 | T461;
  assign T461 = T116 ? reg_scause : 64'h0;
  assign T462 = insn_redirect_trap ? reg_mcause : reg_scause;
  assign T463 = T473 ? T472 : T464;
  assign T464 = T471 ? T915 : T465;
  assign T465 = T469 ? 64'h3 : T466;
  assign T466 = T468 ? 64'h2 : T467;
  assign T467 = T25 ? io_cause : reg_mcause;
  assign T468 = T25 & csr_xcpt;
  assign T469 = T468 & insn_break;
  assign T915 = {60'h0, T470};
  assign T470 = T916 + 4'h8;
  assign T916 = {2'h0, reg_mstatus_prv};
  assign T471 = T468 & insn_call;
  assign T472 = wdata & 64'h800000000000001f;
  assign T473 = wen & T171;
  assign T474 = T478 | T475;
  assign T475 = T118 ? reg_sscratch : 64'h0;
  assign T476 = T477 ? wdata : reg_sscratch;
  assign T477 = wen & T118;
  assign T478 = T496 | T917;
  assign T917 = {56'h0, T479};
  assign T479 = T120 ? T480 : 8'h0;
  assign T480 = T481;
  assign T481 = {T489, T482};
  assign T482 = {T486, T483};
  assign T483 = {T485, T484};
  assign T484 = 1'h0;
  assign T485 = reg_mie_ssip;
  assign T486 = {T488, T487};
  assign T487 = 1'h0;
  assign T488 = 1'h0;
  assign T489 = {T493, T490};
  assign T490 = {T492, T491};
  assign T491 = 1'h0;
  assign T492 = reg_mie_stip;
  assign T493 = {T495, T494};
  assign T494 = 1'h0;
  assign T495 = 1'h0;
  assign T496 = T514 | T918;
  assign T918 = {56'h0, T497};
  assign T497 = T122 ? T498 : 8'h0;
  assign T498 = T499;
  assign T499 = {T507, T500};
  assign T500 = {T504, T501};
  assign T501 = {T503, T502};
  assign T502 = 1'h0;
  assign T503 = reg_mip_ssip;
  assign T504 = {T506, T505};
  assign T505 = 1'h0;
  assign T506 = 1'h0;
  assign T507 = {T511, T508};
  assign T508 = {T510, T509};
  assign T509 = 1'h0;
  assign T510 = reg_mip_stip;
  assign T511 = {T513, T512};
  assign T512 = 1'h0;
  assign T513 = 1'h0;
  assign T514 = T563 | T515;
  assign T515 = T77 ? T516 : 64'h0;
  assign T516 = T517;
  assign T517 = {T548, T518};
  assign T518 = {T541, T519};
  assign T519 = {T539, T520};
  assign T520 = {T538, T521};
  assign T521 = T522;
  assign T522 = read_mstatus[1'h0:1'h0];
  assign read_mstatus = T523;
  assign T523 = {T531, T524};
  assign T524 = {T528, T525};
  assign T525 = {T527, T526};
  assign T526 = {io_status_prv, io_status_ie};
  assign T527 = {io_status_prv1, io_status_ie1};
  assign T528 = {T530, T529};
  assign T529 = {io_status_prv2, io_status_ie2};
  assign T530 = {io_status_prv3, io_status_ie3};
  assign T531 = {T535, T532};
  assign T532 = {T534, T533};
  assign T533 = {io_status_xs, io_status_fs};
  assign T534 = {io_status_vm, io_status_mprv};
  assign T535 = {T537, T536};
  assign T536 = {io_status_sd_rv32, io_status_zero1};
  assign T537 = {io_status_sd, io_status_zero2};
  assign T538 = 2'h0;
  assign T539 = T540;
  assign T540 = read_mstatus[2'h3:2'h3];
  assign T541 = {T546, T542};
  assign T542 = {T545, T543};
  assign T543 = T544;
  assign T544 = read_mstatus[3'h4:3'h4];
  assign T545 = 7'h0;
  assign T546 = T547;
  assign T547 = read_mstatus[4'hd:4'hc];
  assign T548 = {T556, T549};
  assign T549 = {T555, T550};
  assign T550 = {T553, T551};
  assign T551 = T552;
  assign T552 = read_mstatus[4'hf:4'he];
  assign T553 = T554;
  assign T554 = read_mstatus[5'h10:5'h10];
  assign T555 = 14'h0;
  assign T556 = {T561, T557};
  assign T557 = {T560, T558};
  assign T558 = T559;
  assign T559 = read_mstatus[5'h1f:5'h1f];
  assign T560 = 31'h0;
  assign T561 = T562;
  assign T562 = read_mstatus[6'h3f:6'h3f];
  assign T563 = T576 | T564;
  assign T564 = T125 ? T565 : 64'h0;
  assign T565 = {R571, R566};
  assign T919 = reset ? 6'h0 : T567;
  assign T567 = T570 ? T568 : R566;
  assign T568 = T569[3'h5:1'h0];
  assign T569 = T920 + 7'h1;
  assign T920 = {1'h0, R566};
  assign T570 = io_uarch_counters_15 != 1'h0;
  assign T921 = reset ? 58'h0 : T572;
  assign T572 = T574 ? T573 : R571;
  assign T573 = R571 + 58'h1;
  assign T574 = T570 & T575;
  assign T575 = T569[3'h6:3'h6];
  assign T576 = T589 | T577;
  assign T577 = T127 ? T578 : 64'h0;
  assign T578 = {R584, R579};
  assign T922 = reset ? 6'h0 : T580;
  assign T580 = T583 ? T581 : R579;
  assign T581 = T582[3'h5:1'h0];
  assign T582 = T923 + 7'h1;
  assign T923 = {1'h0, R579};
  assign T583 = io_uarch_counters_14 != 1'h0;
  assign T924 = reset ? 58'h0 : T585;
  assign T585 = T587 ? T586 : R584;
  assign T586 = R584 + 58'h1;
  assign T587 = T583 & T588;
  assign T588 = T582[3'h6:3'h6];
  assign T589 = T602 | T590;
  assign T590 = T129 ? T591 : 64'h0;
  assign T591 = {R597, R592};
  assign T925 = reset ? 6'h0 : T593;
  assign T593 = T596 ? T594 : R592;
  assign T594 = T595[3'h5:1'h0];
  assign T595 = T926 + 7'h1;
  assign T926 = {1'h0, R592};
  assign T596 = io_uarch_counters_13 != 1'h0;
  assign T927 = reset ? 58'h0 : T598;
  assign T598 = T600 ? T599 : R597;
  assign T599 = R597 + 58'h1;
  assign T600 = T596 & T601;
  assign T601 = T595[3'h6:3'h6];
  assign T602 = T615 | T603;
  assign T603 = T131 ? T604 : 64'h0;
  assign T604 = {R610, R605};
  assign T928 = reset ? 6'h0 : T606;
  assign T606 = T609 ? T607 : R605;
  assign T607 = T608[3'h5:1'h0];
  assign T608 = T929 + 7'h1;
  assign T929 = {1'h0, R605};
  assign T609 = io_uarch_counters_12 != 1'h0;
  assign T930 = reset ? 58'h0 : T611;
  assign T611 = T613 ? T612 : R610;
  assign T612 = R610 + 58'h1;
  assign T613 = T609 & T614;
  assign T614 = T608[3'h6:3'h6];
  assign T615 = T628 | T616;
  assign T616 = T133 ? T617 : 64'h0;
  assign T617 = {R623, R618};
  assign T931 = reset ? 6'h0 : T619;
  assign T619 = T622 ? T620 : R618;
  assign T620 = T621[3'h5:1'h0];
  assign T621 = T932 + 7'h1;
  assign T932 = {1'h0, R618};
  assign T622 = io_uarch_counters_11 != 1'h0;
  assign T933 = reset ? 58'h0 : T624;
  assign T624 = T626 ? T625 : R623;
  assign T625 = R623 + 58'h1;
  assign T626 = T622 & T627;
  assign T627 = T621[3'h6:3'h6];
  assign T628 = T641 | T629;
  assign T629 = T135 ? T630 : 64'h0;
  assign T630 = {R636, R631};
  assign T934 = reset ? 6'h0 : T632;
  assign T632 = T635 ? T633 : R631;
  assign T633 = T634[3'h5:1'h0];
  assign T634 = T935 + 7'h1;
  assign T935 = {1'h0, R631};
  assign T635 = io_uarch_counters_10 != 1'h0;
  assign T936 = reset ? 58'h0 : T637;
  assign T637 = T639 ? T638 : R636;
  assign T638 = R636 + 58'h1;
  assign T639 = T635 & T640;
  assign T640 = T634[3'h6:3'h6];
  assign T641 = T654 | T642;
  assign T642 = T137 ? T643 : 64'h0;
  assign T643 = {R649, R644};
  assign T937 = reset ? 6'h0 : T645;
  assign T645 = T648 ? T646 : R644;
  assign T646 = T647[3'h5:1'h0];
  assign T647 = T938 + 7'h1;
  assign T938 = {1'h0, R644};
  assign T648 = io_uarch_counters_9 != 1'h0;
  assign T939 = reset ? 58'h0 : T650;
  assign T650 = T652 ? T651 : R649;
  assign T651 = R649 + 58'h1;
  assign T652 = T648 & T653;
  assign T653 = T647[3'h6:3'h6];
  assign T654 = T667 | T655;
  assign T655 = T139 ? T656 : 64'h0;
  assign T656 = {R662, R657};
  assign T940 = reset ? 6'h0 : T658;
  assign T658 = T661 ? T659 : R657;
  assign T659 = T660[3'h5:1'h0];
  assign T660 = T941 + 7'h1;
  assign T941 = {1'h0, R657};
  assign T661 = io_uarch_counters_8 != 1'h0;
  assign T942 = reset ? 58'h0 : T663;
  assign T663 = T665 ? T664 : R662;
  assign T664 = R662 + 58'h1;
  assign T665 = T661 & T666;
  assign T666 = T660[3'h6:3'h6];
  assign T667 = T680 | T668;
  assign T668 = T141 ? T669 : 64'h0;
  assign T669 = {R675, R670};
  assign T943 = reset ? 6'h0 : T671;
  assign T671 = T674 ? T672 : R670;
  assign T672 = T673[3'h5:1'h0];
  assign T673 = T944 + 7'h1;
  assign T944 = {1'h0, R670};
  assign T674 = io_uarch_counters_7 != 1'h0;
  assign T945 = reset ? 58'h0 : T676;
  assign T676 = T678 ? T677 : R675;
  assign T677 = R675 + 58'h1;
  assign T678 = T674 & T679;
  assign T679 = T673[3'h6:3'h6];
  assign T680 = T693 | T681;
  assign T681 = T143 ? T682 : 64'h0;
  assign T682 = {R688, R683};
  assign T946 = reset ? 6'h0 : T684;
  assign T684 = T687 ? T685 : R683;
  assign T685 = T686[3'h5:1'h0];
  assign T686 = T947 + 7'h1;
  assign T947 = {1'h0, R683};
  assign T687 = io_uarch_counters_6 != 1'h0;
  assign T948 = reset ? 58'h0 : T689;
  assign T689 = T691 ? T690 : R688;
  assign T690 = R688 + 58'h1;
  assign T691 = T687 & T692;
  assign T692 = T686[3'h6:3'h6];
  assign T693 = T706 | T694;
  assign T694 = T145 ? T695 : 64'h0;
  assign T695 = {R701, R696};
  assign T949 = reset ? 6'h0 : T697;
  assign T697 = T700 ? T698 : R696;
  assign T698 = T699[3'h5:1'h0];
  assign T699 = T950 + 7'h1;
  assign T950 = {1'h0, R696};
  assign T700 = io_uarch_counters_5 != 1'h0;
  assign T951 = reset ? 58'h0 : T702;
  assign T702 = T704 ? T703 : R701;
  assign T703 = R701 + 58'h1;
  assign T704 = T700 & T705;
  assign T705 = T699[3'h6:3'h6];
  assign T706 = T719 | T707;
  assign T707 = T147 ? T708 : 64'h0;
  assign T708 = {R714, R709};
  assign T952 = reset ? 6'h0 : T710;
  assign T710 = T713 ? T711 : R709;
  assign T711 = T712[3'h5:1'h0];
  assign T712 = T953 + 7'h1;
  assign T953 = {1'h0, R709};
  assign T713 = io_uarch_counters_4 != 1'h0;
  assign T954 = reset ? 58'h0 : T715;
  assign T715 = T717 ? T716 : R714;
  assign T716 = R714 + 58'h1;
  assign T717 = T713 & T718;
  assign T718 = T712[3'h6:3'h6];
  assign T719 = T732 | T720;
  assign T720 = T149 ? T721 : 64'h0;
  assign T721 = {R727, R722};
  assign T955 = reset ? 6'h0 : T723;
  assign T723 = T726 ? T724 : R722;
  assign T724 = T725[3'h5:1'h0];
  assign T725 = T956 + 7'h1;
  assign T956 = {1'h0, R722};
  assign T726 = io_uarch_counters_3 != 1'h0;
  assign T957 = reset ? 58'h0 : T728;
  assign T728 = T730 ? T729 : R727;
  assign T729 = R727 + 58'h1;
  assign T730 = T726 & T731;
  assign T731 = T725[3'h6:3'h6];
  assign T732 = T745 | T733;
  assign T733 = T151 ? T734 : 64'h0;
  assign T734 = {R740, R735};
  assign T958 = reset ? 6'h0 : T736;
  assign T736 = T739 ? T737 : R735;
  assign T737 = T738[3'h5:1'h0];
  assign T738 = T959 + 7'h1;
  assign T959 = {1'h0, R735};
  assign T739 = io_uarch_counters_2 != 1'h0;
  assign T960 = reset ? 58'h0 : T741;
  assign T741 = T743 ? T742 : R740;
  assign T742 = R740 + 58'h1;
  assign T743 = T739 & T744;
  assign T744 = T738[3'h6:3'h6];
  assign T745 = T758 | T746;
  assign T746 = T153 ? T747 : 64'h0;
  assign T747 = {R753, R748};
  assign T961 = reset ? 6'h0 : T749;
  assign T749 = T752 ? T750 : R748;
  assign T750 = T751[3'h5:1'h0];
  assign T751 = T962 + 7'h1;
  assign T962 = {1'h0, R748};
  assign T752 = io_uarch_counters_1 != 1'h0;
  assign T963 = reset ? 58'h0 : T754;
  assign T754 = T756 ? T755 : R753;
  assign T755 = R753 + 58'h1;
  assign T756 = T752 & T757;
  assign T757 = T751[3'h6:3'h6];
  assign T758 = T771 | T759;
  assign T759 = T155 ? T760 : 64'h0;
  assign T760 = {R766, R761};
  assign T964 = reset ? 6'h0 : T762;
  assign T762 = T765 ? T763 : R761;
  assign T763 = T764[3'h5:1'h0];
  assign T764 = T965 + 7'h1;
  assign T965 = {1'h0, R761};
  assign T765 = io_uarch_counters_0 != 1'h0;
  assign T966 = reset ? 58'h0 : T767;
  assign T767 = T769 ? T768 : R766;
  assign T768 = R766 + 58'h1;
  assign T769 = T765 & T770;
  assign T770 = T764[3'h6:3'h6];
  assign T771 = T789 | T772;
  assign T772 = T157 ? T773 : 64'h0;
  assign T773 = {R782, R774};
  assign T967 = reset ? 6'h0 : T775;
  assign T775 = T781 ? T780 : T776;
  assign T776 = T779 ? T777 : R774;
  assign T777 = T778[3'h5:1'h0];
  assign T778 = T968 + 7'h1;
  assign T968 = {1'h0, R774};
  assign T779 = io_retire != 1'h0;
  assign T780 = wdata[3'h5:1'h0];
  assign T781 = wen & T157;
  assign T969 = reset ? 58'h0 : T783;
  assign T783 = T781 ? T788 : T784;
  assign T784 = T786 ? T785 : R782;
  assign T785 = R782 + 58'h1;
  assign T786 = T779 & T787;
  assign T787 = T778[3'h6:3'h6];
  assign T788 = wdata[6'h3f:3'h6];
  assign T789 = T791 | T790;
  assign T790 = T159 ? T773 : 64'h0;
  assign T791 = T793 | T792;
  assign T792 = T161 ? reg_fromhost : 64'h0;
  assign T793 = T804 | T794;
  assign T794 = T163 ? reg_tohost : 64'h0;
  assign T970 = reset ? 64'h0 : T795;
  assign T795 = T800 ? wdata : T796;
  assign T796 = T797 ? 64'h0 : reg_tohost;
  assign T797 = T798 & T163;
  assign T798 = host_csr_req_fire & T799;
  assign T799 = host_csr_bits_rw ^ 1'h1;
  assign T800 = T803 & T801;
  assign T801 = T802 | host_csr_req_fire;
  assign T802 = reg_tohost == 64'h0;
  assign T803 = wen & T163;
  assign T804 = T809 | T971;
  assign T971 = {63'h0, T805};
  assign T805 = T165 ? reg_stats : 1'h0;
  assign T972 = reset ? 1'h0 : T806;
  assign T806 = T808 ? T807 : reg_stats;
  assign T807 = wdata[1'h0:1'h0];
  assign T808 = wen & T165;
  assign T809 = T811 | T973;
  assign T973 = {63'h0, T810};
  assign T810 = T167 ? io_host_id : 1'h0;
  assign T811 = T813 | T812;
  assign T812 = T169 ? reg_mtimecmp : 64'h0;
  assign T813 = T815 | T814;
  assign T814 = T171 ? reg_mcause : 64'h0;
  assign T815 = T820 | T816;
  assign T816 = T173 ? T817 : 64'h0;
  assign T817 = {T818, reg_mbadaddr};
  assign T818 = 24'h0 - T974;
  assign T974 = {23'h0, T819};
  assign T819 = reg_mbadaddr[6'h27:6'h27];
  assign T820 = T825 | T821;
  assign T821 = T175 ? T822 : 64'h0;
  assign T822 = {T823, reg_mepc};
  assign T823 = 24'h0 - T975;
  assign T975 = {23'h0, T824};
  assign T824 = reg_mepc[6'h27:6'h27];
  assign T825 = T829 | T826;
  assign T826 = T177 ? reg_mscratch : 64'h0;
  assign T827 = T828 ? wdata : reg_mscratch;
  assign T828 = wen & T177;
  assign T829 = T839 | T976;
  assign T976 = {56'h0, T830};
  assign T830 = T179 ? T831 : 8'h0;
  assign T831 = T832;
  assign T832 = {T836, T833};
  assign T833 = {T835, T834};
  assign T834 = {reg_mie_ssip, reg_mie_usip};
  assign T977 = reset ? 1'h0 : reg_mie_usip;
  assign T835 = {reg_mie_msip, reg_mie_hsip};
  assign T978 = reset ? 1'h0 : reg_mie_hsip;
  assign T836 = {T838, T837};
  assign T837 = {reg_mie_stip, reg_mie_utip};
  assign T979 = reset ? 1'h0 : reg_mie_utip;
  assign T838 = {reg_mie_mtip, reg_mie_htip};
  assign T980 = reset ? 1'h0 : reg_mie_htip;
  assign T839 = T849 | T981;
  assign T981 = {56'h0, T840};
  assign T840 = T181 ? T841 : 8'h0;
  assign T841 = T842;
  assign T842 = {T846, T843};
  assign T843 = {T845, T844};
  assign T844 = {reg_mip_ssip, reg_mip_usip};
  assign T982 = reset ? 1'h0 : reg_mip_usip;
  assign T845 = {reg_mip_msip, reg_mip_hsip};
  assign T983 = reset ? 1'h0 : reg_mip_hsip;
  assign T846 = {T848, T847};
  assign T847 = {reg_mip_stip, reg_mip_utip};
  assign T984 = reset ? 1'h0 : reg_mip_utip;
  assign T848 = {reg_mip_mtip, reg_mip_htip};
  assign T985 = reset ? 1'h0 : reg_mip_htip;
  assign T849 = T850 | 64'h0;
  assign T850 = T852 | T986;
  assign T986 = {33'h0, T851};
  assign T851 = T185 ? 31'h40000000 : 31'h0;
  assign T852 = T854 | T987;
  assign T987 = {55'h0, T853};
  assign T853 = T187 ? 9'h100 : 9'h0;
  assign T854 = T855 | 64'h0;
  assign T855 = T856 | 64'h0;
  assign T856 = T858 | T857;
  assign T857 = T59 ? read_mstatus : 64'h0;
  assign T858 = T859 | T988;
  assign T988 = {63'h0, T194};
  assign T859 = T861 | T860;
  assign T860 = T196 ? 64'h8000000000041101 : 64'h0;
  assign T861 = T863 | T862;
  assign T862 = T198 ? read_time : 64'h0;
  assign T863 = T865 | T864;
  assign T864 = T200 ? read_time : 64'h0;
  assign T865 = T867 | T866;
  assign T866 = T202 ? read_time : 64'h0;
  assign T867 = T869 | T868;
  assign T868 = T204 ? read_time : 64'h0;
  assign T869 = T871 | T870;
  assign T870 = T206 ? read_time : 64'h0;
  assign T871 = T873 | T872;
  assign T872 = T208 ? T316 : 64'h0;
  assign T873 = 64'h0 | T874;
  assign T874 = T210 ? T316 : 64'h0;
  assign io_host_debug_stats_csr = reg_stats;
  assign io_host_csr_resp_bits = host_csr_bits_data;
  assign io_host_csr_resp_valid = host_csr_rep_valid;
  assign T875 = T877 ? 1'h0 : T876;
  assign T876 = host_csr_req_fire ? 1'h1 : host_csr_rep_valid;
  assign T877 = io_host_csr_resp_ready & io_host_csr_resp_valid;
  assign io_host_csr_req_ready = T878;
  assign T878 = T880 & T879;
  assign T879 = host_csr_rep_valid ^ 1'h1;
  assign T880 = host_csr_req_valid ^ 1'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "these conditions must be mutually exclusive");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      reg_mstatus_prv <= 2'h3;
    end else if(T88) begin
      reg_mstatus_prv <= T87;
    end else if(insn_redirect_trap) begin
      reg_mstatus_prv <= 2'h1;
    end else if(insn_ret) begin
      reg_mstatus_prv <= reg_mstatus_prv1;
    end else if(T25) begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_prv1 <= 2'h3;
    end else if(T76) begin
      reg_mstatus_prv1 <= T881;
    end else if(T69) begin
      reg_mstatus_prv1 <= T68;
    end else if(insn_ret) begin
      reg_mstatus_prv1 <= reg_mstatus_prv2;
    end else if(T25) begin
      reg_mstatus_prv1 <= reg_mstatus_prv;
    end
    if(reset) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T52) begin
      reg_mstatus_prv2 <= T35;
    end else if(insn_ret) begin
      reg_mstatus_prv2 <= 2'h0;
    end else if(T25) begin
      reg_mstatus_prv2 <= reg_mstatus_prv1;
    end
    if(host_csr_req_fire) begin
      host_csr_bits_data <= io_rw_rdata;
    end else if(T40) begin
      host_csr_bits_data <= io_host_csr_req_bits_data;
    end
    if(host_csr_req_fire) begin
      host_csr_req_valid <= 1'h0;
    end else if(T40) begin
      host_csr_req_valid <= 1'h1;
    end
    if(T40) begin
      host_csr_bits_addr <= io_host_csr_req_bits_addr;
    end
    if(T40) begin
      host_csr_bits_rw <= io_host_csr_req_bits_rw;
    end
    if(reset) begin
      reg_mstatus_ie <= 1'h0;
    end else if(T76) begin
      reg_mstatus_ie <= T243;
    end else if(T58) begin
      reg_mstatus_ie <= T242;
    end else if(insn_ret) begin
      reg_mstatus_ie <= reg_mstatus_ie1;
    end else if(T25) begin
      reg_mstatus_ie <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_ie1 <= 1'h0;
    end else if(T76) begin
      reg_mstatus_ie1 <= T241;
    end else if(T58) begin
      reg_mstatus_ie1 <= T240;
    end else if(insn_ret) begin
      reg_mstatus_ie1 <= reg_mstatus_ie2;
    end else if(T25) begin
      reg_mstatus_ie1 <= reg_mstatus_ie;
    end
    if(reset) begin
      reg_mstatus_ie2 <= 1'h0;
    end else if(T58) begin
      reg_mstatus_ie2 <= T239;
    end else if(insn_ret) begin
      reg_mstatus_ie2 <= 1'h1;
    end else if(T25) begin
      reg_mstatus_ie2 <= reg_mstatus_ie1;
    end
    if(reset) begin
      reg_mip_ssip <= 1'h0;
    end else if(T252) begin
      reg_mip_ssip <= T251;
    end else if(T250) begin
      reg_mip_ssip <= T249;
    end
    if(reset) begin
      reg_mie_ssip <= 1'h0;
    end else if(T258) begin
      reg_mie_ssip <= T257;
    end else if(T256) begin
      reg_mie_ssip <= T255;
    end
    if(reset) begin
      reg_mip_msip <= 1'h0;
    end else if(T268) begin
      reg_mip_msip <= 1'h1;
    end else if(T250) begin
      reg_mip_msip <= T267;
    end
    if(reset) begin
      reg_mie_msip <= 1'h0;
    end else if(T256) begin
      reg_mie_msip <= T270;
    end
    if(reset) begin
      reg_mip_stip <= 1'h0;
    end else if(T250) begin
      reg_mip_stip <= T278;
    end
    if(reset) begin
      reg_mie_stip <= 1'h0;
    end else if(T258) begin
      reg_mie_stip <= T282;
    end else if(T256) begin
      reg_mie_stip <= T281;
    end
    if(reset) begin
      reg_mip_mtip <= 1'h0;
    end else if(T295) begin
      reg_mip_mtip <= 1'h0;
    end else if(T291) begin
      reg_mip_mtip <= 1'h1;
    end
    if(T293) begin
      read_time <= wdata;
    end
    if(T295) begin
      reg_mtimecmp <= wdata;
    end
    if(reset) begin
      reg_mie_mtip <= 1'h0;
    end else if(T256) begin
      reg_mie_mtip <= T297;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T305) begin
      reg_fromhost <= wdata;
    end
    reg_frm <= T894;
    if(reset) begin
      R317 <= 6'h0;
    end else begin
      R317 <= T318;
    end
    if(reset) begin
      R320 <= 58'h0;
    end else if(T323) begin
      R320 <= T322;
    end
    reg_sepc <= T900;
    reg_mepc <= T902;
    reg_stvec <= T904;
    if(T363) begin
      reg_sptbr <= T361;
    end
    if(reset) begin
      reg_mstatus_ie3 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_prv3 <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_fs <= 2'h0;
    end else if(T76) begin
      reg_mstatus_fs <= T372;
    end else if(T58) begin
      reg_mstatus_fs <= T371;
    end
    if(reset) begin
      reg_mstatus_xs <= 2'h0;
    end
    if(reset) begin
      reg_mstatus_mprv <= 1'h0;
    end else if(T76) begin
      reg_mstatus_mprv <= T381;
    end else if(T58) begin
      reg_mstatus_mprv <= T380;
    end else if(T25) begin
      reg_mstatus_mprv <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_vm <= 5'h0;
    end else if(T388) begin
      reg_mstatus_vm <= 5'h9;
    end else if(T385) begin
      reg_mstatus_vm <= 5'h0;
    end
    if(reset) begin
      reg_mstatus_zero1 <= 9'h0;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_zero2 <= 31'h0;
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else if(some_interrupt_pending) begin
      reg_wfi <= 1'h0;
    end else if(insn_wfi) begin
      reg_wfi <= 1'h1;
    end
    if(insn_redirect_trap) begin
      reg_sbadaddr <= reg_mbadaddr;
    end
    if(T457) begin
      reg_mbadaddr <= T456;
    end else if(T448) begin
      reg_mbadaddr <= T440;
    end else if(T25) begin
      reg_mbadaddr <= io_pc;
    end
    if(insn_redirect_trap) begin
      reg_scause <= reg_mcause;
    end
    if(T473) begin
      reg_mcause <= T472;
    end else if(T471) begin
      reg_mcause <= T915;
    end else if(T469) begin
      reg_mcause <= 64'h3;
    end else if(T468) begin
      reg_mcause <= 64'h2;
    end else if(T25) begin
      reg_mcause <= io_cause;
    end
    if(T477) begin
      reg_sscratch <= wdata;
    end
    if(reset) begin
      R566 <= 6'h0;
    end else if(T570) begin
      R566 <= T568;
    end
    if(reset) begin
      R571 <= 58'h0;
    end else if(T574) begin
      R571 <= T573;
    end
    if(reset) begin
      R579 <= 6'h0;
    end else if(T583) begin
      R579 <= T581;
    end
    if(reset) begin
      R584 <= 58'h0;
    end else if(T587) begin
      R584 <= T586;
    end
    if(reset) begin
      R592 <= 6'h0;
    end else if(T596) begin
      R592 <= T594;
    end
    if(reset) begin
      R597 <= 58'h0;
    end else if(T600) begin
      R597 <= T599;
    end
    if(reset) begin
      R605 <= 6'h0;
    end else if(T609) begin
      R605 <= T607;
    end
    if(reset) begin
      R610 <= 58'h0;
    end else if(T613) begin
      R610 <= T612;
    end
    if(reset) begin
      R618 <= 6'h0;
    end else if(T622) begin
      R618 <= T620;
    end
    if(reset) begin
      R623 <= 58'h0;
    end else if(T626) begin
      R623 <= T625;
    end
    if(reset) begin
      R631 <= 6'h0;
    end else if(T635) begin
      R631 <= T633;
    end
    if(reset) begin
      R636 <= 58'h0;
    end else if(T639) begin
      R636 <= T638;
    end
    if(reset) begin
      R644 <= 6'h0;
    end else if(T648) begin
      R644 <= T646;
    end
    if(reset) begin
      R649 <= 58'h0;
    end else if(T652) begin
      R649 <= T651;
    end
    if(reset) begin
      R657 <= 6'h0;
    end else if(T661) begin
      R657 <= T659;
    end
    if(reset) begin
      R662 <= 58'h0;
    end else if(T665) begin
      R662 <= T664;
    end
    if(reset) begin
      R670 <= 6'h0;
    end else if(T674) begin
      R670 <= T672;
    end
    if(reset) begin
      R675 <= 58'h0;
    end else if(T678) begin
      R675 <= T677;
    end
    if(reset) begin
      R683 <= 6'h0;
    end else if(T687) begin
      R683 <= T685;
    end
    if(reset) begin
      R688 <= 58'h0;
    end else if(T691) begin
      R688 <= T690;
    end
    if(reset) begin
      R696 <= 6'h0;
    end else if(T700) begin
      R696 <= T698;
    end
    if(reset) begin
      R701 <= 58'h0;
    end else if(T704) begin
      R701 <= T703;
    end
    if(reset) begin
      R709 <= 6'h0;
    end else if(T713) begin
      R709 <= T711;
    end
    if(reset) begin
      R714 <= 58'h0;
    end else if(T717) begin
      R714 <= T716;
    end
    if(reset) begin
      R722 <= 6'h0;
    end else if(T726) begin
      R722 <= T724;
    end
    if(reset) begin
      R727 <= 58'h0;
    end else if(T730) begin
      R727 <= T729;
    end
    if(reset) begin
      R735 <= 6'h0;
    end else if(T739) begin
      R735 <= T737;
    end
    if(reset) begin
      R740 <= 58'h0;
    end else if(T743) begin
      R740 <= T742;
    end
    if(reset) begin
      R748 <= 6'h0;
    end else if(T752) begin
      R748 <= T750;
    end
    if(reset) begin
      R753 <= 58'h0;
    end else if(T756) begin
      R753 <= T755;
    end
    if(reset) begin
      R761 <= 6'h0;
    end else if(T765) begin
      R761 <= T763;
    end
    if(reset) begin
      R766 <= 58'h0;
    end else if(T769) begin
      R766 <= T768;
    end
    if(reset) begin
      R774 <= 6'h0;
    end else if(T781) begin
      R774 <= T780;
    end else if(T779) begin
      R774 <= T777;
    end
    if(reset) begin
      R782 <= 58'h0;
    end else if(T781) begin
      R782 <= T788;
    end else if(T786) begin
      R782 <= T785;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T800) begin
      reg_tohost <= wdata;
    end else if(T797) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T808) begin
      reg_stats <= T807;
    end
    if(T828) begin
      reg_mscratch <= wdata;
    end
    if(reset) begin
      reg_mie_usip <= 1'h0;
    end
    if(reset) begin
      reg_mie_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mie_utip <= 1'h0;
    end
    if(reset) begin
      reg_mie_htip <= 1'h0;
    end
    if(reset) begin
      reg_mip_usip <= 1'h0;
    end
    if(reset) begin
      reg_mip_hsip <= 1'h0;
    end
    if(reset) begin
      reg_mip_utip <= 1'h0;
    end
    if(reset) begin
      reg_mip_htip <= 1'h0;
    end
    if(T877) begin
      host_csr_rep_valid <= 1'h0;
    end else if(host_csr_req_fire) begin
      host_csr_rep_valid <= 1'h1;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] out;
  wire[63:0] T4;
  wire[63:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T136;
  wire cmp;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[63:0] T23;
  wire T24;
  wire[63:0] T25;
  wire T26;
  wire[63:0] T27;
  wire T28;
  wire[63:0] shout_l;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[62:0] T31;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[63:0] T34;
  wire[61:0] T35;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[59:0] T39;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[55:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[47:0] T47;
  wire[63:0] T48;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[31:0] T51;
  wire[63:0] T52;
  wire[63:0] T137;
  wire[31:0] T53;
  wire[63:0] T54;
  wire[63:0] T138;
  wire[47:0] T55;
  wire[63:0] T56;
  wire[63:0] T139;
  wire[55:0] T57;
  wire[63:0] T58;
  wire[63:0] T140;
  wire[59:0] T59;
  wire[63:0] T60;
  wire[63:0] T141;
  wire[61:0] T61;
  wire[63:0] T62;
  wire[63:0] T142;
  wire[62:0] T63;
  wire T64;
  wire[63:0] shout_r;
  wire[64:0] T65;
  wire[5:0] shamt;
  wire[4:0] T66;
  wire[5:0] full_shamt;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[64:0] T71;
  wire[64:0] T72;
  wire[63:0] shin;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  wire[62:0] T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[63:0] T79;
  wire[61:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[59:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] T87;
  wire[55:0] T88;
  wire[63:0] T89;
  wire[63:0] T90;
  wire[63:0] T91;
  wire[47:0] T92;
  wire[63:0] T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[31:0] T96;
  wire[63:0] T97;
  wire[63:0] T143;
  wire[31:0] T98;
  wire[63:0] T99;
  wire[63:0] T144;
  wire[47:0] T100;
  wire[63:0] T101;
  wire[63:0] T145;
  wire[55:0] T102;
  wire[63:0] T103;
  wire[63:0] T146;
  wire[59:0] T104;
  wire[63:0] T105;
  wire[63:0] T147;
  wire[61:0] T106;
  wire[63:0] T107;
  wire[63:0] T148;
  wire[62:0] T108;
  wire[63:0] shin_r;
  wire[31:0] T109;
  wire[31:0] T110;
  wire[31:0] T111;
  wire[31:0] T149;
  wire T112;
  wire T113;
  wire T114;
  wire[31:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire[63:0] T130;
  wire[31:0] T131;
  wire[31:0] T132;
  wire[31:0] T150;
  wire T133;
  wire T134;
  wire T135;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T134 ? T130 : out;
  assign out = T127 ? sum : T4;
  assign T4 = T124 ? shout_r : T5;
  assign T5 = T64 ? shout_l : T6;
  assign T6 = T28 ? T27 : T7;
  assign T7 = T26 ? T25 : T8;
  assign T8 = T24 ? T23 : T136;
  assign T136 = {63'h0, cmp};
  assign cmp = T22 ^ T9;
  assign T9 = T20 ? T19 : T10;
  assign T10 = T16 ? T15 : T11;
  assign T11 = T14 ? T13 : T12;
  assign T12 = io_in1[6'h3f:6'h3f];
  assign T13 = io_in2[6'h3f:6'h3f];
  assign T14 = io_fn[1'h1:1'h1];
  assign T15 = sum[6'h3f:6'h3f];
  assign T16 = T18 == T17;
  assign T17 = io_in2[6'h3f:6'h3f];
  assign T18 = io_in1[6'h3f:6'h3f];
  assign T19 = sum == 64'h0;
  assign T20 = T21 ^ 1'h1;
  assign T21 = io_fn[2'h2:2'h2];
  assign T22 = io_fn[1'h0:1'h0];
  assign T23 = io_in1 ^ io_in2;
  assign T24 = io_fn == 4'h4;
  assign T25 = io_in1 | io_in2;
  assign T26 = io_fn == 4'h6;
  assign T27 = io_in1 & io_in2;
  assign T28 = io_fn == 4'h7;
  assign shout_l = T62 | T29;
  assign T29 = T30 & 64'haaaaaaaaaaaaaaaa;
  assign T30 = T31 << 1'h1;
  assign T31 = T32[6'h3e:1'h0];
  assign T32 = T60 | T33;
  assign T33 = T34 & 64'hcccccccccccccccc;
  assign T34 = T35 << 2'h2;
  assign T35 = T36[6'h3d:1'h0];
  assign T36 = T58 | T37;
  assign T37 = T38 & 64'hf0f0f0f0f0f0f0f0;
  assign T38 = T39 << 3'h4;
  assign T39 = T40[6'h3b:1'h0];
  assign T40 = T56 | T41;
  assign T41 = T42 & 64'hff00ff00ff00ff00;
  assign T42 = T43 << 4'h8;
  assign T43 = T44[6'h37:1'h0];
  assign T44 = T54 | T45;
  assign T45 = T46 & 64'hffff0000ffff0000;
  assign T46 = T47 << 5'h10;
  assign T47 = T48[6'h2f:1'h0];
  assign T48 = T52 | T49;
  assign T49 = T50 & 64'hffffffff00000000;
  assign T50 = T51 << 6'h20;
  assign T51 = shout_r[5'h1f:1'h0];
  assign T52 = T137 & 64'hffffffff;
  assign T137 = {32'h0, T53};
  assign T53 = shout_r >> 6'h20;
  assign T54 = T138 & 64'hffff0000ffff;
  assign T138 = {16'h0, T55};
  assign T55 = T48 >> 5'h10;
  assign T56 = T139 & 64'hff00ff00ff00ff;
  assign T139 = {8'h0, T57};
  assign T57 = T44 >> 4'h8;
  assign T58 = T140 & 64'hf0f0f0f0f0f0f0f;
  assign T140 = {4'h0, T59};
  assign T59 = T40 >> 3'h4;
  assign T60 = T141 & 64'h3333333333333333;
  assign T141 = {2'h0, T61};
  assign T61 = T36 >> 2'h2;
  assign T62 = T142 & 64'h5555555555555555;
  assign T142 = {1'h0, T63};
  assign T63 = T32 >> 1'h1;
  assign T64 = io_fn == 4'h1;
  assign shout_r = T65[6'h3f:1'h0];
  assign T65 = $signed(T71) >>> shamt;
  assign shamt = {T67, T66};
  assign T66 = full_shamt[3'h4:1'h0];
  assign full_shamt = io_in2[3'h5:1'h0];
  assign T67 = T70 & T68;
  assign T68 = 1'h1 == T69;
  assign T69 = io_dw & 1'h1;
  assign T70 = full_shamt[3'h5:3'h5];
  assign T71 = T72;
  assign T72 = {T121, shin};
  assign shin = T118 ? shin_r : T73;
  assign T73 = T107 | T74;
  assign T74 = T75 & 64'haaaaaaaaaaaaaaaa;
  assign T75 = T76 << 1'h1;
  assign T76 = T77[6'h3e:1'h0];
  assign T77 = T105 | T78;
  assign T78 = T79 & 64'hcccccccccccccccc;
  assign T79 = T80 << 2'h2;
  assign T80 = T81[6'h3d:1'h0];
  assign T81 = T103 | T82;
  assign T82 = T83 & 64'hf0f0f0f0f0f0f0f0;
  assign T83 = T84 << 3'h4;
  assign T84 = T85[6'h3b:1'h0];
  assign T85 = T101 | T86;
  assign T86 = T87 & 64'hff00ff00ff00ff00;
  assign T87 = T88 << 4'h8;
  assign T88 = T89[6'h37:1'h0];
  assign T89 = T99 | T90;
  assign T90 = T91 & 64'hffff0000ffff0000;
  assign T91 = T92 << 5'h10;
  assign T92 = T93[6'h2f:1'h0];
  assign T93 = T97 | T94;
  assign T94 = T95 & 64'hffffffff00000000;
  assign T95 = T96 << 6'h20;
  assign T96 = shin_r[5'h1f:1'h0];
  assign T97 = T143 & 64'hffffffff;
  assign T143 = {32'h0, T98};
  assign T98 = shin_r >> 6'h20;
  assign T99 = T144 & 64'hffff0000ffff;
  assign T144 = {16'h0, T100};
  assign T100 = T93 >> 5'h10;
  assign T101 = T145 & 64'hff00ff00ff00ff;
  assign T145 = {8'h0, T102};
  assign T102 = T89 >> 4'h8;
  assign T103 = T146 & 64'hf0f0f0f0f0f0f0f;
  assign T146 = {4'h0, T104};
  assign T104 = T85 >> 3'h4;
  assign T105 = T147 & 64'h3333333333333333;
  assign T147 = {2'h0, T106};
  assign T106 = T81 >> 2'h2;
  assign T107 = T148 & 64'h5555555555555555;
  assign T148 = {1'h0, T108};
  assign T108 = T77 >> 1'h1;
  assign shin_r = {T110, T109};
  assign T109 = io_in1[5'h1f:1'h0];
  assign T110 = T116 ? T115 : T111;
  assign T111 = 32'h0 - T149;
  assign T149 = {31'h0, T112};
  assign T112 = T114 & T113;
  assign T113 = io_in1[5'h1f:5'h1f];
  assign T114 = io_fn[2'h3:2'h3];
  assign T115 = io_in1[6'h3f:6'h20];
  assign T116 = 1'h1 == T117;
  assign T117 = io_dw & 1'h1;
  assign T118 = T120 | T119;
  assign T119 = io_fn == 4'hb;
  assign T120 = io_fn == 4'h5;
  assign T121 = T123 & T122;
  assign T122 = shin[6'h3f:6'h3f];
  assign T123 = io_fn[2'h3:2'h3];
  assign T124 = T126 | T125;
  assign T125 = io_fn == 4'hb;
  assign T126 = io_fn == 4'h5;
  assign T127 = T129 | T128;
  assign T128 = io_fn == 4'ha;
  assign T129 = io_fn == 4'h0;
  assign T130 = {T132, T131};
  assign T131 = out[5'h1f:1'h0];
  assign T132 = 32'h0 - T150;
  assign T150 = {31'h0, T133};
  assign T133 = out[5'h1f:5'h1f];
  assign T134 = 1'h0 == T135;
  assign T135 = io_dw & 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T148;
  wire[63:0] negated_remainder;
  wire[63:0] T95;
  wire T10;
  wire T11;
  reg  isMul;
  wire T12;
  wire cmdMul;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire T19;
  reg [2:0] state;
  wire[2:0] T149;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  reg  neg_out;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  reg  isHi;
  wire T33;
  wire cmdHi;
  wire T34;
  wire T35;
  wire T36;
  wire[3:0] T37;
  wire T38;
  wire[3:0] T39;
  wire T40;
  wire T41;
  wire less;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T42;
  wire[64:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[64:0] T47;
  wire[63:0] rhs_in;
  wire[31:0] T48;
  wire[31:0] T49;
  wire[31:0] T50;
  wire[31:0] T150;
  wire[31:0] T51;
  wire T52;
  wire T53;
  wire rhs_sign;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire rhsSigned;
  wire T59;
  wire T60;
  wire[3:0] T61;
  wire[64:0] T62;
  wire T63;
  reg [6:0] count;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[6:0] T68;
  wire T69;
  wire T70;
  wire T71;
  wire lhs_sign;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire lhsSigned;
  wire T77;
  wire T78;
  wire[3:0] T79;
  wire T80;
  wire T81;
  wire[2:0] T82;
  wire T83;
  wire T84;
  wire[2:0] T85;
  wire[2:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire[129:0] T151;
  wire T96;
  wire[129:0] T152;
  wire[63:0] T97;
  wire T98;
  wire[129:0] T99;
  wire[64:0] T100;
  wire[63:0] T101;
  wire[128:0] T102;
  wire[63:0] T103;
  wire[128:0] T104;
  wire[128:0] T105;
  wire[62:0] T106;
  wire[63:0] T107;
  wire[128:0] T108;
  wire[63:0] T109;
  wire[64:0] T110;
  wire[65:0] T111;
  wire[65:0] T153;
  wire[64:0] T112;
  wire[64:0] T113;
  wire T154;
  wire[65:0] T114;
  wire[1:0] T115;
  wire[1:0] T116;
  wire T117;
  wire[64:0] T118;
  wire[64:0] T119;
  wire[64:0] T120;
  wire T121;
  wire T122;
  wire[129:0] T155;
  wire[128:0] T123;
  wire[64:0] T124;
  wire T125;
  wire[63:0] T126;
  wire[63:0] T127;
  wire[63:0] T128;
  wire[63:0] T129;
  wire T130;
  wire T131;
  wire T132;
  wire[129:0] T156;
  wire[63:0] lhs_in;
  wire[31:0] T133;
  wire[31:0] T134;
  wire[31:0] T135;
  wire[31:0] T157;
  wire[31:0] T136;
  wire T137;
  wire T138;
  wire[63:0] T139;
  wire[31:0] T140;
  wire[31:0] T141;
  wire[31:0] T158;
  wire T142;
  wire T143;
  wire T144;
  reg  req_dw;
  wire T145;
  wire T146;
  wire T147;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T143 ? T139 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T156 : T5;
  assign T5 = T130 ? T155 : T6;
  assign T6 = T121 ? T99 : T7;
  assign T7 = T98 ? T152 : T8;
  assign T8 = T96 ? T151 : T9;
  assign T9 = T10 ? T148 : remainder;
  assign T148 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T95;
  assign T95 = remainder[6'h3f:1'h0];
  assign T10 = T19 & T11;
  assign T11 = T18 | isMul;
  assign T12 = T1 ? cmdMul : isMul;
  assign cmdMul = T13;
  assign T13 = T16 | T14;
  assign T14 = T15 == 4'h8;
  assign T15 = io_req_bits_fn & 4'h8;
  assign T16 = T17 == 4'h0;
  assign T17 = io_req_bits_fn & 4'h4;
  assign T18 = remainder[6'h3f:6'h3f];
  assign T19 = state == 3'h1;
  assign T149 = reset ? 3'h0 : T20;
  assign T20 = T1 ? T91 : T21;
  assign T21 = T89 ? 3'h0 : T22;
  assign T22 = T87 ? T85 : T23;
  assign T23 = T83 ? T82 : T24;
  assign T24 = T98 ? T27 : T25;
  assign T25 = T96 ? 3'h5 : T26;
  assign T26 = T19 ? 3'h2 : state;
  assign T27 = neg_out ? 3'h4 : 3'h5;
  assign T28 = T1 ? T69 : T29;
  assign T29 = T30 ? 1'h0 : neg_out;
  assign T30 = T130 & T31;
  assign T31 = T40 & T32;
  assign T32 = isHi ^ 1'h1;
  assign T33 = T1 ? cmdHi : isHi;
  assign cmdHi = T34;
  assign T34 = T35 | T14;
  assign T35 = T38 | T36;
  assign T36 = T37 == 4'h2;
  assign T37 = io_req_bits_fn & 4'h2;
  assign T38 = T39 == 4'h1;
  assign T39 = io_req_bits_fn & 4'h5;
  assign T40 = T63 & T41;
  assign T41 = less ^ 1'h1;
  assign less = subtractor[7'h40:7'h40];
  assign subtractor = T62 - divisor;
  assign T42 = T1 ? T47 : T43;
  assign T43 = T44 ? subtractor : divisor;
  assign T44 = T19 & T45;
  assign T45 = T46 | isMul;
  assign T46 = divisor[6'h3f:6'h3f];
  assign T47 = {rhs_sign, rhs_in};
  assign rhs_in = {T49, T48};
  assign T48 = io_req_bits_in2[5'h1f:1'h0];
  assign T49 = T52 ? T51 : T50;
  assign T50 = 32'h0 - T150;
  assign T150 = {31'h0, rhs_sign};
  assign T51 = io_req_bits_in2[6'h3f:6'h20];
  assign T52 = 1'h1 == T53;
  assign T53 = io_req_bits_dw & 1'h1;
  assign rhs_sign = rhsSigned & T54;
  assign T54 = T57 ? T56 : T55;
  assign T55 = io_req_bits_in2[5'h1f:5'h1f];
  assign T56 = io_req_bits_in2[6'h3f:6'h3f];
  assign T57 = 1'h1 == T58;
  assign T58 = io_req_bits_dw & 1'h1;
  assign rhsSigned = T59;
  assign T59 = T60 | T16;
  assign T60 = T61 == 4'h0;
  assign T61 = io_req_bits_fn & 4'h9;
  assign T62 = remainder[8'h80:7'h40];
  assign T63 = count == 7'h0;
  assign T64 = T1 ? 7'h0 : T65;
  assign T65 = T130 ? T68 : T66;
  assign T66 = T121 ? T67 : count;
  assign T67 = count + 7'h1;
  assign T68 = count + 7'h1;
  assign T69 = T81 & T70;
  assign T70 = cmdHi ? lhs_sign : T71;
  assign T71 = lhs_sign != rhs_sign;
  assign lhs_sign = lhsSigned & T72;
  assign T72 = T75 ? T74 : T73;
  assign T73 = io_req_bits_in1[5'h1f:5'h1f];
  assign T74 = io_req_bits_in1[6'h3f:6'h3f];
  assign T75 = 1'h1 == T76;
  assign T76 = io_req_bits_dw & 1'h1;
  assign lhsSigned = T77;
  assign T77 = T80 | T78;
  assign T78 = T79 == 4'h0;
  assign T79 = io_req_bits_fn & 4'h3;
  assign T80 = T60 | T16;
  assign T81 = cmdMul ^ 1'h1;
  assign T82 = isHi ? 3'h3 : 3'h5;
  assign T83 = T121 & T84;
  assign T84 = count == 7'h3f;
  assign T85 = isHi ? 3'h3 : T86;
  assign T86 = neg_out ? 3'h4 : 3'h5;
  assign T87 = T130 & T88;
  assign T88 = count == 7'h40;
  assign T89 = T90 | io_kill;
  assign T90 = io_resp_ready & io_resp_valid;
  assign T91 = T92 ? 3'h1 : 3'h2;
  assign T92 = lhs_sign | T93;
  assign T93 = rhs_sign & T94;
  assign T94 = cmdMul ^ 1'h1;
  assign T151 = {66'h0, negated_remainder};
  assign T96 = state == 3'h4;
  assign T152 = {66'h0, T97};
  assign T97 = remainder[8'h80:7'h41];
  assign T98 = state == 3'h3;
  assign T99 = {T120, T100};
  assign T100 = {1'h0, T101};
  assign T101 = T102[6'h3f:1'h0];
  assign T102 = {T119, T103};
  assign T103 = T104[6'h3f:1'h0];
  assign T104 = T105;
  assign T105 = {T111, T106};
  assign T106 = T107[6'h3f:1'h1];
  assign T107 = T108[6'h3f:1'h0];
  assign T108 = {T110, T109};
  assign T109 = remainder[6'h3f:1'h0];
  assign T110 = remainder[8'h81:7'h41];
  assign T111 = T114 + T153;
  assign T153 = {T154, T112};
  assign T112 = T113;
  assign T113 = T108[8'h80:7'h40];
  assign T154 = T112[7'h40:7'h40];
  assign T114 = $signed(T118) * $signed(T115);
  assign T115 = T116;
  assign T116 = {1'h0, T117};
  assign T117 = T107[1'h0:1'h0];
  assign T118 = divisor;
  assign T119 = T104[8'h80:7'h40];
  assign T120 = T102 >> 7'h40;
  assign T121 = T122 & isMul;
  assign T122 = state == 3'h2;
  assign T155 = {1'h0, T123};
  assign T123 = {T127, T124};
  assign T124 = {T126, T125};
  assign T125 = less ^ 1'h1;
  assign T126 = remainder[6'h3f:1'h0];
  assign T127 = less ? T129 : T128;
  assign T128 = subtractor[6'h3f:1'h0];
  assign T129 = remainder[7'h7f:7'h40];
  assign T130 = T132 & T131;
  assign T131 = isMul ^ 1'h1;
  assign T132 = state == 3'h2;
  assign T156 = {66'h0, lhs_in};
  assign lhs_in = {T134, T133};
  assign T133 = io_req_bits_in1[5'h1f:1'h0];
  assign T134 = T137 ? T136 : T135;
  assign T135 = 32'h0 - T157;
  assign T157 = {31'h0, lhs_sign};
  assign T136 = io_req_bits_in1[6'h3f:6'h20];
  assign T137 = 1'h1 == T138;
  assign T138 = io_req_bits_dw & 1'h1;
  assign T139 = {T141, T140};
  assign T140 = remainder[5'h1f:1'h0];
  assign T141 = 32'h0 - T158;
  assign T158 = {31'h0, T142};
  assign T142 = remainder[5'h1f:5'h1f];
  assign T143 = 1'h0 == T144;
  assign T144 = req_dw & 1'h1;
  assign T145 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T146;
  assign T146 = state == 3'h5;
  assign io_req_ready = T147;
  assign T147 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T156;
    end else if(T130) begin
      remainder <= T155;
    end else if(T121) begin
      remainder <= T99;
    end else if(T98) begin
      remainder <= T152;
    end else if(T96) begin
      remainder <= T151;
    end else if(T10) begin
      remainder <= T148;
    end
    if(T1) begin
      isMul <= cmdMul;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T91;
    end else if(T89) begin
      state <= 3'h0;
    end else if(T87) begin
      state <= T85;
    end else if(T83) begin
      state <= T82;
    end else if(T98) begin
      state <= T27;
    end else if(T96) begin
      state <= 3'h5;
    end else if(T19) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T69;
    end else if(T30) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= cmdHi;
    end
    if(T1) begin
      divisor <= T47;
    end else if(T44) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T130) begin
      count <= T68;
    end else if(T121) begin
      count <= T67;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module Rocket(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    output io_imem_req_valid,
    output[39:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [39:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data_0,
    input  io_imem_resp_bits_mask,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input  io_imem_btb_resp_bits_mask,
    input  io_imem_btb_resp_bits_bridx,
    input [38:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_history,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_btb_update_bits_pc,
    output[38:0] io_imem_btb_update_bits_target,
    //output io_imem_btb_update_bits_taken
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output[38:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_bht_update_bits_prediction_bits_target,
    output[2:0] io_imem_bht_update_bits_prediction_bits_entry,
    output[3:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output[38:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output[38:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output[38:0] io_imem_ras_update_bits_prediction_bits_target,
    output[2:0] io_imem_ras_update_bits_prediction_bits_entry,
    output[3:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output[1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    output io_imem_invalidate,
    input [39:0] io_imem_npc,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output[39:0] io_dmem_req_bits_addr,
    output[8:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_kill,
    output io_dmem_req_bits_phys,
    output[63:0] io_dmem_req_bits_data,
    input  io_dmem_resp_valid,
    input [39:0] io_dmem_resp_bits_addr,
    input [8:0] io_dmem_resp_bits_tag,
    input [4:0] io_dmem_resp_bits_cmd,
    input [2:0] io_dmem_resp_bits_typ,
    input [63:0] io_dmem_resp_bits_data,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_word_bypass,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [8:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    output io_dmem_invalidate_lr,
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_status_sd,
    output[30:0] io_ptw_status_zero2,
    output io_ptw_status_sd_rv32,
    output[8:0] io_ptw_status_zero1,
    output[4:0] io_ptw_status_vm,
    output io_ptw_status_mprv,
    output[1:0] io_ptw_status_xs,
    output[1:0] io_ptw_status_fs,
    output[1:0] io_ptw_status_prv3,
    output io_ptw_status_ie3,
    output[1:0] io_ptw_status_prv2,
    output io_ptw_status_ie2,
    output[1:0] io_ptw_status_prv1,
    output io_ptw_status_ie1,
    output[1:0] io_ptw_status_prv,
    output io_ptw_status_ie,
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    output io_fpu_valid,
    //input  io_fpu_fcsr_rdy
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    //input [4:0] io_fpu_dec_cmd
    //input  io_fpu_dec_ldst
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    //input  io_fpu_dec_swap12
    //input  io_fpu_dec_swap23
    //input  io_fpu_dec_single
    //input  io_fpu_dec_fromint
    //input  io_fpu_dec_toint
    //input  io_fpu_dec_fastpipe
    //input  io_fpu_dec_fma
    //input  io_fpu_dec_div
    //input  io_fpu_dec_sqrt
    //input  io_fpu_dec_round
    //input  io_fpu_dec_wflags
    //input  io_fpu_sboard_set
    //input  io_fpu_sboard_clr
    //input [4:0] io_fpu_sboard_clra
    //input  io_fpu_cp_req_ready
    //output io_fpu_cp_req_valid
    //output[4:0] io_fpu_cp_req_bits_cmd
    //output io_fpu_cp_req_bits_ldst
    //output io_fpu_cp_req_bits_wen
    //output io_fpu_cp_req_bits_ren1
    //output io_fpu_cp_req_bits_ren2
    //output io_fpu_cp_req_bits_ren3
    //output io_fpu_cp_req_bits_swap12
    //output io_fpu_cp_req_bits_swap23
    //output io_fpu_cp_req_bits_single
    //output io_fpu_cp_req_bits_fromint
    //output io_fpu_cp_req_bits_toint
    //output io_fpu_cp_req_bits_fastpipe
    //output io_fpu_cp_req_bits_fma
    //output io_fpu_cp_req_bits_div
    //output io_fpu_cp_req_bits_sqrt
    //output io_fpu_cp_req_bits_round
    //output io_fpu_cp_req_bits_wflags
    //output[2:0] io_fpu_cp_req_bits_rm
    //output[1:0] io_fpu_cp_req_bits_typ
    //output[64:0] io_fpu_cp_req_bits_in1
    //output[64:0] io_fpu_cp_req_bits_in2
    //output[64:0] io_fpu_cp_req_bits_in3
    //output io_fpu_cp_resp_ready
    //input  io_fpu_cp_resp_valid
    //input [64:0] io_fpu_cp_resp_bits_data
    //input [4:0] io_fpu_cp_resp_bits_exc
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [8:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_kill,
    input  io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    //output io_rocc_mem_resp_valid
    //output[39:0] io_rocc_mem_resp_bits_addr
    //output[8:0] io_rocc_mem_resp_bits_tag
    //output[4:0] io_rocc_mem_resp_bits_cmd
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output[63:0] io_rocc_mem_resp_bits_data
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data_word_bypass
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[8:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_invalidate_lr,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_autl_acquire_ready
    input  io_rocc_autl_acquire_valid,
    input [25:0] io_rocc_autl_acquire_bits_addr_block,
    input [1:0] io_rocc_autl_acquire_bits_client_xact_id,
    input [1:0] io_rocc_autl_acquire_bits_addr_beat,
    input  io_rocc_autl_acquire_bits_is_builtin_type,
    input [2:0] io_rocc_autl_acquire_bits_a_type,
    input [16:0] io_rocc_autl_acquire_bits_union,
    input [127:0] io_rocc_autl_acquire_bits_data,
    input  io_rocc_autl_grant_ready,
    //output io_rocc_autl_grant_valid
    //output[1:0] io_rocc_autl_grant_bits_addr_beat
    //output[1:0] io_rocc_autl_grant_bits_client_xact_id
    //output[2:0] io_rocc_autl_grant_bits_manager_xact_id
    //output io_rocc_autl_grant_bits_is_builtin_type
    //output[3:0] io_rocc_autl_grant_bits_g_type
    //output[127:0] io_rocc_autl_grant_bits_data
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [26:0] io_rocc_iptw_req_bits_addr,
    input [1:0] io_rocc_iptw_req_bits_prv,
    input  io_rocc_iptw_req_bits_store,
    input  io_rocc_iptw_req_bits_fetch,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[19:0] io_rocc_iptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_iptw_resp_bits_pte_reserved_for_software
    //output io_rocc_iptw_resp_bits_pte_d
    //output io_rocc_iptw_resp_bits_pte_r
    //output[3:0] io_rocc_iptw_resp_bits_pte_typ
    //output io_rocc_iptw_resp_bits_pte_v
    //output io_rocc_iptw_status_sd
    //output[30:0] io_rocc_iptw_status_zero2
    //output io_rocc_iptw_status_sd_rv32
    //output[8:0] io_rocc_iptw_status_zero1
    //output[4:0] io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_mprv
    //output[1:0] io_rocc_iptw_status_xs
    //output[1:0] io_rocc_iptw_status_fs
    //output[1:0] io_rocc_iptw_status_prv3
    //output io_rocc_iptw_status_ie3
    //output[1:0] io_rocc_iptw_status_prv2
    //output io_rocc_iptw_status_ie2
    //output[1:0] io_rocc_iptw_status_prv1
    //output io_rocc_iptw_status_ie1
    //output[1:0] io_rocc_iptw_status_prv
    //output io_rocc_iptw_status_ie
    //output io_rocc_iptw_invalidate
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [26:0] io_rocc_dptw_req_bits_addr,
    input [1:0] io_rocc_dptw_req_bits_prv,
    input  io_rocc_dptw_req_bits_store,
    input  io_rocc_dptw_req_bits_fetch,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[19:0] io_rocc_dptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_dptw_resp_bits_pte_reserved_for_software
    //output io_rocc_dptw_resp_bits_pte_d
    //output io_rocc_dptw_resp_bits_pte_r
    //output[3:0] io_rocc_dptw_resp_bits_pte_typ
    //output io_rocc_dptw_resp_bits_pte_v
    //output io_rocc_dptw_status_sd
    //output[30:0] io_rocc_dptw_status_zero2
    //output io_rocc_dptw_status_sd_rv32
    //output[8:0] io_rocc_dptw_status_zero1
    //output[4:0] io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_mprv
    //output[1:0] io_rocc_dptw_status_xs
    //output[1:0] io_rocc_dptw_status_fs
    //output[1:0] io_rocc_dptw_status_prv3
    //output io_rocc_dptw_status_ie3
    //output[1:0] io_rocc_dptw_status_prv2
    //output io_rocc_dptw_status_ie2
    //output[1:0] io_rocc_dptw_status_prv1
    //output io_rocc_dptw_status_ie1
    //output[1:0] io_rocc_dptw_status_prv
    //output io_rocc_dptw_status_ie
    //output io_rocc_dptw_invalidate
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [26:0] io_rocc_pptw_req_bits_addr,
    input [1:0] io_rocc_pptw_req_bits_prv,
    input  io_rocc_pptw_req_bits_store,
    input  io_rocc_pptw_req_bits_fetch,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[19:0] io_rocc_pptw_resp_bits_pte_ppn
    //output[2:0] io_rocc_pptw_resp_bits_pte_reserved_for_software
    //output io_rocc_pptw_resp_bits_pte_d
    //output io_rocc_pptw_resp_bits_pte_r
    //output[3:0] io_rocc_pptw_resp_bits_pte_typ
    //output io_rocc_pptw_resp_bits_pte_v
    //output io_rocc_pptw_status_sd
    //output[30:0] io_rocc_pptw_status_zero2
    //output io_rocc_pptw_status_sd_rv32
    //output[8:0] io_rocc_pptw_status_zero1
    //output[4:0] io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_mprv
    //output[1:0] io_rocc_pptw_status_xs
    //output[1:0] io_rocc_pptw_status_fs
    //output[1:0] io_rocc_pptw_status_prv3
    //output io_rocc_pptw_status_ie3
    //output[1:0] io_rocc_pptw_status_prv2
    //output io_rocc_pptw_status_ie2
    //output[1:0] io_rocc_pptw_status_prv1
    //output io_rocc_pptw_status_ie1
    //output[1:0] io_rocc_pptw_status_prv
    //output io_rocc_pptw_status_ie
    //output io_rocc_pptw_invalidate
    //output io_rocc_fpu_req_ready
    input  io_rocc_fpu_req_valid,
    input [4:0] io_rocc_fpu_req_bits_cmd,
    input  io_rocc_fpu_req_bits_ldst,
    input  io_rocc_fpu_req_bits_wen,
    input  io_rocc_fpu_req_bits_ren1,
    input  io_rocc_fpu_req_bits_ren2,
    input  io_rocc_fpu_req_bits_ren3,
    input  io_rocc_fpu_req_bits_swap12,
    input  io_rocc_fpu_req_bits_swap23,
    input  io_rocc_fpu_req_bits_single,
    input  io_rocc_fpu_req_bits_fromint,
    input  io_rocc_fpu_req_bits_toint,
    input  io_rocc_fpu_req_bits_fastpipe,
    input  io_rocc_fpu_req_bits_fma,
    input  io_rocc_fpu_req_bits_div,
    input  io_rocc_fpu_req_bits_sqrt,
    input  io_rocc_fpu_req_bits_round,
    input  io_rocc_fpu_req_bits_wflags,
    input [2:0] io_rocc_fpu_req_bits_rm,
    input [1:0] io_rocc_fpu_req_bits_typ,
    input [64:0] io_rocc_fpu_req_bits_in1,
    input [64:0] io_rocc_fpu_req_bits_in2,
    input [64:0] io_rocc_fpu_req_bits_in3,
    input  io_rocc_fpu_resp_ready,
    //output io_rocc_fpu_resp_valid
    //output[64:0] io_rocc_fpu_resp_bits_data
    //output[4:0] io_rocc_fpu_resp_bits_exc
    output io_rocc_exception,
    //output io_rocc_dma_req_ready
    input  io_rocc_dma_req_valid,
    input [1:0] io_rocc_dma_req_bits_client_xact_id,
    input [1:0] io_rocc_dma_req_bits_cmd,
    input [31:0] io_rocc_dma_req_bits_source,
    input [31:0] io_rocc_dma_req_bits_dest,
    input [31:0] io_rocc_dma_req_bits_length,
    input  io_rocc_dma_resp_ready
    //output io_rocc_dma_resp_valid
    //output[1:0] io_rocc_dma_resp_bits_client_xact_id
    //output[1:0] io_rocc_dma_resp_bits_status
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  wire ctrl_killd;
  wire T7;
  wire T8;
  wire ctrl_stalld;
  wire T9;
  wire id_do_fence;
  wire T10;
  wire id_csr_en;
  wire[2:0] id_ctrl_csr;
  wire[2:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire[31:0] T16;
  wire T17;
  wire[31:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire id_ctrl_rocc;
  wire id_ctrl_mem;
  wire T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire[31:0] T38;
  reg  id_reg_fence;
  wire T917;
  wire T39;
  wire T40;
  wire id_fence_next;
  wire T41;
  wire id_amo_rl;
  wire id_ctrl_amo;
  wire T42;
  wire[31:0] T43;
  wire id_ctrl_fence;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire id_ctrl_fence_i;
  wire T47;
  wire[31:0] T48;
  wire T49;
  wire id_amo_aq;
  wire id_mem_busy;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire id_sboard_hazard;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[4:0] T59;
  wire[4:0] T60;
  wire[4:0] id_waddr;
  wire T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[4:0] ll_waddr;
  wire[4:0] T66;
  wire[4:0] dmem_resp_waddr;
  wire[8:0] T67;
  wire T68;
  wire dmem_resp_xpu;
  wire T69;
  wire T70;
  wire dmem_resp_replay;
  wire ll_wen;
  wire T71;
  wire T72;
  reg [31:0] R73;
  wire[31:0] T918;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[31:0] T76;
  wire[31:0] T77;
  wire[31:0] T78;
  wire[4:0] wb_waddr;
  wire T79;
  wire wb_wen;
  reg  wb_ctrl_wxd;
  wire T80;
  reg  mem_ctrl_wxd;
  wire T81;
  reg  ex_ctrl_wxd;
  wire T82;
  wire id_ctrl_wxd;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire[31:0] T91;
  wire T92;
  wire T93;
  wire[31:0] T94;
  wire T95;
  wire T96;
  wire[31:0] T97;
  wire T98;
  wire T99;
  wire[31:0] T100;
  wire T101;
  wire[31:0] T102;
  wire T103;
  wire wb_valid;
  wire T104;
  wire T105;
  wire T106;
  wire replay_wb;
  wire T107;
  wire T108;
  wire T109;
  reg  wb_ctrl_rocc;
  wire T110;
  reg  mem_ctrl_rocc;
  wire T111;
  reg  ex_ctrl_rocc;
  wire T112;
  wire replay_wb_common;
  reg  wb_reg_replay;
  wire T113;
  wire T114;
  wire take_pc_wb;
  wire T115;
  wire T116;
  wire wb_xcpt;
  reg  wb_reg_xcpt;
  wire T117;
  wire T118;
  wire mem_xcpt;
  wire T119;
  wire T120;
  reg  mem_ctrl_mem;
  wire T121;
  reg  ex_ctrl_mem;
  wire T122;
  reg  mem_reg_valid;
  wire T123;
  wire ctrl_killx;
  wire T124;
  reg  ex_reg_valid;
  wire T125;
  wire T126;
  wire replay_ex;
  wire T127;
  wire replay_ex_load_use;
  reg  ex_reg_load_use;
  wire T128;
  wire id_load_use;
  wire T129;
  wire T130;
  wire data_hazard_mem;
  wire T131;
  wire T132;
  wire T133;
  wire[4:0] mem_waddr;
  wire T134;
  wire T135;
  wire T136;
  wire[4:0] id_raddr_1;
  wire T137;
  wire T138;
  wire id_ctrl_rxs2;
  wire T139;
  wire T140;
  wire[31:0] T141;
  wire T142;
  wire T143;
  wire[31:0] T144;
  wire T145;
  wire[31:0] T146;
  wire T147;
  wire T148;
  wire[4:0] id_raddr_0;
  wire T149;
  wire T150;
  wire id_ctrl_rxs1;
  wire T151;
  wire T152;
  wire[31:0] T153;
  wire T154;
  wire T155;
  wire[31:0] T156;
  wire T157;
  wire T158;
  wire[31:0] T159;
  wire T160;
  wire[31:0] T161;
  wire wb_dcache_miss;
  wire T162;
  reg  wb_ctrl_mem;
  wire T163;
  wire replay_ex_structural;
  wire T164;
  wire T165;
  reg  ex_ctrl_div;
  wire T166;
  wire id_ctrl_div;
  wire T167;
  wire[31:0] T168;
  wire T169;
  wire T170;
  wire take_pc;
  wire take_pc_mem;
  wire T171;
  wire T172;
  wire mem_npc_misaligned;
  wire[39:0] mem_npc;
  wire[39:0] T173;
  wire[39:0] T174;
  wire[39:0] mem_br_target;
  wire[39:0] T919;
  wire[21:0] T175;
  wire[21:0] T176;
  wire[21:0] T177;
  wire[21:0] T178;
  wire[11:0] T179;
  wire[4:0] T180;
  wire[3:0] T181;
  wire[6:0] T182;
  wire[5:0] T183;
  wire T184;
  wire T185;
  wire[9:0] T186;
  wire[8:0] T187;
  wire[7:0] T188;
  wire[7:0] T189;
  wire T190;
  wire T191;
  reg  mem_ctrl_jal;
  wire T192;
  reg  ex_ctrl_jal;
  wire T193;
  wire id_ctrl_jal;
  wire[21:0] T920;
  wire[14:0] T194;
  wire[14:0] T195;
  wire[11:0] T196;
  wire[4:0] T197;
  wire[3:0] T198;
  wire[6:0] T199;
  wire[5:0] T200;
  wire T201;
  wire T202;
  wire[2:0] T203;
  wire[1:0] T204;
  wire T205;
  wire T206;
  wire[6:0] T921;
  wire T922;
  wire T207;
  wire mem_br_taken;
  reg [63:0] bypass_mux_1;
  wire[63:0] T208;
  reg  mem_ctrl_branch;
  wire T209;
  reg  ex_ctrl_branch;
  wire T210;
  wire id_ctrl_branch;
  wire T211;
  wire[31:0] T212;
  wire[17:0] T923;
  wire T924;
  wire[39:0] T213;
  reg [39:0] mem_reg_pc;
  wire[39:0] T214;
  reg [39:0] ex_reg_pc;
  wire[39:0] T215;
  wire[39:0] T216;
  wire[39:0] T217;
  wire[38:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire[1:0] T222;
  wire T223;
  wire[1:0] T224;
  wire T225;
  wire T226;
  wire[25:0] T227;
  wire[25:0] T228;
  wire T229;
  wire[25:0] T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  reg  mem_ctrl_jalr;
  wire T235;
  reg  ex_ctrl_jalr;
  wire T236;
  wire id_ctrl_jalr;
  wire T237;
  wire[31:0] T238;
  wire want_take_pc_mem;
  wire T239;
  reg  mem_reg_flush_pipe;
  wire T240;
  reg  ex_reg_flush_pipe;
  wire T241;
  wire T242;
  wire id_csr_flush;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire[11:0] T247;
  wire[11:0] id_csr_addr;
  wire T248;
  wire T249;
  wire id_csr_ren;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire id_system_insn;
  wire mem_misprediction;
  wire T254;
  wire T255;
  wire T256;
  wire mem_wrong_npc;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  reg  mem_reg_xcpt;
  wire T271;
  wire ex_xcpt;
  wire T272;
  reg  ex_ctrl_fp;
  wire T273;
  wire id_ctrl_fp;
  wire T274;
  reg  ex_reg_xcpt;
  wire T275;
  wire id_xcpt;
  wire id_illegal_insn;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire id_ctrl_legal;
  wire T284;
  wire T285;
  wire[31:0] T286;
  wire T287;
  wire T288;
  wire[31:0] T289;
  wire T290;
  wire T291;
  wire[31:0] T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire[31:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire[31:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[31:0] T305;
  wire T306;
  wire T307;
  wire[31:0] T308;
  wire T309;
  wire T310;
  wire[31:0] T311;
  wire T312;
  wire T313;
  wire[31:0] T314;
  wire T315;
  wire T316;
  wire[31:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[31:0] T321;
  wire T322;
  wire T323;
  wire[31:0] T324;
  wire T325;
  wire T326;
  wire[31:0] T327;
  wire T328;
  wire T329;
  wire[31:0] T330;
  wire T331;
  wire T332;
  wire[31:0] T333;
  wire T334;
  wire T335;
  wire[31:0] T336;
  wire T337;
  wire T338;
  wire[31:0] T339;
  wire T340;
  wire T341;
  wire[31:0] T342;
  wire T343;
  wire T344;
  wire[31:0] T345;
  wire T346;
  wire T347;
  wire[31:0] T348;
  wire T349;
  wire T350;
  wire[31:0] T351;
  wire T352;
  wire T353;
  wire[31:0] T354;
  wire T355;
  wire T356;
  wire T357;
  reg  ex_reg_xcpt_interrupt;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg  mem_reg_xcpt_interrupt;
  wire T362;
  wire T363;
  wire replay_mem;
  wire fpu_kill_mem;
  wire T364;
  reg  mem_ctrl_fp;
  wire T365;
  wire T366;
  reg  mem_reg_replay;
  wire T367;
  wire T368;
  wire dcache_kill_mem;
  wire T369;
  reg  wb_reg_valid;
  wire T370;
  wire ctrl_killm;
  wire T371;
  wire killm_common;
  wire T372;
  wire T373;
  wire T374;
  wire wb_set_sboard;
  wire T375;
  reg  wb_ctrl_div;
  wire T376;
  reg  mem_ctrl_div;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire[4:0] T386;
  wire[4:0] T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire[4:0] T393;
  wire[4:0] T394;
  wire T395;
  wire T396;
  wire id_wb_hazard;
  wire T397;
  wire fp_data_hazard_wb;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[4:0] id_raddr3;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  reg  wb_ctrl_wfd;
  wire T409;
  reg  mem_ctrl_wfd;
  wire T410;
  reg  ex_ctrl_wfd;
  wire T411;
  wire id_ctrl_wfd;
  wire T412;
  wire data_hazard_wb;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire id_mem_hazard;
  wire T422;
  wire fp_data_hazard_mem;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire mem_cannot_bypass;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  reg  mem_mem_cmd_bh;
  wire T439;
  wire ex_slow_bypass;
  wire T440;
  wire T441;
  reg [2:0] ex_ctrl_mem_type;
  wire[2:0] T442;
  wire[2:0] id_ctrl_mem_type;
  wire[2:0] T443;
  wire[1:0] T444;
  wire T445;
  wire[31:0] T446;
  wire T447;
  wire[31:0] T448;
  wire T449;
  wire[31:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  reg [4:0] ex_ctrl_mem_cmd;
  wire[4:0] T457;
  wire[4:0] id_ctrl_mem_cmd;
  wire[4:0] T458;
  wire[3:0] T459;
  wire[2:0] T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire[31:0] T464;
  wire T465;
  wire T466;
  wire[31:0] T467;
  wire T468;
  wire[31:0] T469;
  wire T470;
  wire T471;
  wire[31:0] T472;
  wire T473;
  wire[31:0] T474;
  wire T475;
  wire T476;
  wire[31:0] T477;
  wire T478;
  wire T479;
  wire[31:0] T480;
  wire T481;
  wire[31:0] T482;
  wire T483;
  reg [2:0] mem_ctrl_csr;
  wire[2:0] T484;
  reg [2:0] ex_ctrl_csr;
  wire[2:0] T485;
  wire[2:0] T486;
  wire[2:0] id_csr;
  wire id_ex_hazard;
  wire T487;
  wire fp_data_hazard_ex;
  wire T488;
  wire T489;
  wire T490;
  wire[4:0] ex_waddr;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire ex_cannot_bypass;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire data_hazard_ex;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[31:0] T518;
  wire[63:0] T519;
  reg [63:0] R520;
  reg [63:0] R521;
  wire[63:0] ex_rs_1;
  wire[63:0] T522;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire[1:0] T537;
  wire[63:0] id_rs_1;
  wire[63:0] T538;
  wire[63:0] T539;
  reg [63:0] T540 [30:0];
  wire[63:0] T541;
  wire T542;
  wire T543;
  wire[4:0] T544;
  wire T545;
  wire T546;
  wire[4:0] rf_waddr;
  wire rf_wen;
  wire[4:0] T547;
  wire[4:0] T548;
  wire[4:0] T549;
  wire[63:0] rf_wdata;
  wire[63:0] T550;
  wire[63:0] T551;
  reg [63:0] bypass_mux_2;
  wire[63:0] T552;
  wire[63:0] T553;
  wire[63:0] mem_int_wdata;
  wire[63:0] T554;
  wire[63:0] T555;
  wire[63:0] T925;
  wire[23:0] T926;
  wire T927;
  wire T556;
  wire T557;
  reg [2:0] wb_ctrl_csr;
  wire[2:0] T558;
  wire[63:0] ll_wdata;
  wire T559;
  wire dmem_resp_valid;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T571;
  wire[61:0] T572;
  wire[63:0] T573;
  wire[63:0] T574;
  wire T575;
  wire[1:0] T576;
  wire[63:0] T577;
  wire T578;
  wire T579;
  reg  ex_reg_rs_bypass_1;
  wire T580;
  wire[4:0] T581;
  wire[4:0] T582;
  wire[63:0] T583;
  reg [63:0] R584;
  reg [63:0] R585;
  wire[63:0] ex_rs_0;
  wire[63:0] T586;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire[1:0] T597;
  wire[63:0] id_rs_0;
  wire[63:0] T598;
  wire[63:0] T599;
  wire[4:0] T600;
  wire[4:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T612;
  wire[61:0] T613;
  wire[63:0] T614;
  wire[63:0] T615;
  wire T616;
  wire[1:0] T617;
  wire[63:0] T618;
  wire T619;
  wire T620;
  reg  ex_reg_rs_bypass_0;
  wire T621;
  wire[4:0] T622;
  wire[4:0] T623;
  wire T624;
  wire[63:0] T625;
  wire[4:0] T626;
  wire[4:0] T627;
  wire[39:0] T628;
  reg [39:0] wb_reg_pc;
  wire[39:0] T629;
  wire T630;
  wire[32:0] T631;
  wire[32:0] T632;
  wire T633;
  wire[1127:0] T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  reg  R639;
  wire T640;
  reg  ex_ctrl_alu_dw;
  wire T641;
  wire id_ctrl_alu_dw;
  wire T642;
  wire T643;
  wire[31:0] T644;
  wire T645;
  wire[31:0] T646;
  reg [3:0] ex_ctrl_alu_fn;
  wire[3:0] T647;
  wire[3:0] id_ctrl_alu_fn;
  wire[3:0] T648;
  wire[2:0] T649;
  wire[1:0] T650;
  wire T651;
  wire T652;
  wire[31:0] T653;
  wire T654;
  wire T655;
  wire[31:0] T656;
  wire T657;
  wire[31:0] T658;
  wire T659;
  wire T660;
  wire[31:0] T661;
  wire T662;
  wire T663;
  wire[31:0] T664;
  wire T665;
  wire T666;
  wire[31:0] T667;
  wire T668;
  wire T669;
  wire[31:0] T670;
  wire T671;
  wire[31:0] T672;
  wire T673;
  wire T674;
  wire[31:0] T675;
  wire T676;
  wire T677;
  wire[31:0] T678;
  wire T679;
  wire T680;
  wire[31:0] T681;
  wire T682;
  wire[31:0] T683;
  wire T684;
  wire T685;
  wire[31:0] T686;
  wire T687;
  wire T688;
  wire T689;
  wire[31:0] T690;
  wire T691;
  wire[63:0] T692;
  wire[63:0] ex_op1;
  wire[63:0] T928;
  wire[39:0] T693;
  wire[39:0] T694;
  wire T695;
  reg [1:0] ex_ctrl_sel_alu1;
  wire[1:0] T696;
  wire[1:0] id_ctrl_sel_alu1;
  wire[1:0] T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[31:0] T702;
  wire T703;
  wire T704;
  wire[31:0] T705;
  wire[23:0] T929;
  wire T930;
  wire[63:0] T706;
  wire T707;
  wire[63:0] T708;
  wire[63:0] ex_op2;
  wire[63:0] T931;
  wire[31:0] T709;
  wire[31:0] T932;
  wire[3:0] T710;
  wire T711;
  reg [1:0] ex_ctrl_sel_alu2;
  wire[1:0] T712;
  wire[1:0] id_ctrl_sel_alu2;
  wire[1:0] T713;
  wire T714;
  wire T715;
  wire[31:0] T716;
  wire T717;
  wire T718;
  wire T719;
  wire T720;
  wire[31:0] T721;
  wire T722;
  wire[31:0] T723;
  wire T724;
  wire T725;
  wire[31:0] T726;
  wire T727;
  wire T728;
  wire T729;
  wire[31:0] T730;
  wire[27:0] T933;
  wire T934;
  wire[31:0] ex_imm;
  wire[31:0] T731;
  wire[11:0] T732;
  wire[4:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  reg [2:0] ex_ctrl_sel_imm;
  wire[2:0] T739;
  wire[2:0] id_ctrl_sel_imm;
  wire[2:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire[31:0] T744;
  wire T745;
  wire[31:0] T746;
  wire T747;
  wire T748;
  wire[31:0] T749;
  wire T750;
  wire T751;
  wire[31:0] T752;
  wire T753;
  wire T754;
  wire[31:0] T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire[3:0] T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire[3:0] T764;
  wire T765;
  wire[3:0] T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire[6:0] T771;
  wire[5:0] T772;
  wire[5:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire T792;
  wire[19:0] T793;
  wire[18:0] T794;
  wire[7:0] T795;
  wire[7:0] T796;
  wire[7:0] T797;
  wire[7:0] T935;
  wire T798;
  wire T799;
  wire T800;
  wire[10:0] T801;
  wire[10:0] T936;
  wire[10:0] T802;
  wire[10:0] T803;
  wire T804;
  wire T805;
  wire[31:0] T937;
  wire T938;
  wire[63:0] T806;
  wire T807;
  reg [63:0] wb_reg_cause;
  wire[63:0] T808;
  wire[63:0] mem_cause;
  wire[63:0] T939;
  wire[2:0] T809;
  wire[2:0] T810;
  wire[2:0] T811;
  wire[2:0] T812;
  reg [63:0] mem_reg_cause;
  wire[63:0] T813;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T814;
  wire[63:0] id_cause;
  wire[63:0] T940;
  wire[1:0] T815;
  wire[2:0] T816;
  wire[11:0] T817;
  wire T818;
  wire T819;
  wire T820;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T821;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T822;
  wire T823;
  wire T824;
  wire T825;
  reg  ex_ctrl_rxs2;
  wire T826;
  wire T827;
  wire[6:0] T828;
  wire[4:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[4:0] T833;
  wire[4:0] T834;
  wire[6:0] T835;
  wire wb_rocc_val;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire T840;
  wire dmem_resp_fpu;
  wire T841;
  wire[63:0] T842;
  wire T843;
  wire[8:0] T941;
  wire[5:0] T844;
  wire[39:0] T845;
  wire[39:0] T846;
  wire[38:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[1:0] T851;
  wire T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire[25:0] T856;
  wire[25:0] T857;
  wire T858;
  wire[25:0] T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  reg  wb_ctrl_fence_i;
  wire T866;
  reg  mem_ctrl_fence_i;
  wire T867;
  reg  ex_ctrl_fence_i;
  wire T868;
  wire[38:0] T942;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[38:0] T943;
  wire T876;
  wire T877;
  wire T878;
  wire[38:0] T944;
  wire T879;
  wire T880;
  wire[4:0] T881;
  wire[4:0] T882;
  wire T883;
  wire[38:0] T945;
  wire[38:0] T946;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T884;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T885;
  wire T886;
  wire T887;
  reg  ex_reg_btb_hit;
  wire T888;
  reg [3:0] mem_reg_btb_resp_bht_history;
  wire[3:0] T889;
  reg [3:0] ex_reg_btb_resp_bht_history;
  wire[3:0] T890;
  reg [2:0] mem_reg_btb_resp_entry;
  wire[2:0] T891;
  reg [2:0] ex_reg_btb_resp_entry;
  wire[2:0] T892;
  reg [38:0] mem_reg_btb_resp_target;
  wire[38:0] T893;
  reg [38:0] ex_reg_btb_resp_target;
  wire[38:0] T894;
  reg  mem_reg_btb_resp_bridx;
  wire T895;
  reg  ex_reg_btb_resp_bridx;
  wire T896;
  reg  mem_reg_btb_resp_mask;
  wire T897;
  reg  ex_reg_btb_resp_mask;
  wire T898;
  reg  mem_reg_btb_resp_taken;
  wire T899;
  reg  ex_reg_btb_resp_taken;
  wire T900;
  reg  mem_reg_btb_hit;
  wire T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire T912;
  wire[39:0] T913;
  wire[39:0] T914;
  wire[39:0] T915;
  wire T916;
  wire csr_io_host_csr_req_ready;
  wire csr_io_host_csr_resp_valid;
  wire[63:0] csr_io_host_csr_resp_bits;
  wire csr_io_host_debug_stats_csr;
  wire[63:0] csr_io_rw_rdata;
  wire csr_io_csr_stall;
  wire csr_io_csr_xcpt;
  wire csr_io_eret;
  wire csr_io_status_sd;
  wire[30:0] csr_io_status_zero2;
  wire csr_io_status_sd_rv32;
  wire[8:0] csr_io_status_zero1;
  wire[4:0] csr_io_status_vm;
  wire csr_io_status_mprv;
  wire[1:0] csr_io_status_xs;
  wire[1:0] csr_io_status_fs;
  wire[1:0] csr_io_status_prv3;
  wire csr_io_status_ie3;
  wire[1:0] csr_io_status_prv2;
  wire csr_io_status_ie2;
  wire[1:0] csr_io_status_prv1;
  wire csr_io_status_ie1;
  wire[1:0] csr_io_status_prv;
  wire csr_io_status_ie;
  wire[31:0] csr_io_ptbr;
  wire[39:0] csr_io_evec;
  wire csr_io_fatc;
  wire[63:0] csr_io_time;
  wire[2:0] csr_io_fcsr_rm;
  wire csr_io_interrupt;
  wire[63:0] csr_io_interrupt_cause;
  wire[63:0] alu_io_out;
  wire[63:0] alu_io_adder_out;
  wire div_io_req_ready;
  wire div_io_resp_valid;
  wire[63:0] div_io_resp_bits_data;
  wire[4:0] div_io_resp_bits_tag;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    id_reg_fence = {1{$random}};
    R73 = {1{$random}};
    wb_ctrl_wxd = {1{$random}};
    mem_ctrl_wxd = {1{$random}};
    ex_ctrl_wxd = {1{$random}};
    wb_ctrl_rocc = {1{$random}};
    mem_ctrl_rocc = {1{$random}};
    ex_ctrl_rocc = {1{$random}};
    wb_reg_replay = {1{$random}};
    wb_reg_xcpt = {1{$random}};
    mem_ctrl_mem = {1{$random}};
    ex_ctrl_mem = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    ex_reg_load_use = {1{$random}};
    wb_ctrl_mem = {1{$random}};
    ex_ctrl_div = {1{$random}};
    mem_ctrl_jal = {1{$random}};
    ex_ctrl_jal = {1{$random}};
    bypass_mux_1 = {2{$random}};
    mem_ctrl_branch = {1{$random}};
    ex_ctrl_branch = {1{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    mem_ctrl_jalr = {1{$random}};
    ex_ctrl_jalr = {1{$random}};
    mem_reg_flush_pipe = {1{$random}};
    ex_reg_flush_pipe = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_ctrl_fp = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    mem_ctrl_fp = {1{$random}};
    mem_reg_replay = {1{$random}};
    wb_reg_valid = {1{$random}};
    wb_ctrl_div = {1{$random}};
    mem_ctrl_div = {1{$random}};
    wb_ctrl_wfd = {1{$random}};
    mem_ctrl_wfd = {1{$random}};
    ex_ctrl_wfd = {1{$random}};
    mem_mem_cmd_bh = {1{$random}};
    ex_ctrl_mem_type = {1{$random}};
    ex_ctrl_mem_cmd = {1{$random}};
    mem_ctrl_csr = {1{$random}};
    ex_ctrl_csr = {1{$random}};
    R520 = {2{$random}};
    R521 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T540[initvar] = {2{$random}};
    bypass_mux_2 = {2{$random}};
    wb_ctrl_csr = {1{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R584 = {2{$random}};
    R585 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    R639 = {1{$random}};
    ex_ctrl_alu_dw = {1{$random}};
    ex_ctrl_alu_fn = {1{$random}};
    ex_ctrl_sel_alu1 = {1{$random}};
    ex_ctrl_sel_alu2 = {1{$random}};
    ex_ctrl_sel_imm = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
    ex_ctrl_rxs2 = {1{$random}};
    wb_ctrl_fence_i = {1{$random}};
    mem_ctrl_fence_i = {1{$random}};
    ex_ctrl_fence_i = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_history = {1{$random}};
    ex_reg_btb_resp_bht_history = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_bridx = {1{$random}};
    ex_reg_btb_resp_bridx = {1{$random}};
    mem_reg_btb_resp_mask = {1{$random}};
    ex_reg_btb_resp_mask = {1{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_rocc_dma_resp_bits_status = {1{$random}};
//  assign io_rocc_dma_resp_bits_client_xact_id = {1{$random}};
//  assign io_rocc_dma_resp_valid = {1{$random}};
//  assign io_rocc_dma_req_ready = {1{$random}};
//  assign io_rocc_fpu_resp_bits_exc = {1{$random}};
//  assign io_rocc_fpu_resp_bits_data = {3{$random}};
//  assign io_rocc_fpu_resp_valid = {1{$random}};
//  assign io_rocc_fpu_req_ready = {1{$random}};
//  assign io_rocc_pptw_invalidate = {1{$random}};
//  assign io_rocc_pptw_status_ie = {1{$random}};
//  assign io_rocc_pptw_status_prv = {1{$random}};
//  assign io_rocc_pptw_status_ie1 = {1{$random}};
//  assign io_rocc_pptw_status_prv1 = {1{$random}};
//  assign io_rocc_pptw_status_ie2 = {1{$random}};
//  assign io_rocc_pptw_status_prv2 = {1{$random}};
//  assign io_rocc_pptw_status_ie3 = {1{$random}};
//  assign io_rocc_pptw_status_prv3 = {1{$random}};
//  assign io_rocc_pptw_status_fs = {1{$random}};
//  assign io_rocc_pptw_status_xs = {1{$random}};
//  assign io_rocc_pptw_status_mprv = {1{$random}};
//  assign io_rocc_pptw_status_vm = {1{$random}};
//  assign io_rocc_pptw_status_zero1 = {1{$random}};
//  assign io_rocc_pptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_pptw_status_zero2 = {1{$random}};
//  assign io_rocc_pptw_status_sd = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_pptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_pptw_resp_bits_error = {1{$random}};
//  assign io_rocc_pptw_resp_valid = {1{$random}};
//  assign io_rocc_pptw_req_ready = {1{$random}};
//  assign io_rocc_dptw_invalidate = {1{$random}};
//  assign io_rocc_dptw_status_ie = {1{$random}};
//  assign io_rocc_dptw_status_prv = {1{$random}};
//  assign io_rocc_dptw_status_ie1 = {1{$random}};
//  assign io_rocc_dptw_status_prv1 = {1{$random}};
//  assign io_rocc_dptw_status_ie2 = {1{$random}};
//  assign io_rocc_dptw_status_prv2 = {1{$random}};
//  assign io_rocc_dptw_status_ie3 = {1{$random}};
//  assign io_rocc_dptw_status_prv3 = {1{$random}};
//  assign io_rocc_dptw_status_fs = {1{$random}};
//  assign io_rocc_dptw_status_xs = {1{$random}};
//  assign io_rocc_dptw_status_mprv = {1{$random}};
//  assign io_rocc_dptw_status_vm = {1{$random}};
//  assign io_rocc_dptw_status_zero1 = {1{$random}};
//  assign io_rocc_dptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_dptw_status_zero2 = {1{$random}};
//  assign io_rocc_dptw_status_sd = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_dptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_dptw_resp_bits_error = {1{$random}};
//  assign io_rocc_dptw_resp_valid = {1{$random}};
//  assign io_rocc_dptw_req_ready = {1{$random}};
//  assign io_rocc_iptw_invalidate = {1{$random}};
//  assign io_rocc_iptw_status_ie = {1{$random}};
//  assign io_rocc_iptw_status_prv = {1{$random}};
//  assign io_rocc_iptw_status_ie1 = {1{$random}};
//  assign io_rocc_iptw_status_prv1 = {1{$random}};
//  assign io_rocc_iptw_status_ie2 = {1{$random}};
//  assign io_rocc_iptw_status_prv2 = {1{$random}};
//  assign io_rocc_iptw_status_ie3 = {1{$random}};
//  assign io_rocc_iptw_status_prv3 = {1{$random}};
//  assign io_rocc_iptw_status_fs = {1{$random}};
//  assign io_rocc_iptw_status_xs = {1{$random}};
//  assign io_rocc_iptw_status_mprv = {1{$random}};
//  assign io_rocc_iptw_status_vm = {1{$random}};
//  assign io_rocc_iptw_status_zero1 = {1{$random}};
//  assign io_rocc_iptw_status_sd_rv32 = {1{$random}};
//  assign io_rocc_iptw_status_zero2 = {1{$random}};
//  assign io_rocc_iptw_status_sd = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_v = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_typ = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_r = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_d = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_reserved_for_software = {1{$random}};
//  assign io_rocc_iptw_resp_bits_pte_ppn = {1{$random}};
//  assign io_rocc_iptw_resp_bits_error = {1{$random}};
//  assign io_rocc_iptw_resp_valid = {1{$random}};
//  assign io_rocc_iptw_req_ready = {1{$random}};
//  assign io_rocc_autl_grant_bits_data = {4{$random}};
//  assign io_rocc_autl_grant_bits_g_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_is_builtin_type = {1{$random}};
//  assign io_rocc_autl_grant_bits_manager_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_client_xact_id = {1{$random}};
//  assign io_rocc_autl_grant_bits_addr_beat = {1{$random}};
//  assign io_rocc_autl_grant_valid = {1{$random}};
//  assign io_rocc_autl_acquire_ready = {1{$random}};
//  assign io_rocc_mem_ordered = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_st = {1{$random}};
//  assign io_rocc_mem_xcpt_pf_ld = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_st = {1{$random}};
//  assign io_rocc_mem_xcpt_ma_ld = {1{$random}};
//  assign io_rocc_mem_replay_next_bits = {1{$random}};
//  assign io_rocc_mem_replay_next_valid = {1{$random}};
//  assign io_rocc_mem_resp_bits_store_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_data_word_bypass = {2{$random}};
//  assign io_rocc_mem_resp_bits_has_data = {1{$random}};
//  assign io_rocc_mem_resp_bits_replay = {1{$random}};
//  assign io_rocc_mem_resp_bits_nack = {1{$random}};
//  assign io_rocc_mem_resp_bits_data = {2{$random}};
//  assign io_rocc_mem_resp_bits_typ = {1{$random}};
//  assign io_rocc_mem_resp_bits_cmd = {1{$random}};
//  assign io_rocc_mem_resp_bits_tag = {1{$random}};
//  assign io_rocc_mem_resp_bits_addr = {2{$random}};
//  assign io_rocc_mem_resp_valid = {1{$random}};
//  assign io_rocc_mem_req_ready = {1{$random}};
//  assign io_rocc_resp_ready = {1{$random}};
//  assign io_fpu_cp_resp_ready = {1{$random}};
//  assign io_fpu_cp_req_bits_in3 = {3{$random}};
//  assign io_fpu_cp_req_bits_in2 = {3{$random}};
//  assign io_fpu_cp_req_bits_in1 = {3{$random}};
//  assign io_fpu_cp_req_bits_typ = {1{$random}};
//  assign io_fpu_cp_req_bits_rm = {1{$random}};
//  assign io_fpu_cp_req_bits_wflags = {1{$random}};
//  assign io_fpu_cp_req_bits_round = {1{$random}};
//  assign io_fpu_cp_req_bits_sqrt = {1{$random}};
//  assign io_fpu_cp_req_bits_div = {1{$random}};
//  assign io_fpu_cp_req_bits_fma = {1{$random}};
//  assign io_fpu_cp_req_bits_fastpipe = {1{$random}};
//  assign io_fpu_cp_req_bits_toint = {1{$random}};
//  assign io_fpu_cp_req_bits_fromint = {1{$random}};
//  assign io_fpu_cp_req_bits_single = {1{$random}};
//  assign io_fpu_cp_req_bits_swap23 = {1{$random}};
//  assign io_fpu_cp_req_bits_swap12 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren3 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren2 = {1{$random}};
//  assign io_fpu_cp_req_bits_ren1 = {1{$random}};
//  assign io_fpu_cp_req_bits_wen = {1{$random}};
//  assign io_fpu_cp_req_bits_ldst = {1{$random}};
//  assign io_fpu_cp_req_bits_cmd = {1{$random}};
//  assign io_fpu_cp_req_valid = {1{$random}};
//  assign io_imem_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T516 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T515 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign T5 = T6 | csr_io_interrupt;
  assign T6 = ctrl_killd ^ 1'h1;
  assign ctrl_killd = T7;
  assign T7 = T8 | csr_io_interrupt;
  assign T8 = T513 | ctrl_stalld;
  assign ctrl_stalld = T9 | csr_io_csr_stall;
  assign T9 = T51 | id_do_fence;
  assign id_do_fence = id_mem_busy & T10;
  assign T10 = T19 | id_csr_en;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_ctrl_csr = T11;
  assign T11 = {T17, T12};
  assign T12 = {T15, T13};
  assign T13 = T14 == 32'h1050;
  assign T14 = io_imem_resp_bits_data_0 & 32'h1050;
  assign T15 = T16 == 32'h2050;
  assign T16 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T17 = T18 == 32'h50;
  assign T18 = io_imem_resp_bits_data_0 & 32'h3050;
  assign T19 = T46 | T20;
  assign T20 = id_reg_fence & T21;
  assign T21 = id_ctrl_mem | id_ctrl_rocc;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_mem = T22;
  assign T22 = T25 | T23;
  assign T23 = T24 == 32'h1000202f;
  assign T24 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h800202f;
  assign T27 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h202f;
  assign T30 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h3;
  assign T33 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T34 = T37 | T35;
  assign T35 = T36 == 32'h3;
  assign T36 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T37 = T38 == 32'h3;
  assign T38 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T917 = reset ? 1'h0 : T39;
  assign T39 = id_fence_next | T40;
  assign T40 = id_reg_fence & id_mem_busy;
  assign id_fence_next = id_ctrl_fence | T41;
  assign T41 = id_ctrl_amo & id_amo_rl;
  assign id_amo_rl = io_imem_resp_bits_data_0[5'h19:5'h19];
  assign id_ctrl_amo = T42;
  assign T42 = T43 == 32'h2008;
  assign T43 = io_imem_resp_bits_data_0 & 32'h6048;
  assign id_ctrl_fence = T44;
  assign T44 = T45 == 32'h8;
  assign T45 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T46 = T49 | id_ctrl_fence_i;
  assign id_ctrl_fence_i = T47;
  assign T47 = T48 == 32'h1008;
  assign T48 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T49 = id_ctrl_amo & id_amo_aq;
  assign id_amo_aq = io_imem_resp_bits_data_0[5'h1a:5'h1a];
  assign id_mem_busy = T50 | io_dmem_req_valid;
  assign T50 = io_dmem_ordered ^ 1'h1;
  assign T51 = T54 | T52;
  assign T52 = id_ctrl_mem & T53;
  assign T53 = io_dmem_req_ready ^ 1'h1;
  assign T54 = T396 | id_sboard_hazard;
  assign id_sboard_hazard = T381 | T55;
  assign T55 = T379 & T56;
  assign T56 = T61 & T57;
  assign T57 = T58 - 1'h1;
  assign T58 = 1'h1 << T59;
  assign T59 = T60 + 5'h1;
  assign T60 = id_waddr - id_waddr;
  assign id_waddr = io_imem_resp_bits_data_0[4'hb:3'h7];
  assign T61 = T62 >> id_waddr;
  assign T62 = R73 & T63;
  assign T63 = ~ T64;
  assign T64 = ll_wen ? T65 : 32'h0;
  assign T65 = 1'h1 << ll_waddr;
  assign ll_waddr = T66;
  assign T66 = T68 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign dmem_resp_waddr = T67[3'h5:1'h1];
  assign T67 = io_dmem_resp_bits_tag;
  assign T68 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_xpu = T69 ^ 1'h1;
  assign T69 = T70;
  assign T70 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign ll_wen = T71;
  assign T71 = T68 ? 1'h1 : T72;
  assign T72 = T635 & div_io_resp_valid;
  assign T918 = reset ? 32'h0 : T74;
  assign T74 = T378 ? T76 : T75;
  assign T75 = ll_wen ? T62 : R73;
  assign T76 = T62 | T77;
  assign T77 = T79 ? T78 : 32'h0;
  assign T78 = 1'h1 << wb_waddr;
  assign wb_waddr = wb_reg_inst[4'hb:3'h7];
  assign T79 = wb_set_sboard & wb_wen;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign T80 = T516 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign T81 = T515 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign T82 = T103 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign id_ctrl_wxd = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h0;
  assign T85 = io_imem_resp_bits_data_0 & 32'h28;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h2010;
  assign T88 = io_imem_resp_bits_data_0 & 32'h2010;
  assign T89 = T92 | T90;
  assign T90 = T91 == 32'h2008;
  assign T91 = io_imem_resp_bits_data_0 & 32'h2008;
  assign T92 = T95 | T93;
  assign T93 = T94 == 32'h1010;
  assign T94 = io_imem_resp_bits_data_0 & 32'h1010;
  assign T95 = T98 | T96;
  assign T96 = T97 == 32'h48;
  assign T97 = io_imem_resp_bits_data_0 & 32'h48;
  assign T98 = T101 | T99;
  assign T99 = T100 == 32'h10;
  assign T100 = io_imem_resp_bits_data_0 & 32'h50;
  assign T101 = T102 == 32'h4;
  assign T102 = io_imem_resp_bits_data_0 & 32'hc;
  assign T103 = ctrl_killd ^ 1'h1;
  assign wb_valid = T105 & T104;
  assign T104 = csr_io_csr_xcpt ^ 1'h1;
  assign T105 = wb_reg_valid & T106;
  assign T106 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T107;
  assign T107 = T109 & T108;
  assign T108 = io_rocc_cmd_ready ^ 1'h1;
  assign T109 = wb_reg_valid & wb_ctrl_rocc;
  assign T110 = T516 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign T111 = T515 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign T112 = T103 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign replay_wb_common = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T113 = replay_mem & T114;
  assign T114 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T115;
  assign T115 = T116 | csr_io_eret;
  assign T116 = replay_wb | wb_xcpt;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T117 = mem_xcpt & T118;
  assign T118 = take_pc_wb ^ 1'h1;
  assign mem_xcpt = T259 | T119;
  assign T119 = T120 & io_dmem_xcpt_pf_ld;
  assign T120 = mem_reg_valid & mem_ctrl_mem;
  assign T121 = T515 ? ex_ctrl_mem : mem_ctrl_mem;
  assign T122 = T103 ? id_ctrl_mem : ex_ctrl_mem;
  assign T123 = ctrl_killx ^ 1'h1;
  assign ctrl_killx = T126 | T124;
  assign T124 = ex_reg_valid ^ 1'h1;
  assign T125 = ctrl_killd ^ 1'h1;
  assign T126 = take_pc | replay_ex;
  assign replay_ex = ex_reg_valid & T127;
  assign T127 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T128 = T103 ? id_load_use : ex_reg_load_use;
  assign id_load_use = T129;
  assign T129 = T130 & mem_ctrl_mem;
  assign T130 = mem_reg_valid & data_hazard_mem;
  assign data_hazard_mem = mem_ctrl_wxd & T131;
  assign T131 = T134 | T132;
  assign T132 = T379 & T133;
  assign T133 = id_waddr == mem_waddr;
  assign mem_waddr = mem_reg_inst[4'hb:3'h7];
  assign T134 = T147 | T135;
  assign T135 = T137 & T136;
  assign T136 = id_raddr_1 == mem_waddr;
  assign id_raddr_1 = io_imem_resp_bits_data_0[5'h18:5'h14];
  assign T137 = id_ctrl_rxs2 & T138;
  assign T138 = id_raddr_1 != 5'h0;
  assign id_ctrl_rxs2 = T139;
  assign T139 = T142 | T140;
  assign T140 = T141 == 32'h20;
  assign T141 = io_imem_resp_bits_data_0 & 32'h34;
  assign T142 = T145 | T143;
  assign T143 = T144 == 32'h20;
  assign T144 = io_imem_resp_bits_data_0 & 32'h64;
  assign T145 = T146 == 32'h20;
  assign T146 = io_imem_resp_bits_data_0 & 32'h70;
  assign T147 = T149 & T148;
  assign T148 = id_raddr_0 == mem_waddr;
  assign id_raddr_0 = io_imem_resp_bits_data_0[5'h13:4'hf];
  assign T149 = id_ctrl_rxs1 & T150;
  assign T150 = id_raddr_0 != 5'h0;
  assign id_ctrl_rxs1 = T151;
  assign T151 = T154 | T152;
  assign T152 = T153 == 32'h2000;
  assign T153 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T154 = T157 | T155;
  assign T155 = T156 == 32'h0;
  assign T156 = io_imem_resp_bits_data_0 & 32'h18;
  assign T157 = T160 | T158;
  assign T158 = T159 == 32'h0;
  assign T159 = io_imem_resp_bits_data_0 & 32'h44;
  assign T160 = T161 == 32'h0;
  assign T161 = io_imem_resp_bits_data_0 & 32'h4004;
  assign wb_dcache_miss = wb_ctrl_mem & T162;
  assign T162 = io_dmem_resp_valid ^ 1'h1;
  assign T163 = T516 ? mem_ctrl_mem : wb_ctrl_mem;
  assign replay_ex_structural = T169 | T164;
  assign T164 = ex_ctrl_div & T165;
  assign T165 = div_io_req_ready ^ 1'h1;
  assign T166 = T103 ? id_ctrl_div : ex_ctrl_div;
  assign id_ctrl_div = T167;
  assign T167 = T168 == 32'h2000030;
  assign T168 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T169 = ex_ctrl_mem & T170;
  assign T170 = io_dmem_req_ready ^ 1'h1;
  assign take_pc = take_pc_wb | take_pc_mem;
  assign take_pc_mem = T171;
  assign T171 = want_take_pc_mem & T172;
  assign T172 = mem_npc_misaligned ^ 1'h1;
  assign mem_npc_misaligned = mem_npc[1'h1:1'h1];
  assign mem_npc = T173;
  assign T173 = T174 & 40'hfffffffffe;
  assign T174 = mem_ctrl_jalr ? T216 : mem_br_target;
  assign mem_br_target = T213 + T919;
  assign T919 = {T923, T175};
  assign T175 = T207 ? T920 : T176;
  assign T176 = mem_ctrl_jal ? T177 : 22'h4;
  assign T177 = T178;
  assign T178 = {T186, T179};
  assign T179 = {T182, T180};
  assign T180 = {T181, 1'h0};
  assign T181 = mem_reg_inst[5'h18:5'h15];
  assign T182 = {T184, T183};
  assign T183 = mem_reg_inst[5'h1e:5'h19];
  assign T184 = T185;
  assign T185 = mem_reg_inst[5'h14:5'h14];
  assign T186 = {T190, T187};
  assign T187 = {T190, T188};
  assign T188 = T189;
  assign T189 = mem_reg_inst[5'h13:4'hc];
  assign T190 = T191;
  assign T191 = mem_reg_inst[5'h1f:5'h1f];
  assign T192 = T515 ? ex_ctrl_jal : mem_ctrl_jal;
  assign T193 = T103 ? id_ctrl_jal : ex_ctrl_jal;
  assign id_ctrl_jal = T96;
  assign T920 = {T921, T194};
  assign T194 = T195;
  assign T195 = {T203, T196};
  assign T196 = {T199, T197};
  assign T197 = {T198, 1'h0};
  assign T198 = mem_reg_inst[4'hb:4'h8];
  assign T199 = {T201, T200};
  assign T200 = mem_reg_inst[5'h1e:5'h19];
  assign T201 = T202;
  assign T202 = mem_reg_inst[3'h7:3'h7];
  assign T203 = {T205, T204};
  assign T204 = {T205, T205};
  assign T205 = T206;
  assign T206 = mem_reg_inst[5'h1f:5'h1f];
  assign T921 = T922 ? 7'h7f : 7'h0;
  assign T922 = T194[4'he:4'he];
  assign T207 = mem_ctrl_branch & mem_br_taken;
  assign mem_br_taken = bypass_mux_1[1'h0:1'h0];
  assign T208 = T515 ? alu_io_out : bypass_mux_1;
  assign T209 = T515 ? ex_ctrl_branch : mem_ctrl_branch;
  assign T210 = T103 ? id_ctrl_branch : ex_ctrl_branch;
  assign id_ctrl_branch = T211;
  assign T211 = T212 == 32'h40;
  assign T212 = io_imem_resp_bits_data_0 & 32'h54;
  assign T923 = T924 ? 18'h3ffff : 18'h0;
  assign T924 = T175[5'h15:5'h15];
  assign T213 = mem_reg_pc;
  assign T214 = T515 ? ex_reg_pc : mem_reg_pc;
  assign T215 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T216 = T217;
  assign T217 = {T219, T218};
  assign T218 = bypass_mux_1[6'h26:1'h0];
  assign T219 = T232 ? T231 : T220;
  assign T220 = T225 ? T223 : T221;
  assign T221 = T222[1'h0:1'h0];
  assign T222 = bypass_mux_1[6'h27:6'h26];
  assign T223 = T224 == 2'h3;
  assign T224 = T222;
  assign T225 = T229 | T226;
  assign T226 = T227 == 26'h3fffffe;
  assign T227 = T228;
  assign T228 = bypass_mux_1 >> 6'h26;
  assign T229 = T230 == 26'h3ffffff;
  assign T230 = T228;
  assign T231 = T222 != 2'h0;
  assign T232 = T234 | T233;
  assign T233 = T228 == 26'h1;
  assign T234 = T228 == 26'h0;
  assign T235 = T515 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign T236 = T103 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign id_ctrl_jalr = T237;
  assign T237 = T238 == 32'h4;
  assign T238 = io_imem_resp_bits_data_0 & 32'h1c;
  assign want_take_pc_mem = mem_reg_valid & T239;
  assign T239 = mem_misprediction | mem_reg_flush_pipe;
  assign T240 = T515 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign T241 = T103 ? T242 : ex_reg_flush_pipe;
  assign T242 = id_ctrl_fence_i | id_csr_flush;
  assign id_csr_flush = id_system_insn | T243;
  assign T243 = T248 & T244;
  assign T244 = T245 ^ 1'h1;
  assign T245 = T246;
  assign T246 = T247 == 12'h40;
  assign T247 = id_csr_addr & 12'h8c4;
  assign id_csr_addr = io_imem_resp_bits_data_0[5'h1f:5'h14];
  assign T248 = id_csr_en & T249;
  assign T249 = id_csr_ren ^ 1'h1;
  assign id_csr_ren = T251 & T250;
  assign T250 = id_raddr_0 == 5'h0;
  assign T251 = T253 | T252;
  assign T252 = id_ctrl_csr == 3'h3;
  assign T253 = id_ctrl_csr == 3'h2;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign mem_misprediction = T256 & T254;
  assign T254 = T255 | mem_ctrl_jal;
  assign T255 = mem_ctrl_branch | mem_ctrl_jalr;
  assign T256 = mem_wrong_npc & mem_reg_valid;
  assign mem_wrong_npc = T258 | T257;
  assign T257 = ex_reg_valid ^ 1'h1;
  assign T258 = mem_npc != ex_reg_pc;
  assign T259 = T262 | T260;
  assign T260 = T261 & io_dmem_xcpt_pf_st;
  assign T261 = mem_reg_valid & mem_ctrl_mem;
  assign T262 = T265 | T263;
  assign T263 = T264 & io_dmem_xcpt_ma_ld;
  assign T264 = mem_reg_valid & mem_ctrl_mem;
  assign T265 = T268 | T266;
  assign T266 = T267 & io_dmem_xcpt_ma_st;
  assign T267 = mem_reg_valid & mem_ctrl_mem;
  assign T268 = T270 | T269;
  assign T269 = want_take_pc_mem & mem_npc_misaligned;
  assign T270 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T271 = T361 & ex_xcpt;
  assign ex_xcpt = T274 | T272;
  assign T272 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign T273 = T103 ? id_ctrl_fp : ex_ctrl_fp;
  assign id_ctrl_fp = 1'h0;
  assign T274 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T275 = T357 & id_xcpt;
  assign id_xcpt = T356 | id_illegal_insn;
  assign id_illegal_insn = T279 | T276;
  assign T276 = id_ctrl_rocc & T277;
  assign T277 = T278 ^ 1'h1;
  assign T278 = csr_io_status_xs != 2'h0;
  assign T279 = T283 | T280;
  assign T280 = id_ctrl_fp & T281;
  assign T281 = T282 ^ 1'h1;
  assign T282 = csr_io_status_fs != 2'h0;
  assign T283 = id_ctrl_legal ^ 1'h1;
  assign id_ctrl_legal = T284;
  assign T284 = T287 | T285;
  assign T285 = T286 == 32'h33;
  assign T286 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T287 = T290 | T288;
  assign T288 = T289 == 32'h4063;
  assign T289 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T290 = T293 | T291;
  assign T291 = T292 == 32'h1063;
  assign T292 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T293 = T295 | T294;
  assign T294 = io_imem_resp_bits_data_0 == 32'h30500073;
  assign T295 = T298 | T296;
  assign T296 = T297 == 32'h10100073;
  assign T297 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T298 = T299 | T23;
  assign T299 = T302 | T300;
  assign T300 = T301 == 32'h10000073;
  assign T301 = io_imem_resp_bits_data_0 & 32'hffdfffff;
  assign T302 = T303 | T26;
  assign T303 = T306 | T304;
  assign T304 = T305 == 32'h2004033;
  assign T305 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T306 = T309 | T307;
  assign T307 = T308 == 32'h5033;
  assign T308 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T309 = T312 | T310;
  assign T310 = T311 == 32'h501b;
  assign T311 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T312 = T315 | T313;
  assign T313 = T314 == 32'h5013;
  assign T314 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T315 = T318 | T316;
  assign T316 = T317 == 32'h2073;
  assign T317 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T318 = T319 | T29;
  assign T319 = T322 | T320;
  assign T320 = T321 == 32'h2013;
  assign T321 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T322 = T325 | T323;
  assign T323 = T324 == 32'h101b;
  assign T324 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T325 = T328 | T326;
  assign T326 = T327 == 32'h1013;
  assign T327 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T328 = T331 | T329;
  assign T329 = T330 == 32'h73;
  assign T330 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T331 = T334 | T332;
  assign T332 = T333 == 32'h6f;
  assign T333 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T334 = T337 | T335;
  assign T335 = T336 == 32'h63;
  assign T336 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T337 = T340 | T338;
  assign T338 = T339 == 32'h33;
  assign T339 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T340 = T343 | T341;
  assign T341 = T342 == 32'h33;
  assign T342 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T343 = T346 | T344;
  assign T344 = T345 == 32'h17;
  assign T345 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T346 = T349 | T347;
  assign T347 = T348 == 32'h13;
  assign T348 = io_imem_resp_bits_data_0 & 32'h7077;
  assign T349 = T352 | T350;
  assign T350 = T351 == 32'hf;
  assign T351 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T352 = T355 | T353;
  assign T353 = T354 == 32'h3;
  assign T354 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T355 = T37 | T35;
  assign T356 = csr_io_interrupt | io_imem_resp_bits_xcpt_if;
  assign T357 = ctrl_killd ^ 1'h1;
  assign T358 = T359 & io_imem_resp_valid;
  assign T359 = csr_io_interrupt & T360;
  assign T360 = take_pc ^ 1'h1;
  assign T361 = ctrl_killx ^ 1'h1;
  assign T362 = T363 & ex_reg_xcpt_interrupt;
  assign T363 = take_pc ^ 1'h1;
  assign replay_mem = T366 | fpu_kill_mem;
  assign fpu_kill_mem = T364 & io_fpu_nack_mem;
  assign T364 = mem_reg_valid & mem_ctrl_fp;
  assign T365 = T515 ? ex_ctrl_fp : mem_ctrl_fp;
  assign T366 = dcache_kill_mem | mem_reg_replay;
  assign T367 = T368 & replay_ex;
  assign T368 = take_pc ^ 1'h1;
  assign dcache_kill_mem = T369 & io_dmem_replay_next_valid;
  assign T369 = mem_reg_valid & mem_ctrl_wxd;
  assign T370 = ctrl_killm ^ 1'h1;
  assign ctrl_killm = T371 | fpu_kill_mem;
  assign T371 = killm_common | mem_xcpt;
  assign killm_common = T373 | T372;
  assign T372 = mem_reg_valid ^ 1'h1;
  assign T373 = T374 | mem_reg_xcpt;
  assign T374 = dcache_kill_mem | take_pc_wb;
  assign wb_set_sboard = T375 | wb_ctrl_rocc;
  assign T375 = wb_ctrl_div | wb_dcache_miss;
  assign T376 = T516 ? mem_ctrl_div : wb_ctrl_div;
  assign T377 = T515 ? ex_ctrl_div : mem_ctrl_div;
  assign T378 = ll_wen | T79;
  assign T379 = id_ctrl_wxd & T380;
  assign T380 = id_waddr != 5'h0;
  assign T381 = T389 | T382;
  assign T382 = T137 & T383;
  assign T383 = T388 & T384;
  assign T384 = T385 - 1'h1;
  assign T385 = 1'h1 << T386;
  assign T386 = T387 + 5'h1;
  assign T387 = id_raddr_1 - id_raddr_1;
  assign T388 = T62 >> id_raddr_1;
  assign T389 = T149 & T390;
  assign T390 = T395 & T391;
  assign T391 = T392 - 1'h1;
  assign T392 = 1'h1 << T393;
  assign T393 = T394 + 5'h1;
  assign T394 = id_raddr_0 - id_raddr_0;
  assign T395 = T62 >> id_raddr_0;
  assign T396 = T421 | id_wb_hazard;
  assign id_wb_hazard = wb_reg_valid & T397;
  assign T397 = T412 | fp_data_hazard_wb;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T398;
  assign T398 = T401 | T399;
  assign T399 = io_fpu_dec_wen & T400;
  assign T400 = id_waddr == wb_waddr;
  assign T401 = T404 | T402;
  assign T402 = io_fpu_dec_ren3 & T403;
  assign T403 = id_raddr3 == wb_waddr;
  assign id_raddr3 = io_imem_resp_bits_data_0[5'h1f:5'h1b];
  assign T404 = T407 | T405;
  assign T405 = io_fpu_dec_ren2 & T406;
  assign T406 = id_raddr_1 == wb_waddr;
  assign T407 = io_fpu_dec_ren1 & T408;
  assign T408 = id_raddr_0 == wb_waddr;
  assign T409 = T516 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign T410 = T515 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign T411 = T103 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign id_ctrl_wfd = 1'h0;
  assign T412 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_ctrl_wxd & T413;
  assign T413 = T416 | T414;
  assign T414 = T379 & T415;
  assign T415 = id_waddr == wb_waddr;
  assign T416 = T419 | T417;
  assign T417 = T137 & T418;
  assign T418 = id_raddr_1 == wb_waddr;
  assign T419 = T149 & T420;
  assign T420 = id_raddr_0 == wb_waddr;
  assign T421 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = mem_reg_valid & T422;
  assign T422 = T434 | fp_data_hazard_mem;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T423;
  assign T423 = T426 | T424;
  assign T424 = io_fpu_dec_wen & T425;
  assign T425 = id_waddr == mem_waddr;
  assign T426 = T429 | T427;
  assign T427 = io_fpu_dec_ren3 & T428;
  assign T428 = id_raddr3 == mem_waddr;
  assign T429 = T432 | T430;
  assign T430 = io_fpu_dec_ren2 & T431;
  assign T431 = id_raddr_1 == mem_waddr;
  assign T432 = io_fpu_dec_ren1 & T433;
  assign T433 = id_raddr_0 == mem_waddr;
  assign T434 = data_hazard_mem & mem_cannot_bypass;
  assign mem_cannot_bypass = T435 | mem_ctrl_rocc;
  assign T435 = T436 | mem_ctrl_fp;
  assign T436 = T437 | mem_ctrl_div;
  assign T437 = T483 | T438;
  assign T438 = mem_ctrl_mem & mem_mem_cmd_bh;
  assign T439 = T515 ? ex_slow_bypass : mem_mem_cmd_bh;
  assign ex_slow_bypass = T456 | T440;
  assign T440 = T451 | T441;
  assign T441 = 3'h5 == ex_ctrl_mem_type;
  assign T442 = T103 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign id_ctrl_mem_type = T443;
  assign T443 = {T449, T444};
  assign T444 = {T447, T445};
  assign T445 = T446 == 32'h1000;
  assign T446 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T447 = T448 == 32'h2000;
  assign T448 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T449 = T450 == 32'h4000;
  assign T450 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T451 = T453 | T452;
  assign T452 = 3'h1 == ex_ctrl_mem_type;
  assign T453 = T455 | T454;
  assign T454 = 3'h4 == ex_ctrl_mem_type;
  assign T455 = 3'h0 == ex_ctrl_mem_type;
  assign T456 = ex_ctrl_mem_cmd == 5'h7;
  assign T457 = T103 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign id_ctrl_mem_cmd = T458;
  assign T458 = {1'h0, T459};
  assign T459 = {T481, T460};
  assign T460 = {T475, T461};
  assign T461 = {T470, T462};
  assign T462 = T465 | T463;
  assign T463 = T464 == 32'h20000020;
  assign T464 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T465 = T468 | T466;
  assign T466 = T467 == 32'h18000020;
  assign T467 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T468 = T469 == 32'h20;
  assign T469 = io_imem_resp_bits_data_0 & 32'h28;
  assign T470 = T473 | T471;
  assign T471 = T472 == 32'h40000008;
  assign T472 = io_imem_resp_bits_data_0 & 32'h40000008;
  assign T473 = T474 == 32'h10000008;
  assign T474 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T475 = T478 | T476;
  assign T476 = T477 == 32'h80000008;
  assign T477 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T478 = T479 | T473;
  assign T479 = T480 == 32'h8000008;
  assign T480 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T481 = T482 == 32'h8;
  assign T482 = io_imem_resp_bits_data_0 & 32'h18000008;
  assign T483 = mem_ctrl_csr != 3'h0;
  assign T484 = T515 ? ex_ctrl_csr : mem_ctrl_csr;
  assign T485 = T103 ? id_csr : T486;
  assign T486 = T103 ? id_ctrl_csr : ex_ctrl_csr;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_ex_hazard = ex_reg_valid & T487;
  assign T487 = T499 | fp_data_hazard_ex;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T488;
  assign T488 = T491 | T489;
  assign T489 = io_fpu_dec_wen & T490;
  assign T490 = id_waddr == ex_waddr;
  assign ex_waddr = ex_reg_inst[4'hb:3'h7];
  assign T491 = T494 | T492;
  assign T492 = io_fpu_dec_ren3 & T493;
  assign T493 = id_raddr3 == ex_waddr;
  assign T494 = T497 | T495;
  assign T495 = io_fpu_dec_ren2 & T496;
  assign T496 = id_raddr_1 == ex_waddr;
  assign T497 = io_fpu_dec_ren1 & T498;
  assign T498 = id_raddr_0 == ex_waddr;
  assign T499 = data_hazard_ex & ex_cannot_bypass;
  assign ex_cannot_bypass = T500 | ex_ctrl_rocc;
  assign T500 = T501 | ex_ctrl_fp;
  assign T501 = T502 | ex_ctrl_div;
  assign T502 = T503 | ex_ctrl_mem;
  assign T503 = T504 | ex_ctrl_jalr;
  assign T504 = ex_ctrl_csr != 3'h0;
  assign data_hazard_ex = ex_ctrl_wxd & T505;
  assign T505 = T508 | T506;
  assign T506 = T379 & T507;
  assign T507 = id_waddr == ex_waddr;
  assign T508 = T511 | T509;
  assign T509 = T137 & T510;
  assign T510 = id_raddr_1 == ex_waddr;
  assign T511 = T149 & T512;
  assign T512 = id_raddr_0 == ex_waddr;
  assign T513 = T514 | take_pc;
  assign T514 = io_imem_resp_valid ^ 1'h1;
  assign T515 = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T516 = T517 | mem_reg_xcpt_interrupt;
  assign T517 = mem_reg_valid | mem_reg_replay;
  assign T518 = wb_reg_inst;
  assign T519 = R520;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T573 : T522;
  assign T522 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T523 = T562 ? T537 : T524;
  assign T524 = T103 ? T525 : ex_reg_rs_lsb_1;
  assign T525 = T536 ? 2'h0 : T526;
  assign T526 = T533 ? 2'h1 : T527;
  assign T527 = T528 ? 2'h2 : 2'h3;
  assign T528 = T530 & T529;
  assign T529 = mem_waddr == id_raddr_1;
  assign T530 = T532 & T531;
  assign T531 = mem_ctrl_mem ^ 1'h1;
  assign T532 = mem_reg_valid & mem_ctrl_wxd;
  assign T533 = T535 & T534;
  assign T534 = ex_waddr == id_raddr_1;
  assign T535 = ex_reg_valid & ex_ctrl_wxd;
  assign T536 = 5'h0 == id_raddr_1;
  assign T537 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T538;
  assign T538 = T560 ? rf_wdata : T539;
  assign T539 = T540[T548];
  assign T542 = T545 & T543;
  assign T543 = T544 < 5'h1f;
  assign T544 = T547[3'h4:1'h0];
  assign T545 = rf_wen & T546;
  assign T546 = rf_waddr != 5'h0;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign rf_wen = wb_wen | ll_wen;
  assign T547 = ~ rf_waddr;
  assign T548 = ~ T549;
  assign T549 = id_raddr_1[3'h4:1'h0];
  assign rf_wdata = T559 ? io_dmem_resp_bits_data : T550;
  assign T550 = ll_wen ? ll_wdata : T551;
  assign T551 = T557 ? csr_io_rw_rdata : bypass_mux_2;
  assign T552 = T516 ? T553 : bypass_mux_2;
  assign T553 = T556 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = T554;
  assign T554 = mem_ctrl_jalr ? T925 : T555;
  assign T555 = bypass_mux_1;
  assign T925 = {T926, mem_br_target};
  assign T926 = T927 ? 24'hffffff : 24'h0;
  assign T927 = mem_br_target[6'h27:6'h27];
  assign T556 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T557 = wb_ctrl_csr != 3'h0;
  assign T558 = T516 ? mem_ctrl_csr : wb_ctrl_csr;
  assign ll_wdata = div_io_resp_bits_data;
  assign T559 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T560 = T545 & T561;
  assign T561 = rf_waddr == id_raddr_1;
  assign T562 = T103 & T563;
  assign T563 = id_ctrl_rxs2 & T564;
  assign T564 = T565 ^ 1'h1;
  assign T565 = T569 | T566;
  assign T566 = T568 & T567;
  assign T567 = mem_waddr == id_raddr_1;
  assign T568 = mem_reg_valid & mem_ctrl_wxd;
  assign T569 = T570 | T528;
  assign T570 = T536 | T533;
  assign T571 = T562 ? T572 : ex_reg_rs_msb_1;
  assign T572 = id_rs_1 >> 2'h2;
  assign T573 = T579 ? T577 : T574;
  assign T574 = T575 ? bypass_mux_1 : 64'h0;
  assign T575 = T576[1'h0:1'h0];
  assign T576 = ex_reg_rs_lsb_1;
  assign T577 = T578 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T578 = T576[1'h0:1'h0];
  assign T579 = T576[1'h1:1'h1];
  assign T580 = T103 ? T565 : ex_reg_rs_bypass_1;
  assign T581 = T582;
  assign T582 = wb_reg_inst[5'h18:5'h14];
  assign T583 = R584;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T614 : T586;
  assign T586 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T587 = T604 ? T597 : T588;
  assign T588 = T103 ? T589 : ex_reg_rs_lsb_0;
  assign T589 = T596 ? 2'h0 : T590;
  assign T590 = T594 ? 2'h1 : T591;
  assign T591 = T592 ? 2'h2 : 2'h3;
  assign T592 = T530 & T593;
  assign T593 = mem_waddr == id_raddr_0;
  assign T594 = T535 & T595;
  assign T595 = ex_waddr == id_raddr_0;
  assign T596 = 5'h0 == id_raddr_0;
  assign T597 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T598;
  assign T598 = T602 ? rf_wdata : T599;
  assign T599 = T540[T600];
  assign T600 = ~ T601;
  assign T601 = id_raddr_0[3'h4:1'h0];
  assign T602 = T545 & T603;
  assign T603 = rf_waddr == id_raddr_0;
  assign T604 = T103 & T605;
  assign T605 = id_ctrl_rxs1 & T606;
  assign T606 = T607 ^ 1'h1;
  assign T607 = T610 | T608;
  assign T608 = T568 & T609;
  assign T609 = mem_waddr == id_raddr_0;
  assign T610 = T611 | T592;
  assign T611 = T596 | T594;
  assign T612 = T604 ? T613 : ex_reg_rs_msb_0;
  assign T613 = id_rs_0 >> 2'h2;
  assign T614 = T620 ? T618 : T615;
  assign T615 = T616 ? bypass_mux_1 : 64'h0;
  assign T616 = T617[1'h0:1'h0];
  assign T617 = ex_reg_rs_lsb_0;
  assign T618 = T619 ? io_dmem_resp_bits_data_word_bypass : bypass_mux_2;
  assign T619 = T617[1'h0:1'h0];
  assign T620 = T617[1'h1:1'h1];
  assign T621 = T103 ? T607 : ex_reg_rs_bypass_0;
  assign T622 = T623;
  assign T623 = wb_reg_inst[5'h13:4'hf];
  assign T624 = rf_wen;
  assign T625 = rf_wdata;
  assign T626 = T627;
  assign T627 = rf_wen ? rf_waddr : 5'h0;
  assign T628 = wb_reg_pc;
  assign T629 = T516 ? mem_reg_pc : wb_reg_pc;
  assign T630 = wb_valid;
  assign T631 = T632;
  assign T632 = csr_io_time[6'h20:1'h0];
  assign T633 = io_host_id;
  assign T635 = T68 ? 1'h0 : T636;
  assign T636 = T637 ^ 1'h1;
  assign T637 = wb_reg_valid & wb_ctrl_wxd;
  assign T638 = killm_common & R639;
  assign T640 = div_io_req_ready & T691;
  assign T641 = T103 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign id_ctrl_alu_dw = T642;
  assign T642 = T645 | T643;
  assign T643 = T644 == 32'h0;
  assign T644 = io_imem_resp_bits_data_0 & 32'h8;
  assign T645 = T646 == 32'h0;
  assign T646 = io_imem_resp_bits_data_0 & 32'h10;
  assign T647 = T103 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign id_ctrl_alu_fn = T648;
  assign T648 = {T684, T649};
  assign T649 = {T673, T650};
  assign T650 = {T659, T651};
  assign T651 = T654 | T652;
  assign T652 = T653 == 32'h7000;
  assign T653 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T654 = T657 | T655;
  assign T655 = T656 == 32'h1040;
  assign T656 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T657 = T658 == 32'h1010;
  assign T658 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T659 = T662 | T660;
  assign T660 = T661 == 32'h40001010;
  assign T661 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T662 = T665 | T663;
  assign T663 = T664 == 32'h40000030;
  assign T664 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T665 = T668 | T666;
  assign T666 = T667 == 32'h6010;
  assign T667 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T668 = T671 | T669;
  assign T669 = T670 == 32'h3010;
  assign T670 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T671 = T672 == 32'h2040;
  assign T672 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T673 = T676 | T674;
  assign T674 = T675 == 32'h4040;
  assign T675 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T676 = T679 | T677;
  assign T677 = T678 == 32'h4010;
  assign T678 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T679 = T682 | T680;
  assign T680 = T681 == 32'h4010;
  assign T681 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T682 = T683 == 32'h2010;
  assign T683 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T684 = T687 | T685;
  assign T685 = T686 == 32'h40001010;
  assign T686 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T687 = T688 | T663;
  assign T688 = T211 | T689;
  assign T689 = T690 == 32'h2010;
  assign T690 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T691 = ex_reg_valid & ex_ctrl_div;
  assign T692 = ex_op1;
  assign ex_op1 = T707 ? T706 : T928;
  assign T928 = {T929, T693};
  assign T693 = T695 ? T694 : 40'h0;
  assign T694 = ex_reg_pc;
  assign T695 = ex_ctrl_sel_alu1 == 2'h2;
  assign T696 = T103 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign id_ctrl_sel_alu1 = T697;
  assign T697 = {T703, T698};
  assign T698 = T699 | T155;
  assign T699 = T700 | T158;
  assign T700 = T160 | T701;
  assign T701 = T702 == 32'h0;
  assign T702 = io_imem_resp_bits_data_0 & 32'h50;
  assign T703 = T704 | T96;
  assign T704 = T705 == 32'h4;
  assign T705 = io_imem_resp_bits_data_0 & 32'h24;
  assign T929 = T930 ? 24'hffffff : 24'h0;
  assign T930 = T693[6'h27:6'h27];
  assign T706 = ex_rs_0;
  assign T707 = ex_ctrl_sel_alu1 == 2'h1;
  assign T708 = ex_op2;
  assign ex_op2 = T807 ? T806 : T931;
  assign T931 = {T937, T709};
  assign T709 = T805 ? ex_imm : T932;
  assign T932 = {T933, T710};
  assign T710 = T711 ? 4'h4 : 4'h0;
  assign T711 = ex_ctrl_sel_alu2 == 2'h1;
  assign T712 = T103 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign id_ctrl_sel_alu2 = T713;
  assign T713 = {T724, T714};
  assign T714 = T717 | T715;
  assign T715 = T716 == 32'h4050;
  assign T716 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T717 = T718 | T96;
  assign T718 = T719 | T101;
  assign T719 = T722 | T720;
  assign T720 = T721 == 32'h0;
  assign T721 = io_imem_resp_bits_data_0 & 32'h20;
  assign T722 = T723 == 32'h0;
  assign T723 = io_imem_resp_bits_data_0 & 32'h58;
  assign T724 = T727 | T725;
  assign T725 = T726 == 32'h4000;
  assign T726 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T727 = T728 | T155;
  assign T728 = T729 | T158;
  assign T729 = T730 == 32'h0;
  assign T730 = io_imem_resp_bits_data_0 & 32'h48;
  assign T933 = T934 ? 28'hfffffff : 28'h0;
  assign T934 = T710[2'h3:2'h3];
  assign ex_imm = T731;
  assign T731 = {T793, T732};
  assign T732 = {T771, T733};
  assign T733 = {T760, T734};
  assign T734 = T759 ? T758 : T735;
  assign T735 = T757 ? T756 : T736;
  assign T736 = T738 ? T737 : 1'h0;
  assign T737 = ex_reg_inst[4'hf:4'hf];
  assign T738 = ex_ctrl_sel_imm == 3'h5;
  assign T739 = T103 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign id_ctrl_sel_imm = T740;
  assign T740 = {T750, T741};
  assign T741 = {T747, T742};
  assign T742 = T745 | T743;
  assign T743 = T744 == 32'h40;
  assign T744 = io_imem_resp_bits_data_0 & 32'h44;
  assign T745 = T746 == 32'h8;
  assign T746 = io_imem_resp_bits_data_0 & 32'h18;
  assign T747 = T748 | T745;
  assign T748 = T749 == 32'h4;
  assign T749 = io_imem_resp_bits_data_0 & 32'h44;
  assign T750 = T753 | T751;
  assign T751 = T752 == 32'h10;
  assign T752 = io_imem_resp_bits_data_0 & 32'h14;
  assign T753 = T754 | T237;
  assign T754 = T755 == 32'h0;
  assign T755 = io_imem_resp_bits_data_0 & 32'h24;
  assign T756 = ex_reg_inst[5'h14:5'h14];
  assign T757 = ex_ctrl_sel_imm == 3'h4;
  assign T758 = ex_reg_inst[3'h7:3'h7];
  assign T759 = ex_ctrl_sel_imm == 3'h0;
  assign T760 = T770 ? 4'h0 : T761;
  assign T761 = T767 ? T766 : T762;
  assign T762 = T765 ? T764 : T763;
  assign T763 = ex_reg_inst[5'h18:5'h15];
  assign T764 = ex_reg_inst[5'h13:5'h10];
  assign T765 = ex_ctrl_sel_imm == 3'h5;
  assign T766 = ex_reg_inst[4'hb:4'h8];
  assign T767 = T769 | T768;
  assign T768 = ex_ctrl_sel_imm == 3'h1;
  assign T769 = ex_ctrl_sel_imm == 3'h0;
  assign T770 = ex_ctrl_sel_imm == 3'h2;
  assign T771 = {T777, T772};
  assign T772 = T774 ? 6'h0 : T773;
  assign T773 = ex_reg_inst[5'h1e:5'h19];
  assign T774 = T776 | T775;
  assign T775 = ex_ctrl_sel_imm == 3'h5;
  assign T776 = ex_ctrl_sel_imm == 3'h2;
  assign T777 = T790 ? 1'h0 : T778;
  assign T778 = T789 ? T787 : T779;
  assign T779 = T786 ? T784 : T780;
  assign T780 = T783 ? 1'h0 : T781;
  assign T781 = T782;
  assign T782 = ex_reg_inst[5'h1f:5'h1f];
  assign T783 = ex_ctrl_sel_imm == 3'h5;
  assign T784 = T785;
  assign T785 = ex_reg_inst[3'h7:3'h7];
  assign T786 = ex_ctrl_sel_imm == 3'h1;
  assign T787 = T788;
  assign T788 = ex_reg_inst[5'h14:5'h14];
  assign T789 = ex_ctrl_sel_imm == 3'h3;
  assign T790 = T792 | T791;
  assign T791 = ex_ctrl_sel_imm == 3'h5;
  assign T792 = ex_ctrl_sel_imm == 3'h2;
  assign T793 = {T780, T794};
  assign T794 = {T801, T795};
  assign T795 = T798 ? T935 : T796;
  assign T796 = T797;
  assign T797 = ex_reg_inst[5'h13:4'hc];
  assign T935 = T780 ? 8'hff : 8'h0;
  assign T798 = T800 & T799;
  assign T799 = ex_ctrl_sel_imm != 3'h3;
  assign T800 = ex_ctrl_sel_imm != 3'h2;
  assign T801 = T804 ? T802 : T936;
  assign T936 = T780 ? 11'h7ff : 11'h0;
  assign T802 = T803;
  assign T803 = ex_reg_inst[5'h1e:5'h14];
  assign T804 = ex_ctrl_sel_imm == 3'h2;
  assign T805 = ex_ctrl_sel_alu2 == 2'h3;
  assign T937 = T938 ? 32'hffffffff : 32'h0;
  assign T938 = T709[5'h1f:5'h1f];
  assign T806 = ex_rs_1;
  assign T807 = ex_ctrl_sel_alu2 == 2'h2;
  assign T808 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T270 ? mem_reg_cause : T939;
  assign T939 = {61'h0, T809};
  assign T809 = T269 ? 3'h0 : T810;
  assign T810 = T266 ? 3'h6 : T811;
  assign T811 = T263 ? 3'h4 : T812;
  assign T812 = T260 ? 3'h7 : 3'h5;
  assign T813 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T274 ? ex_reg_cause : 64'h2;
  assign T814 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : T940;
  assign T940 = {62'h0, T815};
  assign T815 = io_imem_resp_bits_xcpt_if ? 2'h1 : 2'h2;
  assign T816 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T817 = wb_reg_inst[5'h1f:5'h14];
  assign io_rocc_exception = T818;
  assign T818 = wb_xcpt & T819;
  assign T819 = csr_io_status_xs != 2'h0;
  assign io_rocc_s = T820;
  assign T820 = csr_io_status_prv != 2'h0;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T821 = T827 ? mem_reg_rs2 : wb_reg_rs2;
  assign T822 = T823 ? ex_rs_1 : mem_reg_rs2;
  assign T823 = T515 & T824;
  assign T824 = ex_ctrl_rxs2 & T825;
  assign T825 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T826 = T103 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign T827 = T516 & mem_ctrl_rocc;
  assign io_rocc_cmd_bits_rs1 = bypass_mux_2;
  assign io_rocc_cmd_bits_inst_opcode = T828;
  assign T828 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T829;
  assign T829 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T830;
  assign T830 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T831;
  assign T831 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T832;
  assign T832 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T833;
  assign T833 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T834;
  assign T834 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T835;
  assign T835 = wb_reg_inst[5'h1f:5'h19];
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = T837 & T836;
  assign T836 = replay_wb_common ^ 1'h1;
  assign T837 = wb_reg_valid & wb_ctrl_rocc;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T838;
  assign T838 = T839 & id_ctrl_fp;
  assign T839 = ctrl_killd ^ 1'h1;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T840;
  assign T840 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T841;
  assign T841 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_ptw_status_ie = csr_io_status_ie;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_ie1 = csr_io_status_ie1;
  assign io_ptw_status_prv1 = csr_io_status_prv1;
  assign io_ptw_status_ie2 = csr_io_status_ie2;
  assign io_ptw_status_prv2 = csr_io_status_prv2;
  assign io_ptw_status_ie3 = csr_io_status_ie3;
  assign io_ptw_status_prv3 = csr_io_status_prv3;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_ptbr = csr_io_ptbr;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_dmem_req_bits_data = T842;
  assign T842 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_kill = T843;
  assign T843 = killm_common | mem_xcpt;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_tag = T941;
  assign T941 = {3'h0, T844};
  assign T844 = {ex_waddr, ex_ctrl_fp};
  assign io_dmem_req_bits_addr = T845;
  assign T845 = T846;
  assign T846 = {T848, T847};
  assign T847 = alu_io_adder_out[6'h26:1'h0];
  assign T848 = T861 ? T860 : T849;
  assign T849 = T854 ? T852 : T850;
  assign T850 = T851[1'h0:1'h0];
  assign T851 = alu_io_adder_out[6'h27:6'h26];
  assign T852 = T853 == 2'h3;
  assign T853 = T851;
  assign T854 = T858 | T855;
  assign T855 = T856 == 26'h3fffffe;
  assign T856 = T857;
  assign T857 = ex_rs_0 >> 6'h26;
  assign T858 = T859 == 26'h3ffffff;
  assign T859 = T857;
  assign T860 = T851 != 2'h0;
  assign T861 = T863 | T862;
  assign T862 = T857 == 26'h1;
  assign T863 = T857 == 26'h0;
  assign io_dmem_req_valid = T864;
  assign T864 = ex_reg_valid & ex_ctrl_mem;
  assign io_imem_invalidate = T865;
  assign T865 = wb_reg_valid & wb_ctrl_fence_i;
  assign T866 = T516 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign T867 = T515 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign T868 = T103 ? id_ctrl_fence_i : ex_ctrl_fence_i;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_returnAddr = T942;
  assign T942 = mem_int_wdata[6'h26:1'h0];
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_isCall = T869;
  assign T869 = mem_ctrl_wxd & T870;
  assign T870 = mem_waddr[1'h0:1'h0];
  assign io_imem_ras_update_valid = T871;
  assign T871 = T873 & T872;
  assign T872 = take_pc_wb ^ 1'h1;
  assign T873 = T875 & T874;
  assign T874 = mem_npc_misaligned ^ 1'h1;
  assign T875 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_pc = T943;
  assign T943 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_valid = T876;
  assign T876 = T878 & T877;
  assign T877 = take_pc_wb ^ 1'h1;
  assign T878 = mem_reg_valid & mem_ctrl_branch;
  assign io_imem_btb_update_bits_br_pc = T944;
  assign T944 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_isReturn = T879;
  assign T879 = mem_ctrl_jalr & T880;
  assign T880 = 5'h1 == T881;
  assign T881 = T882 & 5'h19;
  assign T882 = mem_reg_inst[5'h13:4'hf];
  assign io_imem_btb_update_bits_isJump = T883;
  assign T883 = mem_ctrl_jal | mem_ctrl_jalr;
  assign io_imem_btb_update_bits_target = T945;
  assign T945 = io_imem_req_bits_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_pc = T946;
  assign T946 = mem_reg_pc[6'h26:1'h0];
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T884 = T887 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T885 = T886 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T886 = T103 & io_imem_btb_resp_valid;
  assign T887 = T515 & ex_reg_btb_hit;
  assign T888 = T103 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign T889 = T887 ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign T890 = T886 ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T891 = T887 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T892 = T886 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T893 = T887 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T894 = T886 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign T895 = T887 ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign T896 = T886 ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign T897 = T887 ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign T898 = T886 ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T899 = T887 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T900 = T886 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T901 = T515 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T902;
  assign T902 = T904 & T903;
  assign T903 = take_pc_wb ^ 1'h1;
  assign T904 = T908 & T905;
  assign T905 = T906 | mem_ctrl_jal;
  assign T906 = T907 | mem_ctrl_jalr;
  assign T907 = mem_ctrl_branch & mem_br_taken;
  assign T908 = T909 & mem_wrong_npc;
  assign T909 = mem_reg_valid & T910;
  assign T910 = mem_npc_misaligned ^ 1'h1;
  assign io_imem_resp_ready = T911;
  assign T911 = T912 | csr_io_interrupt;
  assign T912 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_bits_pc = T913;
  assign T913 = T914;
  assign T914 = T916 ? csr_io_evec : T915;
  assign T915 = replay_wb ? wb_reg_pc : mem_npc;
  assign T916 = wb_xcpt | csr_io_eret;
  assign io_imem_req_valid = take_pc;
  assign io_host_debug_stats_csr = csr_io_host_debug_stats_csr;
  assign io_host_csr_resp_bits = csr_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = csr_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = csr_io_host_csr_req_ready;
  CSRFile csr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( csr_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( csr_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( csr_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( csr_io_host_debug_stats_csr ),
       .io_rw_addr( T817 ),
       .io_rw_cmd( T816 ),
       .io_rw_rdata( csr_io_rw_rdata ),
       .io_rw_wdata( bypass_mux_2 ),
       .io_csr_stall( csr_io_csr_stall ),
       .io_csr_xcpt( csr_io_csr_xcpt ),
       .io_eret( csr_io_eret ),
       .io_status_sd( csr_io_status_sd ),
       .io_status_zero2( csr_io_status_zero2 ),
       .io_status_sd_rv32( csr_io_status_sd_rv32 ),
       .io_status_zero1( csr_io_status_zero1 ),
       .io_status_vm( csr_io_status_vm ),
       .io_status_mprv( csr_io_status_mprv ),
       .io_status_xs( csr_io_status_xs ),
       .io_status_fs( csr_io_status_fs ),
       .io_status_prv3( csr_io_status_prv3 ),
       .io_status_ie3( csr_io_status_ie3 ),
       .io_status_prv2( csr_io_status_prv2 ),
       .io_status_ie2( csr_io_status_ie2 ),
       .io_status_prv1( csr_io_status_prv1 ),
       .io_status_ie1( csr_io_status_ie1 ),
       .io_status_prv( csr_io_status_prv ),
       .io_status_ie( csr_io_status_ie ),
       .io_ptbr( csr_io_ptbr ),
       .io_evec( csr_io_evec ),
       .io_exception( wb_reg_xcpt ),
       .io_retire( wb_valid ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( wb_reg_cause ),
       .io_pc( wb_reg_pc ),
       .io_fatc( csr_io_fatc ),
       .io_time( csr_io_time ),
       .io_fcsr_rm( csr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_invalidate_lr( io_rocc_mem_invalidate_lr ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_autl_acquire_ready(  )
       .io_rocc_autl_acquire_valid( io_rocc_autl_acquire_valid ),
       .io_rocc_autl_acquire_bits_addr_block( io_rocc_autl_acquire_bits_addr_block ),
       .io_rocc_autl_acquire_bits_client_xact_id( io_rocc_autl_acquire_bits_client_xact_id ),
       .io_rocc_autl_acquire_bits_addr_beat( io_rocc_autl_acquire_bits_addr_beat ),
       .io_rocc_autl_acquire_bits_is_builtin_type( io_rocc_autl_acquire_bits_is_builtin_type ),
       .io_rocc_autl_acquire_bits_a_type( io_rocc_autl_acquire_bits_a_type ),
       .io_rocc_autl_acquire_bits_union( io_rocc_autl_acquire_bits_union ),
       .io_rocc_autl_acquire_bits_data( io_rocc_autl_acquire_bits_data ),
       .io_rocc_autl_grant_ready( io_rocc_autl_grant_ready ),
       //.io_rocc_autl_grant_valid(  )
       //.io_rocc_autl_grant_bits_addr_beat(  )
       //.io_rocc_autl_grant_bits_client_xact_id(  )
       //.io_rocc_autl_grant_bits_manager_xact_id(  )
       //.io_rocc_autl_grant_bits_is_builtin_type(  )
       //.io_rocc_autl_grant_bits_g_type(  )
       //.io_rocc_autl_grant_bits_data(  )
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits_addr( io_rocc_iptw_req_bits_addr ),
       .io_rocc_iptw_req_bits_prv( io_rocc_iptw_req_bits_prv ),
       .io_rocc_iptw_req_bits_store( io_rocc_iptw_req_bits_store ),
       .io_rocc_iptw_req_bits_fetch( io_rocc_iptw_req_bits_fetch ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits_addr( io_rocc_dptw_req_bits_addr ),
       .io_rocc_dptw_req_bits_prv( io_rocc_dptw_req_bits_prv ),
       .io_rocc_dptw_req_bits_store( io_rocc_dptw_req_bits_store ),
       .io_rocc_dptw_req_bits_fetch( io_rocc_dptw_req_bits_fetch ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits_addr( io_rocc_pptw_req_bits_addr ),
       .io_rocc_pptw_req_bits_prv( io_rocc_pptw_req_bits_prv ),
       .io_rocc_pptw_req_bits_store( io_rocc_pptw_req_bits_store ),
       .io_rocc_pptw_req_bits_fetch( io_rocc_pptw_req_bits_fetch ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_fpu_req_ready(  )
       .io_rocc_fpu_req_valid( io_rocc_fpu_req_valid ),
       .io_rocc_fpu_req_bits_cmd( io_rocc_fpu_req_bits_cmd ),
       .io_rocc_fpu_req_bits_ldst( io_rocc_fpu_req_bits_ldst ),
       .io_rocc_fpu_req_bits_wen( io_rocc_fpu_req_bits_wen ),
       .io_rocc_fpu_req_bits_ren1( io_rocc_fpu_req_bits_ren1 ),
       .io_rocc_fpu_req_bits_ren2( io_rocc_fpu_req_bits_ren2 ),
       .io_rocc_fpu_req_bits_ren3( io_rocc_fpu_req_bits_ren3 ),
       .io_rocc_fpu_req_bits_swap12( io_rocc_fpu_req_bits_swap12 ),
       .io_rocc_fpu_req_bits_swap23( io_rocc_fpu_req_bits_swap23 ),
       .io_rocc_fpu_req_bits_single( io_rocc_fpu_req_bits_single ),
       .io_rocc_fpu_req_bits_fromint( io_rocc_fpu_req_bits_fromint ),
       .io_rocc_fpu_req_bits_toint( io_rocc_fpu_req_bits_toint ),
       .io_rocc_fpu_req_bits_fastpipe( io_rocc_fpu_req_bits_fastpipe ),
       .io_rocc_fpu_req_bits_fma( io_rocc_fpu_req_bits_fma ),
       .io_rocc_fpu_req_bits_div( io_rocc_fpu_req_bits_div ),
       .io_rocc_fpu_req_bits_sqrt( io_rocc_fpu_req_bits_sqrt ),
       .io_rocc_fpu_req_bits_round( io_rocc_fpu_req_bits_round ),
       .io_rocc_fpu_req_bits_wflags( io_rocc_fpu_req_bits_wflags ),
       .io_rocc_fpu_req_bits_rm( io_rocc_fpu_req_bits_rm ),
       .io_rocc_fpu_req_bits_typ( io_rocc_fpu_req_bits_typ ),
       .io_rocc_fpu_req_bits_in1( io_rocc_fpu_req_bits_in1 ),
       .io_rocc_fpu_req_bits_in2( io_rocc_fpu_req_bits_in2 ),
       .io_rocc_fpu_req_bits_in3( io_rocc_fpu_req_bits_in3 ),
       .io_rocc_fpu_resp_ready( io_rocc_fpu_resp_ready ),
       //.io_rocc_fpu_resp_valid(  )
       //.io_rocc_fpu_resp_bits_data(  )
       //.io_rocc_fpu_resp_bits_exc(  )
       //.io_rocc_exception(  )
       //.io_rocc_dma_req_ready(  )
       .io_rocc_dma_req_valid( io_rocc_dma_req_valid ),
       .io_rocc_dma_req_bits_client_xact_id( io_rocc_dma_req_bits_client_xact_id ),
       .io_rocc_dma_req_bits_cmd( io_rocc_dma_req_bits_cmd ),
       .io_rocc_dma_req_bits_source( io_rocc_dma_req_bits_source ),
       .io_rocc_dma_req_bits_dest( io_rocc_dma_req_bits_dest ),
       .io_rocc_dma_req_bits_length( io_rocc_dma_req_bits_length ),
       .io_rocc_dma_resp_ready( io_rocc_dma_resp_ready ),
       //.io_rocc_dma_resp_valid(  )
       //.io_rocc_dma_resp_bits_client_xact_id(  )
       //.io_rocc_dma_resp_bits_status(  )
       .io_interrupt( csr_io_interrupt ),
       .io_interrupt_cause( csr_io_interrupt_cause )
  );
  ALU alu(
       .io_dw( ex_ctrl_alu_dw ),
       .io_fn( ex_ctrl_alu_fn ),
       .io_in2( T708 ),
       .io_in1( T692 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( T691 ),
       .io_req_bits_fn( ex_ctrl_alu_fn ),
       .io_req_bits_dw( ex_ctrl_alu_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( ex_waddr ),
       .io_kill( T638 ),
       .io_resp_ready( T635 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );

  always @(posedge clk) begin
    if(T516) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T515) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data_0;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T39;
    end
    if(reset) begin
      R73 <= 32'h0;
    end else if(T378) begin
      R73 <= T76;
    end else if(ll_wen) begin
      R73 <= T62;
    end
    if(T516) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if(T515) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if(T103) begin
      ex_ctrl_wxd <= id_ctrl_wxd;
    end
    if(T516) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if(T515) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if(T103) begin
      ex_ctrl_rocc <= id_ctrl_rocc;
    end
    wb_reg_replay <= T113;
    wb_reg_xcpt <= T117;
    if(T515) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_mem <= id_ctrl_mem;
    end
    mem_reg_valid <= T123;
    ex_reg_valid <= T125;
    if(T103) begin
      ex_reg_load_use <= id_load_use;
    end
    if(T516) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if(T103) begin
      ex_ctrl_div <= id_ctrl_div;
    end
    if(T515) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if(T103) begin
      ex_ctrl_jal <= id_ctrl_jal;
    end
    if(T515) begin
      bypass_mux_1 <= alu_io_out;
    end
    if(T515) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if(T103) begin
      ex_ctrl_branch <= id_ctrl_branch;
    end
    if(T515) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T515) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if(T103) begin
      ex_ctrl_jalr <= id_ctrl_jalr;
    end
    if(T515) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if(T103) begin
      ex_reg_flush_pipe <= T242;
    end
    mem_reg_xcpt <= T271;
    if(T103) begin
      ex_ctrl_fp <= id_ctrl_fp;
    end
    ex_reg_xcpt <= T275;
    ex_reg_xcpt_interrupt <= T358;
    mem_reg_xcpt_interrupt <= T362;
    if(T515) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    mem_reg_replay <= T367;
    wb_reg_valid <= T370;
    if(T516) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if(T515) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if(T516) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if(T515) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if(T103) begin
      ex_ctrl_wfd <= id_ctrl_wfd;
    end
    if(T515) begin
      mem_mem_cmd_bh <= ex_slow_bypass;
    end
    if(T103) begin
      ex_ctrl_mem_type <= id_ctrl_mem_type;
    end
    if(T103) begin
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
    end
    if(T515) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if(T103) begin
      ex_ctrl_csr <= id_csr;
    end else if(T103) begin
      ex_ctrl_csr <= id_ctrl_csr;
    end
    R520 <= R521;
    if(ex_reg_rs_bypass_1) begin
      R521 <= T573;
    end else begin
      R521 <= T522;
    end
    if(T562) begin
      ex_reg_rs_lsb_1 <= T537;
    end else if(T103) begin
      ex_reg_rs_lsb_1 <= T525;
    end
    if (T542)
      T540[T547] <= rf_wdata;
    if(T516) begin
      bypass_mux_2 <= T553;
    end
    if(T516) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if(T562) begin
      ex_reg_rs_msb_1 <= T572;
    end
    if(T103) begin
      ex_reg_rs_bypass_1 <= T565;
    end
    R584 <= R585;
    if(ex_reg_rs_bypass_0) begin
      R585 <= T614;
    end else begin
      R585 <= T586;
    end
    if(T604) begin
      ex_reg_rs_lsb_0 <= T597;
    end else if(T103) begin
      ex_reg_rs_lsb_0 <= T589;
    end
    if(T604) begin
      ex_reg_rs_msb_0 <= T613;
    end
    if(T103) begin
      ex_reg_rs_bypass_0 <= T607;
    end
    if(T516) begin
      wb_reg_pc <= mem_reg_pc;
    end
    R639 <= T640;
    if(T103) begin
      ex_ctrl_alu_dw <= id_ctrl_alu_dw;
    end
    if(T103) begin
      ex_ctrl_alu_fn <= id_ctrl_alu_fn;
    end
    if(T103) begin
      ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
    end
    if(T103) begin
      ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
    end
    if(T103) begin
      ex_ctrl_sel_imm <= id_ctrl_sel_imm;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(T827) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(T823) begin
      mem_reg_rs2 <= ex_rs_1;
    end
    if(T103) begin
      ex_ctrl_rxs2 <= id_ctrl_rxs2;
    end
    if(T516) begin
      wb_ctrl_fence_i <= mem_ctrl_fence_i;
    end
    if(T515) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if(T103) begin
      ex_ctrl_fence_i <= id_ctrl_fence_i;
    end
    if(T887) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T886) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(T103) begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T887) begin
      mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
    end
    if(T886) begin
      ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
    end
    if(T887) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T886) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T887) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T886) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T887) begin
      mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
    end
    if(T886) begin
      ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
    end
    if(T887) begin
      mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
    end
    if(T886) begin
      ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
    end
    if(T887) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T886) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T515) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
`ifndef SYNTHESIS
// synthesis translate_off
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T633, T631, T630, T628, T626, T625, T624, T622, T583, T581, T519, T518, T1);
// synthesis translate_on
`endif
  end
endmodule

module BTB(input clk, input reset,
    input  io_req_valid,
    input [38:0] io_req_bits_addr,
    output io_resp_valid,
    output io_resp_bits_taken,
    output io_resp_bits_mask,
    output io_resp_bits_bridx,
    output[38:0] io_resp_bits_target,
    output[2:0] io_resp_bits_entry,
    output[3:0] io_resp_bits_bht_history,
    output[1:0] io_resp_bits_bht_value,
    input  io_btb_update_valid,
    input  io_btb_update_bits_prediction_valid,
    input  io_btb_update_bits_prediction_bits_taken,
    input  io_btb_update_bits_prediction_bits_mask,
    input  io_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_btb_update_bits_prediction_bits_target,
    input [2:0] io_btb_update_bits_prediction_bits_entry,
    input [3:0] io_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_btb_update_bits_pc,
    input [38:0] io_btb_update_bits_target,
    input  io_btb_update_bits_taken,
    input  io_btb_update_bits_isJump,
    input  io_btb_update_bits_isReturn,
    input [38:0] io_btb_update_bits_br_pc,
    input  io_bht_update_valid,
    input  io_bht_update_bits_prediction_valid,
    input  io_bht_update_bits_prediction_bits_taken,
    input  io_bht_update_bits_prediction_bits_mask,
    input  io_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_bht_update_bits_prediction_bits_target,
    input [2:0] io_bht_update_bits_prediction_bits_entry,
    input [3:0] io_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_bht_update_bits_pc,
    input  io_bht_update_bits_taken,
    input  io_bht_update_bits_mispredict,
    input  io_ras_update_valid,
    input  io_ras_update_bits_isCall,
    input  io_ras_update_bits_isReturn,
    input [38:0] io_ras_update_bits_returnAddr,
    input  io_ras_update_bits_prediction_valid,
    input  io_ras_update_bits_prediction_bits_taken,
    input  io_ras_update_bits_prediction_bits_mask,
    input  io_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_ras_update_bits_prediction_bits_target,
    input [2:0] io_ras_update_bits_prediction_bits_entry,
    input [3:0] io_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_ras_update_bits_prediction_bits_bht_value,
    input  io_invalidate
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg [38:0] R4;
  wire[38:0] T5;
  wire T6;
  reg  R7;
  wire T464;
  wire[1:0] T8;
  wire[1:0] T9;
  reg [1:0] T10 [15:0];
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire[3:0] T24;
  reg [3:0] R25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[2:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg  isJump_7;
  wire T35;
  reg  R36;
  wire T37;
  wire T38;
  wire T39;
  wire[7:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  reg [2:0] nextRepl;
  wire[2:0] T465;
  wire[2:0] T43;
  wire[2:0] T44;
  wire T45;
  wire T46;
  reg [2:0] R47;
  wire[2:0] T48;
  reg  updateHit;
  wire T49;
  wire T50;
  wire[7:0] hits;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[3:0] T53;
  wire[1:0] T54;
  wire T55;
  wire[3:0] T56;
  wire[3:0] pageHit;
  reg [3:0] pageValid;
  wire[3:0] T466;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[3:0] pageReplEn;
  wire[3:0] tgtPageReplEn;
  wire[3:0] tgtPageRepl;
  wire[3:0] T60;
  wire[3:0] T467;
  wire T61;
  wire[3:0] T62;
  wire[2:0] T63;
  wire[3:0] idxPageUpdateOH;
  wire[3:0] idxPageRepl;
  wire[3:0] T64;
  reg [1:0] R65;
  wire[1:0] T468;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire doPageRepl;
  wire doIdxPageRepl;
  wire[3:0] updatePageHit;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[1:0] T71;
  wire T72;
  wire[26:0] T73;
  reg [38:0] R74;
  wire[38:0] T75;
  wire[26:0] T76;
  reg [26:0] pages [3:0];
  wire[26:0] T77;
  wire[26:0] T78;
  wire[26:0] T79;
  wire[26:0] T80;
  wire T81;
  wire[3:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[26:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[26:0] T91;
  wire[26:0] T92;
  wire[26:0] T93;
  wire[26:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[26:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire[26:0] T104;
  wire[1:0] T105;
  wire T106;
  wire[26:0] T107;
  wire T108;
  wire[26:0] T109;
  wire useUpdatePageHit;
  wire samePage;
  wire[26:0] T110;
  wire[26:0] T111;
  wire doTgtPageRepl;
  wire T112;
  wire usePageHit;
  wire[3:0] T113;
  wire[3:0] T114;
  wire T115;
  wire[3:0] idxPageReplEn;
  wire T116;
  wire[3:0] T117;
  wire[3:0] T118;
  wire[1:0] T119;
  wire T120;
  wire[26:0] T121;
  wire[26:0] T122;
  wire T123;
  wire[26:0] T124;
  wire[1:0] T125;
  wire T126;
  wire[26:0] T127;
  wire T128;
  wire[26:0] T129;
  wire[3:0] idxPagesOH_0;
  wire[3:0] T130;
  wire[1:0] T131;
  reg [1:0] idxPages [7:0];
  wire[1:0] T132;
  wire[1:0] T469;
  wire T470;
  wire[1:0] T471;
  wire[1:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T133;
  wire[3:0] T134;
  wire[3:0] idxPagesOH_1;
  wire[3:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire[3:0] T139;
  wire[3:0] idxPagesOH_2;
  wire[3:0] T140;
  wire[1:0] T141;
  wire T142;
  wire[3:0] T143;
  wire[3:0] idxPagesOH_3;
  wire[3:0] T144;
  wire[1:0] T145;
  wire[3:0] T146;
  wire[1:0] T147;
  wire T148;
  wire[3:0] T149;
  wire[3:0] idxPagesOH_4;
  wire[3:0] T150;
  wire[1:0] T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] idxPagesOH_5;
  wire[3:0] T154;
  wire[1:0] T155;
  wire[1:0] T156;
  wire T157;
  wire[3:0] T158;
  wire[3:0] idxPagesOH_6;
  wire[3:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[3:0] T162;
  wire[3:0] idxPagesOH_7;
  wire[3:0] T163;
  wire[1:0] T164;
  wire[7:0] T165;
  wire[7:0] T166;
  wire[7:0] T167;
  wire[3:0] T168;
  wire[1:0] T169;
  wire T170;
  wire[11:0] T171;
  wire[11:0] T172;
  reg [11:0] idxs [7:0];
  wire[11:0] T173;
  wire[11:0] T475;
  wire T174;
  wire[11:0] T175;
  wire[1:0] T176;
  wire T177;
  wire[11:0] T178;
  wire T179;
  wire[11:0] T180;
  wire[3:0] T181;
  wire[1:0] T182;
  wire T183;
  wire[11:0] T184;
  wire T185;
  wire[11:0] T186;
  wire[1:0] T187;
  wire T188;
  wire[11:0] T189;
  wire T190;
  wire[11:0] T191;
  reg [7:0] idxValid;
  wire[7:0] T476;
  wire[7:0] T192;
  wire[7:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[7:0] T196;
  wire[7:0] T197;
  wire[7:0] T198;
  wire[7:0] T199;
  wire[3:0] T200;
  wire[1:0] T201;
  wire T202;
  wire[3:0] T203;
  wire[3:0] T204;
  wire[3:0] tgtPagesOH_0;
  wire[3:0] T205;
  wire[1:0] T206;
  reg [1:0] tgtPages [7:0];
  wire[1:0] T207;
  wire[1:0] T477;
  wire T478;
  wire[1:0] T479;
  wire[1:0] T480;
  wire[3:0] T208;
  wire[1:0] T481;
  wire T482;
  wire T209;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[3:0] tgtPagesOH_1;
  wire[3:0] T212;
  wire[1:0] T213;
  wire[1:0] T214;
  wire T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] tgtPagesOH_2;
  wire[3:0] T218;
  wire[1:0] T219;
  wire T220;
  wire[3:0] T221;
  wire[3:0] T222;
  wire[3:0] tgtPagesOH_3;
  wire[3:0] T223;
  wire[1:0] T224;
  wire[3:0] T225;
  wire[1:0] T226;
  wire T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[3:0] tgtPagesOH_4;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] tgtPagesOH_5;
  wire[3:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire T238;
  wire[3:0] T239;
  wire[3:0] T240;
  wire[3:0] tgtPagesOH_6;
  wire[3:0] T241;
  wire[1:0] T242;
  wire T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[3:0] tgtPagesOH_7;
  wire[3:0] T246;
  wire[1:0] T247;
  wire T248;
  wire T249;
  reg  isJump_6;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  reg  isJump_5;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  reg  isJump_4;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  reg  isJump_3;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  reg  isJump_2;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  reg  isJump_1;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  reg  isJump_0;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire[3:0] T290;
  wire[2:0] T291;
  wire T292;
  wire[3:0] T293;
  wire[3:0] T294;
  wire[2:0] T483;
  wire[1:0] T484;
  wire T485;
  wire[1:0] T486;
  wire[1:0] T487;
  wire[3:0] T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[1:0] T491;
  wire T492;
  wire T493;
  wire[38:0] T296;
  wire[38:0] T297;
  wire[38:0] T298;
  wire[11:0] T299;
  wire[11:0] T300;
  wire[11:0] T301;
  reg [11:0] tgts [7:0];
  wire[11:0] T302;
  wire[11:0] T494;
  wire T303;
  wire[11:0] T304;
  wire[11:0] T305;
  wire[11:0] T306;
  wire T307;
  wire[11:0] T308;
  wire[11:0] T309;
  wire[11:0] T310;
  wire T311;
  wire[11:0] T312;
  wire[11:0] T313;
  wire[11:0] T314;
  wire T315;
  wire[11:0] T316;
  wire[11:0] T317;
  wire[11:0] T318;
  wire T319;
  wire[11:0] T320;
  wire[11:0] T321;
  wire[11:0] T322;
  wire T323;
  wire[11:0] T324;
  wire[11:0] T325;
  wire[11:0] T326;
  wire T327;
  wire[11:0] T328;
  wire[11:0] T329;
  wire T330;
  wire[26:0] T331;
  wire[26:0] T332;
  wire[26:0] T333;
  wire T334;
  wire[3:0] T335;
  wire[3:0] T336;
  wire T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire T340;
  wire[3:0] T341;
  wire[3:0] T342;
  wire T343;
  wire[3:0] T344;
  wire[3:0] T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire T349;
  wire[3:0] T350;
  wire[3:0] T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire T355;
  wire[3:0] T356;
  wire T357;
  wire[26:0] T358;
  wire[26:0] T359;
  wire[26:0] T360;
  wire T361;
  wire[26:0] T362;
  wire[26:0] T363;
  wire[26:0] T364;
  wire T365;
  wire[26:0] T366;
  wire[26:0] T367;
  wire T368;
  wire[38:0] T369;
  reg [38:0] R370;
  wire[38:0] T371;
  wire T372;
  wire T373;
  wire[1:0] T374;
  wire T375;
  wire T376;
  reg  R377;
  wire T495;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  reg [1:0] R384;
  wire[1:0] T496;
  wire[1:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire T389;
  wire T390;
  wire[1:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  reg [38:0] R397;
  wire[38:0] T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  reg  useRAS_7;
  wire T405;
  reg  R406;
  wire T407;
  wire T408;
  wire T409;
  wire[7:0] T410;
  wire[2:0] T411;
  wire T412;
  wire T413;
  wire T414;
  reg  useRAS_6;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  reg  useRAS_5;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  reg  useRAS_4;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg  useRAS_3;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  reg  useRAS_2;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg  useRAS_1;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  reg  useRAS_0;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  reg [0:0] brIdx [7:0];
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {2{$random}};
    R7 = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      T10[initvar] = {1{$random}};
    R25 = {1{$random}};
    isJump_7 = {1{$random}};
    R36 = {1{$random}};
    nextRepl = {1{$random}};
    R47 = {1{$random}};
    updateHit = {1{$random}};
    pageValid = {1{$random}};
    R65 = {1{$random}};
    R74 = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    isJump_6 = {1{$random}};
    isJump_5 = {1{$random}};
    isJump_4 = {1{$random}};
    isJump_3 = {1{$random}};
    isJump_2 = {1{$random}};
    isJump_1 = {1{$random}};
    isJump_0 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R370 = {2{$random}};
    R377 = {1{$random}};
    R384 = {1{$random}};
    R397 = {2{$random}};
    useRAS_7 = {1{$random}};
    R406 = {1{$random}};
    useRAS_6 = {1{$random}};
    useRAS_5 = {1{$random}};
    useRAS_4 = {1{$random}};
    useRAS_3 = {1{$random}};
    useRAS_2 = {1{$random}};
    useRAS_1 = {1{$random}};
    useRAS_0 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      brIdx[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req_bits_addr == R4;
  assign T5 = io_btb_update_valid ? io_btb_update_bits_target : R4;
  assign T6 = R7 ^ 1'h1;
  assign T464 = reset ? 1'h0 : io_btb_update_valid;
  assign io_resp_bits_bht_value = T8;
  assign T8 = T9;
  assign T9 = T10[T24];
  assign T12 = {io_bht_update_bits_taken, T13};
  assign T13 = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = T17 | T16;
  assign T16 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T17 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T18 = T20 & T19;
  assign T19 = io_bht_update_bits_prediction_bits_bht_value[1'h0:1'h0];
  assign T20 = io_bht_update_bits_prediction_bits_bht_value[1'h1:1'h1];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22 = T23 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T23 = io_bht_update_bits_pc[3'h5:2'h2];
  assign T24 = T293 ^ R25;
  assign T26 = T292 ? T290 : T27;
  assign T27 = T31 ? T28 : R25;
  assign T28 = {T30, T29};
  assign T29 = R25[2'h3:1'h1];
  assign T30 = T8[1'h0:1'h0];
  assign T31 = T289 & T32;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T248 | T34;
  assign T34 = T50 ? isJump_7 : 1'h0;
  assign T35 = T38 ? R36 : isJump_7;
  assign T37 = io_btb_update_valid ? io_btb_update_bits_isJump : R36;
  assign T38 = R7 & T39;
  assign T39 = T40[3'h7:3'h7];
  assign T40 = 1'h1 << T41;
  assign T41 = T42;
  assign T42 = updateHit ? R47 : nextRepl;
  assign T465 = reset ? 3'h0 : T43;
  assign T43 = T45 ? T44 : nextRepl;
  assign T44 = nextRepl + 3'h1;
  assign T45 = R7 & T46;
  assign T46 = updateHit ^ 1'h1;
  assign T48 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : R47;
  assign T49 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : updateHit;
  assign T50 = hits[3'h7:3'h7];
  assign hits = T165 & T51;
  assign T51 = T52;
  assign T52 = {T146, T53};
  assign T53 = {T137, T54};
  assign T54 = {T133, T55};
  assign T55 = T56 != 4'h0;
  assign T56 = idxPagesOH_0 & pageHit;
  assign pageHit = T117 & pageValid;
  assign T466 = reset ? 4'h0 : T57;
  assign T57 = io_invalidate ? 4'h0 : T58;
  assign T58 = T116 ? T59 : pageValid;
  assign T59 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 4'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T60;
  assign T60 = T62 | T467;
  assign T467 = {3'h0, T61};
  assign T61 = idxPageUpdateOH[2'h3:2'h3];
  assign T62 = T63 << 1'h1;
  assign T63 = idxPageUpdateOH[2'h2:1'h0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T64;
  assign T64 = 1'h1 << R65;
  assign T468 = reset ? 2'h0 : T66;
  assign T66 = T68 ? T67 : R65;
  assign T67 = R65 + 2'h1;
  assign T68 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = useUpdatePageHit ^ 1'h1;
  assign updatePageHit = T69 & pageValid;
  assign T69 = T70;
  assign T70 = {T105, T71};
  assign T71 = {T103, T72};
  assign T72 = T76 == T73;
  assign T73 = R74 >> 4'hc;
  assign T75 = io_btb_update_valid ? io_btb_update_bits_pc : R74;
  assign T76 = pages[2'h0];
  assign T78 = T81 ? T80 : T79;
  assign T79 = R74 >> 4'hc;
  assign T80 = io_req_bits_addr >> 4'hc;
  assign T81 = T82 != 4'h0;
  assign T82 = idxPageUpdateOH & 4'h5;
  assign T83 = R7 & T84;
  assign T84 = T86 & T85;
  assign T85 = pageReplEn[2'h3:2'h3];
  assign T86 = T81 ? doTgtPageRepl : doIdxPageRepl;
  assign T88 = R7 & T89;
  assign T89 = T86 & T90;
  assign T90 = pageReplEn[1'h1:1'h1];
  assign T92 = T81 ? T94 : T93;
  assign T93 = io_req_bits_addr >> 4'hc;
  assign T94 = R74 >> 4'hc;
  assign T95 = R7 & T96;
  assign T96 = T98 & T97;
  assign T97 = pageReplEn[2'h2:2'h2];
  assign T98 = T81 ? doIdxPageRepl : doTgtPageRepl;
  assign T100 = R7 & T101;
  assign T101 = T98 & T102;
  assign T102 = pageReplEn[1'h0:1'h0];
  assign T103 = T104 == T73;
  assign T104 = pages[2'h1];
  assign T105 = {T108, T106};
  assign T106 = T107 == T73;
  assign T107 = pages[2'h2];
  assign T108 = T109 == T73;
  assign T109 = pages[2'h3];
  assign useUpdatePageHit = updatePageHit != 4'h0;
  assign samePage = T111 == T110;
  assign T110 = io_req_bits_addr >> 4'hc;
  assign T111 = R74 >> 4'hc;
  assign doTgtPageRepl = T115 & T112;
  assign T112 = usePageHit ^ 1'h1;
  assign usePageHit = T113 != 4'h0;
  assign T113 = pageHit & T114;
  assign T114 = ~ idxPageReplEn;
  assign T115 = samePage ^ 1'h1;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 4'h0;
  assign T116 = R7 & doPageRepl;
  assign T117 = T118;
  assign T118 = {T125, T119};
  assign T119 = {T123, T120};
  assign T120 = T122 == T121;
  assign T121 = io_req_bits_addr >> 4'hc;
  assign T122 = pages[2'h0];
  assign T123 = T124 == T121;
  assign T124 = pages[2'h1];
  assign T125 = {T128, T126};
  assign T126 = T127 == T121;
  assign T127 = pages[2'h2];
  assign T128 = T129 == T121;
  assign T129 = pages[2'h3];
  assign idxPagesOH_0 = T130[2'h3:1'h0];
  assign T130 = 1'h1 << T131;
  assign T131 = idxPages[3'h0];
  assign T469 = {T474, T470};
  assign T470 = T471[1'h1:1'h1];
  assign T471 = T473 | T472;
  assign T472 = idxPageUpdateOH[1'h1:1'h0];
  assign T473 = idxPageUpdateOH[2'h3:2'h2];
  assign T474 = T473 != 2'h0;
  assign T133 = T134 != 4'h0;
  assign T134 = idxPagesOH_1 & pageHit;
  assign idxPagesOH_1 = T135[2'h3:1'h0];
  assign T135 = 1'h1 << T136;
  assign T136 = idxPages[3'h1];
  assign T137 = {T142, T138};
  assign T138 = T139 != 4'h0;
  assign T139 = idxPagesOH_2 & pageHit;
  assign idxPagesOH_2 = T140[2'h3:1'h0];
  assign T140 = 1'h1 << T141;
  assign T141 = idxPages[3'h2];
  assign T142 = T143 != 4'h0;
  assign T143 = idxPagesOH_3 & pageHit;
  assign idxPagesOH_3 = T144[2'h3:1'h0];
  assign T144 = 1'h1 << T145;
  assign T145 = idxPages[3'h3];
  assign T146 = {T156, T147};
  assign T147 = {T152, T148};
  assign T148 = T149 != 4'h0;
  assign T149 = idxPagesOH_4 & pageHit;
  assign idxPagesOH_4 = T150[2'h3:1'h0];
  assign T150 = 1'h1 << T151;
  assign T151 = idxPages[3'h4];
  assign T152 = T153 != 4'h0;
  assign T153 = idxPagesOH_5 & pageHit;
  assign idxPagesOH_5 = T154[2'h3:1'h0];
  assign T154 = 1'h1 << T155;
  assign T155 = idxPages[3'h5];
  assign T156 = {T161, T157};
  assign T157 = T158 != 4'h0;
  assign T158 = idxPagesOH_6 & pageHit;
  assign idxPagesOH_6 = T159[2'h3:1'h0];
  assign T159 = 1'h1 << T160;
  assign T160 = idxPages[3'h6];
  assign T161 = T162 != 4'h0;
  assign T162 = idxPagesOH_7 & pageHit;
  assign idxPagesOH_7 = T163[2'h3:1'h0];
  assign T163 = 1'h1 << T164;
  assign T164 = idxPages[3'h7];
  assign T165 = idxValid & T166;
  assign T166 = T167;
  assign T167 = {T181, T168};
  assign T168 = {T176, T169};
  assign T169 = {T174, T170};
  assign T170 = T172 == T171;
  assign T171 = io_req_bits_addr[4'hb:1'h0];
  assign T172 = idxs[3'h0];
  assign T475 = R74[4'hb:1'h0];
  assign T174 = T175 == T171;
  assign T175 = idxs[3'h1];
  assign T176 = {T179, T177};
  assign T177 = T178 == T171;
  assign T178 = idxs[3'h2];
  assign T179 = T180 == T171;
  assign T180 = idxs[3'h3];
  assign T181 = {T187, T182};
  assign T182 = {T185, T183};
  assign T183 = T184 == T171;
  assign T184 = idxs[3'h4];
  assign T185 = T186 == T171;
  assign T186 = idxs[3'h5];
  assign T187 = {T190, T188};
  assign T188 = T189 == T171;
  assign T189 = idxs[3'h6];
  assign T190 = T191 == T171;
  assign T191 = idxs[3'h7];
  assign T476 = reset ? 8'h0 : T192;
  assign T192 = io_invalidate ? 8'h0 : T193;
  assign T193 = R7 ? T194 : idxValid;
  assign T194 = T196 | T195;
  assign T195 = 1'h1 << T42;
  assign T196 = idxValid & T197;
  assign T197 = ~ T198;
  assign T198 = T199;
  assign T199 = {T225, T200};
  assign T200 = {T214, T201};
  assign T201 = {T209, T202};
  assign T202 = T203 != 4'h0;
  assign T203 = pageReplEn & T204;
  assign T204 = idxPagesOH_0 | tgtPagesOH_0;
  assign tgtPagesOH_0 = T205[2'h3:1'h0];
  assign T205 = 1'h1 << T206;
  assign T206 = tgtPages[3'h0];
  assign T477 = {T482, T478};
  assign T478 = T479[1'h1:1'h1];
  assign T479 = T481 | T480;
  assign T480 = T208[1'h1:1'h0];
  assign T208 = usePageHit ? pageHit : tgtPageRepl;
  assign T481 = T208[2'h3:2'h2];
  assign T482 = T481 != 2'h0;
  assign T209 = T210 != 4'h0;
  assign T210 = pageReplEn & T211;
  assign T211 = idxPagesOH_1 | tgtPagesOH_1;
  assign tgtPagesOH_1 = T212[2'h3:1'h0];
  assign T212 = 1'h1 << T213;
  assign T213 = tgtPages[3'h1];
  assign T214 = {T220, T215};
  assign T215 = T216 != 4'h0;
  assign T216 = pageReplEn & T217;
  assign T217 = idxPagesOH_2 | tgtPagesOH_2;
  assign tgtPagesOH_2 = T218[2'h3:1'h0];
  assign T218 = 1'h1 << T219;
  assign T219 = tgtPages[3'h2];
  assign T220 = T221 != 4'h0;
  assign T221 = pageReplEn & T222;
  assign T222 = idxPagesOH_3 | tgtPagesOH_3;
  assign tgtPagesOH_3 = T223[2'h3:1'h0];
  assign T223 = 1'h1 << T224;
  assign T224 = tgtPages[3'h3];
  assign T225 = {T237, T226};
  assign T226 = {T232, T227};
  assign T227 = T228 != 4'h0;
  assign T228 = pageReplEn & T229;
  assign T229 = idxPagesOH_4 | tgtPagesOH_4;
  assign tgtPagesOH_4 = T230[2'h3:1'h0];
  assign T230 = 1'h1 << T231;
  assign T231 = tgtPages[3'h4];
  assign T232 = T233 != 4'h0;
  assign T233 = pageReplEn & T234;
  assign T234 = idxPagesOH_5 | tgtPagesOH_5;
  assign tgtPagesOH_5 = T235[2'h3:1'h0];
  assign T235 = 1'h1 << T236;
  assign T236 = tgtPages[3'h5];
  assign T237 = {T243, T238};
  assign T238 = T239 != 4'h0;
  assign T239 = pageReplEn & T240;
  assign T240 = idxPagesOH_6 | tgtPagesOH_6;
  assign tgtPagesOH_6 = T241[2'h3:1'h0];
  assign T241 = 1'h1 << T242;
  assign T242 = tgtPages[3'h6];
  assign T243 = T244 != 4'h0;
  assign T244 = pageReplEn & T245;
  assign T245 = idxPagesOH_7 | tgtPagesOH_7;
  assign tgtPagesOH_7 = T246[2'h3:1'h0];
  assign T246 = 1'h1 << T247;
  assign T247 = tgtPages[3'h7];
  assign T248 = T254 | T249;
  assign T249 = T253 ? isJump_6 : 1'h0;
  assign T250 = T251 ? R36 : isJump_6;
  assign T251 = R7 & T252;
  assign T252 = T40[3'h6:3'h6];
  assign T253 = hits[3'h6:3'h6];
  assign T254 = T260 | T255;
  assign T255 = T259 ? isJump_5 : 1'h0;
  assign T256 = T257 ? R36 : isJump_5;
  assign T257 = R7 & T258;
  assign T258 = T40[3'h5:3'h5];
  assign T259 = hits[3'h5:3'h5];
  assign T260 = T266 | T261;
  assign T261 = T265 ? isJump_4 : 1'h0;
  assign T262 = T263 ? R36 : isJump_4;
  assign T263 = R7 & T264;
  assign T264 = T40[3'h4:3'h4];
  assign T265 = hits[3'h4:3'h4];
  assign T266 = T272 | T267;
  assign T267 = T271 ? isJump_3 : 1'h0;
  assign T268 = T269 ? R36 : isJump_3;
  assign T269 = R7 & T270;
  assign T270 = T40[2'h3:2'h3];
  assign T271 = hits[2'h3:2'h3];
  assign T272 = T278 | T273;
  assign T273 = T277 ? isJump_2 : 1'h0;
  assign T274 = T275 ? R36 : isJump_2;
  assign T275 = R7 & T276;
  assign T276 = T40[2'h2:2'h2];
  assign T277 = hits[2'h2:2'h2];
  assign T278 = T284 | T279;
  assign T279 = T283 ? isJump_1 : 1'h0;
  assign T280 = T281 ? R36 : isJump_1;
  assign T281 = R7 & T282;
  assign T282 = T40[1'h1:1'h1];
  assign T283 = hits[1'h1:1'h1];
  assign T284 = T288 ? isJump_0 : 1'h0;
  assign T285 = T286 ? R36 : isJump_0;
  assign T286 = R7 & T287;
  assign T287 = T40[1'h0:1'h0];
  assign T288 = hits[1'h0:1'h0];
  assign T289 = io_req_valid & io_resp_valid;
  assign T290 = {io_bht_update_bits_taken, T291};
  assign T291 = io_bht_update_bits_prediction_bits_bht_history[2'h3:1'h1];
  assign T292 = T21 & io_bht_update_bits_mispredict;
  assign T293 = io_req_bits_addr[3'h5:2'h2];
  assign io_resp_bits_bht_history = T294;
  assign T294 = R25;
  assign io_resp_bits_entry = T483;
  assign T483 = {T493, T484};
  assign T484 = {T492, T485};
  assign T485 = T486[1'h1:1'h1];
  assign T486 = T491 | T487;
  assign T487 = T488[1'h1:1'h0];
  assign T488 = T490 | T489;
  assign T489 = hits[2'h3:1'h0];
  assign T490 = hits[3'h7:3'h4];
  assign T491 = T488[2'h3:2'h2];
  assign T492 = T491 != 2'h0;
  assign T493 = T490 != 4'h0;
  assign io_resp_bits_target = T296;
  assign T296 = T456 ? io_ras_update_bits_returnAddr : T297;
  assign T297 = T402 ? T369 : T298;
  assign T298 = {T331, T299};
  assign T299 = T304 | T300;
  assign T300 = T303 ? T301 : 12'h0;
  assign T301 = tgts[3'h7];
  assign T494 = io_req_bits_addr[4'hb:1'h0];
  assign T303 = hits[3'h7:3'h7];
  assign T304 = T308 | T305;
  assign T305 = T307 ? T306 : 12'h0;
  assign T306 = tgts[3'h6];
  assign T307 = hits[3'h6:3'h6];
  assign T308 = T312 | T309;
  assign T309 = T311 ? T310 : 12'h0;
  assign T310 = tgts[3'h5];
  assign T311 = hits[3'h5:3'h5];
  assign T312 = T316 | T313;
  assign T313 = T315 ? T314 : 12'h0;
  assign T314 = tgts[3'h4];
  assign T315 = hits[3'h4:3'h4];
  assign T316 = T320 | T317;
  assign T317 = T319 ? T318 : 12'h0;
  assign T318 = tgts[3'h3];
  assign T319 = hits[2'h3:2'h3];
  assign T320 = T324 | T321;
  assign T321 = T323 ? T322 : 12'h0;
  assign T322 = tgts[3'h2];
  assign T323 = hits[2'h2:2'h2];
  assign T324 = T328 | T325;
  assign T325 = T327 ? T326 : 12'h0;
  assign T326 = tgts[3'h1];
  assign T327 = hits[1'h1:1'h1];
  assign T328 = T330 ? T329 : 12'h0;
  assign T329 = tgts[3'h0];
  assign T330 = hits[1'h0:1'h0];
  assign T331 = T358 | T332;
  assign T332 = T334 ? T333 : 27'h0;
  assign T333 = pages[2'h3];
  assign T334 = T335[2'h3:2'h3];
  assign T335 = T338 | T336;
  assign T336 = T337 ? tgtPagesOH_7 : 4'h0;
  assign T337 = hits[3'h7:3'h7];
  assign T338 = T341 | T339;
  assign T339 = T340 ? tgtPagesOH_6 : 4'h0;
  assign T340 = hits[3'h6:3'h6];
  assign T341 = T344 | T342;
  assign T342 = T343 ? tgtPagesOH_5 : 4'h0;
  assign T343 = hits[3'h5:3'h5];
  assign T344 = T347 | T345;
  assign T345 = T346 ? tgtPagesOH_4 : 4'h0;
  assign T346 = hits[3'h4:3'h4];
  assign T347 = T350 | T348;
  assign T348 = T349 ? tgtPagesOH_3 : 4'h0;
  assign T349 = hits[2'h3:2'h3];
  assign T350 = T353 | T351;
  assign T351 = T352 ? tgtPagesOH_2 : 4'h0;
  assign T352 = hits[2'h2:2'h2];
  assign T353 = T356 | T354;
  assign T354 = T355 ? tgtPagesOH_1 : 4'h0;
  assign T355 = hits[1'h1:1'h1];
  assign T356 = T357 ? tgtPagesOH_0 : 4'h0;
  assign T357 = hits[1'h0:1'h0];
  assign T358 = T362 | T359;
  assign T359 = T361 ? T360 : 27'h0;
  assign T360 = pages[2'h2];
  assign T361 = T335[2'h2:2'h2];
  assign T362 = T366 | T363;
  assign T363 = T365 ? T364 : 27'h0;
  assign T364 = pages[2'h1];
  assign T365 = T335[1'h1:1'h1];
  assign T366 = T368 ? T367 : 27'h0;
  assign T367 = pages[2'h0];
  assign T368 = T335[1'h0:1'h0];
  assign T369 = T401 ? R397 : R370;
  assign T371 = T372 ? io_ras_update_bits_returnAddr : R370;
  assign T372 = T396 & T373;
  assign T373 = T374[1'h0:1'h0];
  assign T374 = 1'h1 << T375;
  assign T375 = T376;
  assign T376 = R377 + 1'h1;
  assign T495 = reset ? 1'h0 : T378;
  assign T378 = T381 ? T380 : T379;
  assign T379 = T396 ? T376 : R377;
  assign T380 = R377 - 1'h1;
  assign T381 = T392 & T382;
  assign T382 = T383 ^ 1'h1;
  assign T383 = R384 == 2'h0;
  assign T496 = reset ? 2'h0 : T385;
  assign T385 = io_invalidate ? 2'h0 : T386;
  assign T386 = T381 ? T391 : T387;
  assign T387 = T389 ? T388 : R384;
  assign T388 = R384 + 2'h1;
  assign T389 = T396 & T390;
  assign T390 = R384 < 2'h2;
  assign T391 = R384 - 2'h1;
  assign T392 = io_ras_update_valid & T393;
  assign T393 = T395 & T394;
  assign T394 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T395 = io_ras_update_bits_isCall ^ 1'h1;
  assign T396 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T398 = T399 ? io_ras_update_bits_returnAddr : R397;
  assign T399 = T396 & T400;
  assign T400 = T374[1'h1:1'h1];
  assign T401 = R377;
  assign T402 = T454 & T403;
  assign T403 = T413 | T404;
  assign T404 = T412 ? useRAS_7 : 1'h0;
  assign T405 = T408 ? R406 : useRAS_7;
  assign T407 = io_btb_update_valid ? io_btb_update_bits_isReturn : R406;
  assign T408 = R7 & T409;
  assign T409 = T410[3'h7:3'h7];
  assign T410 = 1'h1 << T411;
  assign T411 = T42;
  assign T412 = hits[3'h7:3'h7];
  assign T413 = T419 | T414;
  assign T414 = T418 ? useRAS_6 : 1'h0;
  assign T415 = T416 ? R406 : useRAS_6;
  assign T416 = R7 & T417;
  assign T417 = T410[3'h6:3'h6];
  assign T418 = hits[3'h6:3'h6];
  assign T419 = T425 | T420;
  assign T420 = T424 ? useRAS_5 : 1'h0;
  assign T421 = T422 ? R406 : useRAS_5;
  assign T422 = R7 & T423;
  assign T423 = T410[3'h5:3'h5];
  assign T424 = hits[3'h5:3'h5];
  assign T425 = T431 | T426;
  assign T426 = T430 ? useRAS_4 : 1'h0;
  assign T427 = T428 ? R406 : useRAS_4;
  assign T428 = R7 & T429;
  assign T429 = T410[3'h4:3'h4];
  assign T430 = hits[3'h4:3'h4];
  assign T431 = T437 | T432;
  assign T432 = T436 ? useRAS_3 : 1'h0;
  assign T433 = T434 ? R406 : useRAS_3;
  assign T434 = R7 & T435;
  assign T435 = T410[2'h3:2'h3];
  assign T436 = hits[2'h3:2'h3];
  assign T437 = T443 | T438;
  assign T438 = T442 ? useRAS_2 : 1'h0;
  assign T439 = T440 ? R406 : useRAS_2;
  assign T440 = R7 & T441;
  assign T441 = T410[2'h2:2'h2];
  assign T442 = hits[2'h2:2'h2];
  assign T443 = T449 | T444;
  assign T444 = T448 ? useRAS_1 : 1'h0;
  assign T445 = T446 ? R406 : useRAS_1;
  assign T446 = R7 & T447;
  assign T447 = T410[1'h1:1'h1];
  assign T448 = hits[1'h1:1'h1];
  assign T449 = T453 ? useRAS_0 : 1'h0;
  assign T450 = T451 ? R406 : useRAS_0;
  assign T451 = R7 & T452;
  assign T452 = T410[1'h0:1'h0];
  assign T453 = hits[1'h0:1'h0];
  assign T454 = T455 ^ 1'h1;
  assign T455 = R384 == 2'h0;
  assign T456 = T396 & T403;
  assign io_resp_bits_bridx = T457;
  assign T457 = brIdx[io_resp_bits_entry];
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_taken = T459;
  assign T459 = T460 ? 1'h0 : io_resp_valid;
  assign T460 = T461 & T32;
  assign T461 = T462 ^ 1'h1;
  assign T462 = T8[1'h0:1'h0];
  assign io_resp_valid = T463;
  assign T463 = hits != 8'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
// synthesis translate_on
`endif
    if(io_btb_update_valid) begin
      R4 <= io_btb_update_bits_target;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_btb_update_valid;
    end
    if (T21)
      T10[T22] <= T12;
    if(T292) begin
      R25 <= T290;
    end else if(T31) begin
      R25 <= T28;
    end
    if(T38) begin
      isJump_7 <= R36;
    end
    if(io_btb_update_valid) begin
      R36 <= io_btb_update_bits_isJump;
    end
    if(reset) begin
      nextRepl <= 3'h0;
    end else if(T45) begin
      nextRepl <= T44;
    end
    if(io_btb_update_valid) begin
      R47 <= io_btb_update_bits_prediction_bits_entry;
    end
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end
    if(reset) begin
      pageValid <= 4'h0;
    end else if(io_invalidate) begin
      pageValid <= 4'h0;
    end else if(T116) begin
      pageValid <= T59;
    end
    if(reset) begin
      R65 <= 2'h0;
    end else if(T68) begin
      R65 <= T67;
    end
    if(io_btb_update_valid) begin
      R74 <= io_btb_update_bits_pc;
    end
    if (T83)
      pages[2'h3] <= T78;
    if (T88)
      pages[2'h1] <= T78;
    if (T95)
      pages[2'h2] <= T92;
    if (T100)
      pages[2'h0] <= T92;
    if (R7)
      idxPages[T42] <= T469;
    if (R7)
      idxs[T42] <= T475;
    if(reset) begin
      idxValid <= 8'h0;
    end else if(io_invalidate) begin
      idxValid <= 8'h0;
    end else if(R7) begin
      idxValid <= T194;
    end
    if (R7)
      tgtPages[T42] <= T477;
    if(T251) begin
      isJump_6 <= R36;
    end
    if(T257) begin
      isJump_5 <= R36;
    end
    if(T263) begin
      isJump_4 <= R36;
    end
    if(T269) begin
      isJump_3 <= R36;
    end
    if(T275) begin
      isJump_2 <= R36;
    end
    if(T281) begin
      isJump_1 <= R36;
    end
    if(T286) begin
      isJump_0 <= R36;
    end
    if (R7)
      tgts[T42] <= T494;
    if(T372) begin
      R370 <= io_ras_update_bits_returnAddr;
    end
    if(reset) begin
      R377 <= 1'h0;
    end else if(T381) begin
      R377 <= T380;
    end else if(T396) begin
      R377 <= T376;
    end
    if(reset) begin
      R384 <= 2'h0;
    end else if(io_invalidate) begin
      R384 <= 2'h0;
    end else if(T381) begin
      R384 <= T391;
    end else if(T389) begin
      R384 <= T388;
    end
    if(T399) begin
      R397 <= io_ras_update_bits_returnAddr;
    end
    if(T408) begin
      useRAS_7 <= R406;
    end
    if(io_btb_update_valid) begin
      R406 <= io_btb_update_bits_isReturn;
    end
    if(T416) begin
      useRAS_6 <= R406;
    end
    if(T422) begin
      useRAS_5 <= R406;
    end
    if(T428) begin
      useRAS_4 <= R406;
    end
    if(T434) begin
      useRAS_3 <= R406;
    end
    if(T440) begin
      useRAS_2 <= R406;
    end
    if(T446) begin
      useRAS_1 <= R406;
    end
    if(T451) begin
      useRAS_0 <= R406;
    end
    if (R7)
      brIdx[T42] <= 1'h0;
  end
endmodule

module FlowThroughSerializer(
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_addr_beat,
    input [1:0] io_in_bits_client_xact_id,
    input [2:0] io_in_bits_manager_xact_id,
    input  io_in_bits_is_builtin_type,
    input [3:0] io_in_bits_g_type,
    input [127:0] io_in_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_manager_xact_id,
    output io_out_bits_is_builtin_type,
    output[3:0] io_out_bits_g_type,
    output[127:0] io_out_bits_data,
    output io_cnt,
    output io_done
);



  assign io_done = 1'h1;
  assign io_cnt = 1'h0;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_valid = io_in_valid;
  assign io_in_ready = io_out_ready;
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [11:0] io_req_bits_idx,
    input [19:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    //output[31:0] io_resp_bits_data
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data
);

  wire[127:0] T0;
  wire[16:0] T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[25:0] T7;
  reg [31:0] refill_addr;
  wire[31:0] T8;
  wire[31:0] s1_addr;
  wire[31:0] T9;
  reg [11:0] s1_pgoff;
  wire[11:0] T10;
  wire T11;
  wire rdy;
  wire T12;
  wire T13;
  wire s1_miss;
  wire T14;
  wire s1_any_tag_hit;
  wire T15;
  wire T16;
  wire s1_disparity_0;
  wire s1_tag_hit_0;
  wire T17;
  wire s1_tag_match_0;
  wire T18;
  wire[19:0] s1_tag;
  wire[19:0] T19;
  wire[19:0] T20;
  wire T51;
  wire s0_valid;
  wire T52;
  wire stall;
  reg  s1_valid;
  wire T109;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T53;
  wire refill_done;
  wire refill_wrap;
  wire T25;
  reg [1:0] refill_cnt;
  wire[1:0] T110;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire T29;
  reg [1:0] state;
  wire[1:0] T111;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[5:0] T44;
  wire[11:0] s0_pgoff;
  wire T45;
  wire[19:0] T21;
  wire[19:0] T22;
  wire[19:0] T23;
  wire[19:0] T24;
  wire[19:0] refill_tag;
  wire[5:0] s1_idx;
  reg [5:0] R42;
  wire[5:0] T43;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[5:0] T62;
  wire T63;
  reg [63:0] vb_array;
  wire[63:0] T112;
  wire[127:0] T113;
  wire[127:0] T64;
  wire[127:0] T65;
  wire[127:0] T66;
  wire[127:0] T114;
  wire[127:0] T67;
  wire[127:0] T68;
  wire[127:0] T69;
  wire[6:0] T70;
  wire[127:0] T115;
  wire T71;
  wire[127:0] T72;
  wire[127:0] T73;
  wire[127:0] T116;
  wire T74;
  wire T75;
  reg  invalidated;
  wire T76;
  wire T77;
  wire[127:0] T78;
  wire[127:0] T79;
  wire[127:0] T80;
  wire[6:0] T81;
  wire[127:0] T117;
  wire T82;
  wire[127:0] T83;
  wire[127:0] T84;
  wire[127:0] T118;
  wire T85;
  wire T86;
  wire out_valid;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire[127:0] s1_dout_0;
  wire[127:0] T95;
  wire[127:0] T96;
  wire T104;
  wire T105;
  wire[7:0] T103;
  wire[127:0] T98;
  wire[127:0] T99;
  wire[7:0] T100;
  reg [7:0] R101;
  wire[7:0] T102;
  wire T106;
  wire T107;
  wire T108;
  wire s1_hit;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    refill_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    s1_valid = {1{$random}};
    refill_cnt = {1{$random}};
    state = {1{$random}};
    R42 = {1{$random}};
    vb_array = {2{$random}};
    invalidated = {1{$random}};
    R101 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_resp_bits_data = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = T0;
  assign T0 = 128'h0;
  assign io_mem_acquire_bits_union = T1;
  assign T1 = 17'h1c1;
  assign io_mem_acquire_bits_a_type = T2;
  assign T2 = 3'h1;
  assign io_mem_acquire_bits_is_builtin_type = T3;
  assign T3 = 1'h1;
  assign io_mem_acquire_bits_addr_beat = T4;
  assign T4 = 2'h0;
  assign io_mem_acquire_bits_client_xact_id = T5;
  assign T5 = 2'h0;
  assign io_mem_acquire_bits_addr_block = T6;
  assign T6 = T7;
  assign T7 = refill_addr >> 3'h6;
  assign T8 = T91 ? s1_addr : refill_addr;
  assign s1_addr = T9;
  assign T9 = {io_req_bits_ppn, s1_pgoff};
  assign T10 = T11 ? io_req_bits_idx : s1_pgoff;
  assign T11 = io_req_valid & rdy;
  assign rdy = T12;
  assign T12 = T90 & T13;
  assign T13 = s1_miss ^ 1'h1;
  assign s1_miss = out_valid & T14;
  assign T14 = s1_any_tag_hit ^ 1'h1;
  assign s1_any_tag_hit = T15;
  assign T15 = s1_tag_hit_0 & T16;
  assign T16 = s1_disparity_0 ^ 1'h1;
  assign s1_disparity_0 = 1'h0;
  assign s1_tag_hit_0 = T17;
  assign T17 = T54 & s1_tag_match_0;
  assign s1_tag_match_0 = T18;
  assign T18 = T19 == s1_tag;
  assign s1_tag = s1_addr[5'h1f:4'hc];
  assign T19 = T20[5'h13:1'h0];
  assign T51 = T53 & s0_valid;
  assign s0_valid = io_req_valid | T52;
  assign T52 = s1_valid & stall;
  assign stall = io_resp_ready ^ 1'h1;
  assign T109 = reset ? 1'h0 : T46;
  assign T46 = T50 | T47;
  assign T47 = T49 & T48;
  assign T48 = io_req_bits_kill ^ 1'h1;
  assign T49 = s1_valid & stall;
  assign T50 = io_req_valid & rdy;
  assign T53 = refill_done ^ 1'h1;
  assign refill_done = T29 & refill_wrap;
  assign refill_wrap = T28 & T25;
  assign T25 = refill_cnt == 2'h3;
  assign T110 = reset ? 2'h0 : T26;
  assign T26 = T28 ? T27 : refill_cnt;
  assign T27 = refill_cnt + 2'h1;
  assign T28 = 1'h1 & FlowThroughSerializer_io_out_valid;
  assign T29 = state == 2'h3;
  assign T111 = reset ? 2'h0 : T30;
  assign T30 = T40 ? 2'h0 : T31;
  assign T31 = T38 ? 2'h3 : T32;
  assign T32 = T36 ? 2'h2 : T33;
  assign T33 = T34 ? 2'h1 : state;
  assign T34 = T35 & s1_miss;
  assign T35 = 2'h0 == state;
  assign T36 = T37 & io_mem_acquire_ready;
  assign T37 = 2'h1 == state;
  assign T38 = T39 & io_mem_grant_valid;
  assign T39 = 2'h2 == state;
  assign T40 = T41 & refill_done;
  assign T41 = 2'h3 == state;
  assign T44 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T45 ? s1_pgoff : io_req_bits_idx;
  assign T45 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(refill_done ? s1_idx : T44),
    .RW0E(T51 || refill_done),
    .RW0W(refill_done),
    .RW0I(T23),
    .RW0M(T22),
    .RW0O(T20)
  );
  assign T22 = 20'hfffff;
  assign T23 = T24;
  assign T24 = refill_tag;
  assign refill_tag = refill_addr[5'h1f:4'hc];
  assign s1_idx = s1_addr[4'hb:3'h6];
  assign T43 = T51 ? T44 : R42;
  assign T54 = T86 & T55;
  assign T55 = T56;
  assign T56 = T63 & T57;
  assign T57 = T58 - 1'h1;
  assign T58 = 1'h1 << T59;
  assign T59 = T60 + 7'h1;
  assign T60 = T61 - T61;
  assign T61 = {1'h0, T62};
  assign T62 = s1_pgoff[4'hb:3'h6];
  assign T63 = vb_array >> T61;
  assign T112 = T113[6'h3f:1'h0];
  assign T113 = reset ? 128'h0 : T64;
  assign T64 = T85 ? T78 : T65;
  assign T65 = io_invalidate ? 128'h0 : T66;
  assign T66 = T74 ? T67 : T114;
  assign T114 = {64'h0, vb_array};
  assign T67 = T72 | T68;
  assign T68 = T115 & T69;
  assign T69 = 1'h1 << T70;
  assign T70 = {1'h0, s1_idx};
  assign T115 = T71 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T71 = 1'h1;
  assign T72 = T116 & T73;
  assign T73 = ~ T69;
  assign T116 = {64'h0, vb_array};
  assign T74 = refill_done & T75;
  assign T75 = invalidated ^ 1'h1;
  assign T76 = T35 ? 1'h0 : T77;
  assign T77 = io_invalidate ? 1'h1 : invalidated;
  assign T78 = T83 | T79;
  assign T79 = T117 & T80;
  assign T80 = 1'h1 << T81;
  assign T81 = {1'h0, s1_idx};
  assign T117 = T82 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T82 = 1'h0;
  assign T83 = T118 & T84;
  assign T84 = ~ T80;
  assign T118 = {64'h0, vb_array};
  assign T85 = s1_valid & s1_disparity_0;
  assign T86 = io_invalidate ^ 1'h1;
  assign out_valid = T88 & T87;
  assign T87 = state == 2'h0;
  assign T88 = s1_valid & T89;
  assign T89 = io_req_bits_kill ^ 1'h1;
  assign T90 = state == 2'h0;
  assign T91 = T92 & s1_miss;
  assign T92 = s1_valid & T93;
  assign T93 = state == 2'h0;
  assign io_mem_acquire_valid = T94;
  assign T94 = state == 2'h1;
  assign io_resp_bits_datablock = s1_dout_0;
  assign s1_dout_0 = T95;
  assign T95 = T106 ? T96 : 128'h0;
  assign T104 = T105 & s0_valid;
  assign T105 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T103 = s0_pgoff[4'hb:3'h4];
  ICache_T97 T97 (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_io_out_valid ? T100 : T103),
    .RW0E(T104 || FlowThroughSerializer_io_out_valid),
    .RW0W(FlowThroughSerializer_io_out_valid),
    .RW0I(T99),
    .RW0O(T96)
  );
  assign T99 = FlowThroughSerializer_io_out_bits_data;
  assign T100 = {s1_idx, refill_cnt};
  assign T102 = T104 ? T103 : R101;
  assign T106 = T108 & T107;
  assign T107 = stall ^ 1'h1;
  assign T108 = s1_valid & rdy;
  assign io_resp_valid = s1_hit;
  assign s1_hit = out_valid & s1_any_tag_hit;
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       //.io_out_bits_addr_beat(  )
       //.io_out_bits_client_xact_id(  )
       //.io_out_bits_manager_xact_id(  )
       //.io_out_bits_is_builtin_type(  )
       //.io_out_bits_g_type(  )
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );

  always @(posedge clk) begin
    if(T91) begin
      refill_addr <= s1_addr;
    end
    if(T11) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T46;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T28) begin
      refill_cnt <= T27;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T40) begin
      state <= 2'h0;
    end else if(T38) begin
      state <= 2'h3;
    end else if(T36) begin
      state <= 2'h2;
    end else if(T34) begin
      state <= 2'h1;
    end
    if(T51) begin
      R42 <= T44;
    end
    vb_array <= T112;
    if(T35) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(T104) begin
      R101 <= T103;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input [3:0] io_clear_mask,
    input [33:0] io_tag,
    output io_hit,
    output[3:0] io_hits,
    output[3:0] io_valid_bits,
    input  io_write,
    input [33:0] io_write_tag,
    input [1:0] io_write_addr
);

  reg [3:0] vb_array;
  wire[3:0] T28;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T29;
  wire T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[1:0] T12;
  wire hits_0;
  wire T13;
  wire[33:0] T14;
  reg [33:0] cam_tags [3:0];
  wire[33:0] T15;
  wire T16;
  wire hits_1;
  wire T17;
  wire[33:0] T18;
  wire T19;
  wire[1:0] T20;
  wire hits_2;
  wire T21;
  wire[33:0] T22;
  wire T23;
  wire hits_3;
  wire T24;
  wire[33:0] T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_valid_bits = vb_array;
  assign T28 = reset ? 4'h0 : T0;
  assign T0 = io_clear ? T8 : T1;
  assign T1 = io_write ? T2 : vb_array;
  assign T2 = T6 | T3;
  assign T3 = T29 & T4;
  assign T4 = 1'h1 << io_write_addr;
  assign T29 = T5 ? 4'hf : 4'h0;
  assign T5 = 1'h1;
  assign T6 = vb_array & T7;
  assign T7 = ~ T4;
  assign T8 = vb_array & T9;
  assign T9 = ~ io_clear_mask;
  assign io_hits = T10;
  assign T10 = T11;
  assign T11 = {T20, T12};
  assign T12 = {hits_1, hits_0};
  assign hits_0 = T16 & T13;
  assign T13 = T14 == io_tag;
  assign T14 = cam_tags[2'h0];
  assign T16 = vb_array[1'h0:1'h0];
  assign hits_1 = T19 & T17;
  assign T17 = T18 == io_tag;
  assign T18 = cam_tags[2'h1];
  assign T19 = vb_array[1'h1:1'h1];
  assign T20 = {hits_3, hits_2};
  assign hits_2 = T23 & T21;
  assign T21 = T22 == io_tag;
  assign T22 = cam_tags[2'h2];
  assign T23 = vb_array[2'h2:2'h2];
  assign hits_3 = T26 & T24;
  assign T24 = T25 == io_tag;
  assign T25 = cam_tags[2'h3];
  assign T26 = vb_array[2'h3:2'h3];
  assign io_hit = T27;
  assign T27 = io_hits != 4'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 4'h0;
    end else if(io_clear) begin
      vb_array <= T8;
    end else if(io_write) begin
      vb_array <= T2;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [27:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    input  io_req_bits_store,
    output io_resp_miss,
    output[19:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    output[3:0] io_resp_hit_idx,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate
);

  reg [1:0] r_refill_waddr;
  wire[1:0] T0;
  wire[1:0] repl_waddr;
  wire[1:0] T1;
  wire[2:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  reg [3:0] R9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[6:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T349;
  wire T350;
  wire[1:0] T351;
  wire[1:0] T352;
  wire[1:0] T353;
  wire T354;
  wire T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire[3:0] T22;
  wire[3:0] T23;
  wire T24;
  wire tlb_hit;
  wire tag_hit;
  wire[3:0] tag_hits;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] w_array;
  wire[3:0] T28;
  wire[3:0] T29;
  wire[1:0] T30;
  reg  uw_array_0;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire[3:0] T42;
  wire[1:0] T43;
  reg  uw_array_1;
  wire T44;
  wire T45;
  wire T46;
  wire[1:0] T47;
  reg  uw_array_2;
  wire T48;
  wire T49;
  wire T50;
  reg  uw_array_3;
  wire T51;
  wire T52;
  wire T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[1:0] T56;
  reg  sw_array_0;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[1:0] T67;
  reg  sw_array_1;
  wire T68;
  wire T69;
  wire T70;
  wire[1:0] T71;
  reg  sw_array_2;
  wire T72;
  wire T73;
  wire T74;
  reg  sw_array_3;
  wire T75;
  wire T76;
  wire T77;
  wire priv_s;
  wire[1:0] priv;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[1:0] T82;
  reg  dirty_array_0;
  wire T83;
  wire T84;
  wire T85;
  wire[3:0] T86;
  wire[1:0] T87;
  reg  dirty_array_1;
  wire T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  reg  dirty_array_2;
  wire T92;
  wire T93;
  wire T94;
  reg  dirty_array_3;
  wire T95;
  wire T96;
  wire T97;
  wire vm_enabled;
  wire T98;
  wire T99;
  wire priv_uses_vm;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire T358;
  wire[3:0] T103;
  wire T359;
  wire T360;
  wire has_invalid_entry;
  wire T104;
  wire T105;
  wire tlb_miss;
  wire T106;
  wire bad_va;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire[33:0] T361;
  reg [34:0] r_refill_tag;
  wire[34:0] T112;
  wire[34:0] lookup_tag;
  wire[34:0] T113;
  wire T114;
  wire T115;
  reg [1:0] state;
  wire[1:0] T362;
  wire[1:0] T116;
  wire[1:0] T117;
  wire[1:0] T118;
  wire[1:0] T119;
  wire[1:0] T120;
  wire[1:0] T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire[33:0] T363;
  wire[3:0] T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[3:0] T132;
  wire[3:0] T133;
  wire[3:0] T134;
  wire[1:0] T135;
  reg  valid_array_0;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[3:0] T140;
  wire[1:0] T141;
  reg  valid_array_1;
  wire T142;
  wire T143;
  wire T144;
  wire[1:0] T145;
  reg  valid_array_2;
  wire T146;
  wire T147;
  wire T148;
  reg  valid_array_3;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  reg  r_req_instruction;
  wire T154;
  reg  r_req_store;
  wire T155;
  wire[26:0] T364;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[3:0] T161;
  wire[3:0] x_array;
  wire[3:0] T162;
  wire[3:0] T163;
  wire[1:0] T164;
  reg  ux_array_0;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire[3:0] T176;
  wire[1:0] T177;
  reg  ux_array_1;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  reg  ux_array_2;
  wire T182;
  wire T183;
  wire T184;
  reg  ux_array_3;
  wire T185;
  wire T186;
  wire T187;
  wire[3:0] T188;
  wire[3:0] T189;
  wire[1:0] T190;
  reg  sx_array_0;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[3:0] T200;
  wire[1:0] T201;
  reg  sx_array_1;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  reg  sx_array_2;
  wire T206;
  wire T207;
  wire T208;
  reg  sx_array_3;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[2:0] T216;
  wire[2:0] T217;
  wire[2:0] T218;
  wire T219;
  wire T220;
  wire[32:0] T365;
  wire[31:0] paddr;
  wire T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire[2:0] T224;
  wire T225;
  wire T226;
  wire T227;
  wire[2:0] T228;
  wire[2:0] T229;
  wire[2:0] T230;
  wire T231;
  wire T232;
  wire T233;
  wire[2:0] T234;
  wire[2:0] T235;
  wire[2:0] T236;
  wire T237;
  wire T238;
  wire T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire addr_ok;
  wire T246;
  wire T247;
  wire[32:0] T366;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[3:0] T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[3:0] T278;
  wire[3:0] r_array;
  wire[3:0] T279;
  wire[3:0] T280;
  wire[1:0] T281;
  reg  ur_array_0;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[1:0] T292;
  reg  ur_array_1;
  wire T293;
  wire T294;
  wire T295;
  wire[1:0] T296;
  reg  ur_array_2;
  wire T297;
  wire T298;
  wire T299;
  reg  ur_array_3;
  wire T300;
  wire T301;
  wire T302;
  wire[3:0] T303;
  wire[3:0] T304;
  wire[1:0] T305;
  reg  sr_array_0;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[1:0] T314;
  reg  sr_array_1;
  wire T315;
  wire T316;
  wire T317;
  wire[1:0] T318;
  reg  sr_array_2;
  wire T319;
  wire T320;
  wire T321;
  reg  sr_array_3;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[19:0] T330;
  wire[19:0] T331;
  wire[19:0] T332;
  wire[19:0] T333;
  wire[19:0] T334;
  reg [19:0] tag_ram [3:0];
  wire[19:0] T335;
  wire T336;
  wire[19:0] T337;
  wire[19:0] T338;
  wire[19:0] T339;
  wire T340;
  wire[19:0] T341;
  wire[19:0] T342;
  wire[19:0] T343;
  wire T344;
  wire[19:0] T345;
  wire[19:0] T346;
  wire T347;
  wire T348;
  wire[3:0] tag_cam_io_hits;
  wire[3:0] tag_cam_io_valid_bits;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R9 = {1{$random}};
    uw_array_0 = {1{$random}};
    uw_array_1 = {1{$random}};
    uw_array_2 = {1{$random}};
    uw_array_3 = {1{$random}};
    sw_array_0 = {1{$random}};
    sw_array_1 = {1{$random}};
    sw_array_2 = {1{$random}};
    sw_array_3 = {1{$random}};
    dirty_array_0 = {1{$random}};
    dirty_array_1 = {1{$random}};
    dirty_array_2 = {1{$random}};
    dirty_array_3 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    valid_array_0 = {1{$random}};
    valid_array_1 = {1{$random}};
    valid_array_2 = {1{$random}};
    valid_array_3 = {1{$random}};
    r_req_instruction = {1{$random}};
    r_req_store = {1{$random}};
    ux_array_0 = {1{$random}};
    ux_array_1 = {1{$random}};
    ux_array_2 = {1{$random}};
    ux_array_3 = {1{$random}};
    sx_array_0 = {1{$random}};
    sx_array_1 = {1{$random}};
    sx_array_2 = {1{$random}};
    sx_array_3 = {1{$random}};
    ur_array_0 = {1{$random}};
    ur_array_1 = {1{$random}};
    ur_array_2 = {1{$random}};
    ur_array_3 = {1{$random}};
    sr_array_0 = {1{$random}};
    sr_array_1 = {1{$random}};
    sr_array_2 = {1{$random}};
    sr_array_3 = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T105 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T355 : T1;
  assign T1 = T2[1'h1:1'h0];
  assign T2 = {T101, T3};
  assign T3 = T8 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 2'h1;
  assign T7 = T101 - T101;
  assign T8 = R9 >> T101;
  assign T10 = T24 ? T11 : R9;
  assign T11 = T19 | T12;
  assign T12 = T18 ? 4'h0 : T13;
  assign T13 = T14[2'h3:1'h0];
  assign T14 = 4'h1 << T15;
  assign T15 = {1'h1, T16};
  assign T16 = T349[1'h1:1'h1];
  assign T349 = {T354, T350};
  assign T350 = T351[1'h1:1'h1];
  assign T351 = T353 | T352;
  assign T352 = tag_cam_io_hits[1'h1:1'h0];
  assign T353 = tag_cam_io_hits[2'h3:2'h2];
  assign T354 = T353 != 2'h0;
  assign T18 = T349[1'h0:1'h0];
  assign T19 = T21 & T20;
  assign T20 = ~ T13;
  assign T21 = T23 | T22;
  assign T22 = T16 ? 4'h0 : 4'h2;
  assign T23 = R9 & 4'hd;
  assign T24 = io_req_valid & tlb_hit;
  assign tlb_hit = vm_enabled & tag_hit;
  assign tag_hit = tag_hits != 4'h0;
  assign tag_hits = tag_cam_io_hits & T25;
  assign T25 = T80 | T26;
  assign T26 = ~ T27;
  assign T27 = io_req_bits_store ? w_array : 4'h0;
  assign w_array = priv_s ? T54 : T28;
  assign T28 = T29;
  assign T29 = {T47, T30};
  assign T30 = {uw_array_1, uw_array_0};
  assign T31 = T40 ? T32 : uw_array_0;
  assign T32 = T34 & T33;
  assign T33 = io_ptw_resp_bits_error ^ 1'h1;
  assign T34 = T36 & T35;
  assign T35 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T36 = T38 & T37;
  assign T37 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T38 = io_ptw_resp_bits_pte_v & T39;
  assign T39 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T40 = io_ptw_resp_valid & T41;
  assign T41 = T42[1'h0:1'h0];
  assign T42 = 1'h1 << T43;
  assign T43 = r_refill_waddr;
  assign T44 = T45 ? T32 : uw_array_1;
  assign T45 = io_ptw_resp_valid & T46;
  assign T46 = T42[1'h1:1'h1];
  assign T47 = {uw_array_3, uw_array_2};
  assign T48 = T49 ? T32 : uw_array_2;
  assign T49 = io_ptw_resp_valid & T50;
  assign T50 = T42[2'h2:2'h2];
  assign T51 = T52 ? T32 : uw_array_3;
  assign T52 = io_ptw_resp_valid & T53;
  assign T53 = T42[2'h3:2'h3];
  assign T54 = T55;
  assign T55 = {T71, T56};
  assign T56 = {sw_array_1, sw_array_0};
  assign T57 = T64 ? T58 : sw_array_0;
  assign T58 = T60 & T59;
  assign T59 = io_ptw_resp_bits_error ^ 1'h1;
  assign T60 = T62 & T61;
  assign T61 = io_ptw_resp_bits_pte_typ[1'h0:1'h0];
  assign T62 = io_ptw_resp_bits_pte_v & T63;
  assign T63 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T64 = io_ptw_resp_valid & T65;
  assign T65 = T66[1'h0:1'h0];
  assign T66 = 1'h1 << T67;
  assign T67 = r_refill_waddr;
  assign T68 = T69 ? T58 : sw_array_1;
  assign T69 = io_ptw_resp_valid & T70;
  assign T70 = T66[1'h1:1'h1];
  assign T71 = {sw_array_3, sw_array_2};
  assign T72 = T73 ? T58 : sw_array_2;
  assign T73 = io_ptw_resp_valid & T74;
  assign T74 = T66[2'h2:2'h2];
  assign T75 = T76 ? T58 : sw_array_3;
  assign T76 = io_ptw_resp_valid & T77;
  assign T77 = T66[2'h3:2'h3];
  assign priv_s = priv == 2'h1;
  assign priv = T78 ? io_ptw_status_prv1 : io_ptw_status_prv;
  assign T78 = io_ptw_status_mprv & T79;
  assign T79 = io_req_bits_instruction ^ 1'h1;
  assign T80 = T81;
  assign T81 = {T91, T82};
  assign T82 = {dirty_array_1, dirty_array_0};
  assign T83 = T84 ? io_ptw_resp_bits_pte_d : dirty_array_0;
  assign T84 = io_ptw_resp_valid & T85;
  assign T85 = T86[1'h0:1'h0];
  assign T86 = 1'h1 << T87;
  assign T87 = r_refill_waddr;
  assign T88 = T89 ? io_ptw_resp_bits_pte_d : dirty_array_1;
  assign T89 = io_ptw_resp_valid & T90;
  assign T90 = T86[1'h1:1'h1];
  assign T91 = {dirty_array_3, dirty_array_2};
  assign T92 = T93 ? io_ptw_resp_bits_pte_d : dirty_array_2;
  assign T93 = io_ptw_resp_valid & T94;
  assign T94 = T86[2'h2:2'h2];
  assign T95 = T96 ? io_ptw_resp_bits_pte_d : dirty_array_3;
  assign T96 = io_ptw_resp_valid & T97;
  assign T97 = T86[2'h3:2'h3];
  assign vm_enabled = T99 & T98;
  assign T98 = io_req_bits_passthrough ^ 1'h1;
  assign T99 = T100 & priv_uses_vm;
  assign priv_uses_vm = priv <= 2'h1;
  assign T100 = io_ptw_status_vm[2'h3:2'h3];
  assign T101 = {1'h1, T102};
  assign T102 = R9[1'h1:1'h1];
  assign T355 = T360 ? 1'h0 : T356;
  assign T356 = T359 ? 1'h1 : T357;
  assign T357 = T358 ? 2'h2 : 2'h3;
  assign T358 = T103[2'h2:2'h2];
  assign T103 = ~ tag_cam_io_valid_bits;
  assign T359 = T103[1'h1:1'h1];
  assign T360 = T103[1'h0:1'h0];
  assign has_invalid_entry = T104 ^ 1'h1;
  assign T104 = tag_cam_io_valid_bits == 4'hf;
  assign T105 = T111 & tlb_miss;
  assign tlb_miss = T109 & T106;
  assign T106 = bad_va ^ 1'h1;
  assign bad_va = T108 != T107;
  assign T107 = io_req_bits_vpn[5'h1a:5'h1a];
  assign T108 = io_req_bits_vpn[5'h1b:5'h1b];
  assign T109 = vm_enabled & T110;
  assign T110 = tag_hit ^ 1'h1;
  assign T111 = io_req_ready & io_req_valid;
  assign T361 = r_refill_tag[6'h21:1'h0];
  assign T112 = T105 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T113;
  assign T113 = {io_req_bits_asid, io_req_bits_vpn};
  assign T114 = T115 & io_ptw_resp_valid;
  assign T115 = state == 2'h2;
  assign T362 = reset ? 2'h0 : T116;
  assign T116 = io_ptw_resp_valid ? 2'h0 : T117;
  assign T117 = T126 ? 2'h3 : T118;
  assign T118 = T125 ? 2'h3 : T119;
  assign T119 = T124 ? 2'h2 : T120;
  assign T120 = T122 ? 2'h0 : T121;
  assign T121 = T105 ? 2'h1 : state;
  assign T122 = T123 & io_ptw_invalidate;
  assign T123 = state == 2'h1;
  assign T124 = T123 & io_ptw_req_ready;
  assign T125 = T124 & io_ptw_invalidate;
  assign T126 = T127 & io_ptw_invalidate;
  assign T127 = state == 2'h2;
  assign T363 = lookup_tag[6'h21:1'h0];
  assign T128 = io_ptw_invalidate ? 4'hf : T129;
  assign T129 = T132 | T130;
  assign T130 = tag_cam_io_hits & T131;
  assign T131 = ~ tag_hits;
  assign T132 = ~ T133;
  assign T133 = T134;
  assign T134 = {T145, T135};
  assign T135 = {valid_array_1, valid_array_0};
  assign T136 = T138 ? T137 : valid_array_0;
  assign T137 = io_ptw_resp_bits_error ^ 1'h1;
  assign T138 = io_ptw_resp_valid & T139;
  assign T139 = T140[1'h0:1'h0];
  assign T140 = 1'h1 << T141;
  assign T141 = r_refill_waddr;
  assign T142 = T143 ? T137 : valid_array_1;
  assign T143 = io_ptw_resp_valid & T144;
  assign T144 = T140[1'h1:1'h1];
  assign T145 = {valid_array_3, valid_array_2};
  assign T146 = T147 ? T137 : valid_array_2;
  assign T147 = io_ptw_resp_valid & T148;
  assign T148 = T140[2'h2:2'h2];
  assign T149 = T150 ? T137 : valid_array_3;
  assign T150 = io_ptw_resp_valid & T151;
  assign T151 = T140[2'h3:2'h3];
  assign T152 = io_ptw_invalidate | T153;
  assign T153 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T154 = T105 ? io_req_bits_instruction : r_req_instruction;
  assign io_ptw_req_bits_store = r_req_store;
  assign T155 = T105 ? io_req_bits_store : r_req_store;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_addr = T364;
  assign T364 = r_refill_tag[5'h1a:1'h0];
  assign io_ptw_req_valid = T156;
  assign T156 = state == 2'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_xcpt_if = T157;
  assign T157 = T212 | T158;
  assign T158 = tlb_hit & T159;
  assign T159 = T160 ^ 1'h1;
  assign T160 = T161 != 4'h0;
  assign T161 = x_array & tag_cam_io_hits;
  assign x_array = priv_s ? T188 : T162;
  assign T162 = T163;
  assign T163 = {T181, T164};
  assign T164 = {ux_array_1, ux_array_0};
  assign T165 = T174 ? T166 : ux_array_0;
  assign T166 = T168 & T167;
  assign T167 = io_ptw_resp_bits_error ^ 1'h1;
  assign T168 = T170 & T169;
  assign T169 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T170 = T172 & T171;
  assign T171 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T172 = io_ptw_resp_bits_pte_v & T173;
  assign T173 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T174 = io_ptw_resp_valid & T175;
  assign T175 = T176[1'h0:1'h0];
  assign T176 = 1'h1 << T177;
  assign T177 = r_refill_waddr;
  assign T178 = T179 ? T166 : ux_array_1;
  assign T179 = io_ptw_resp_valid & T180;
  assign T180 = T176[1'h1:1'h1];
  assign T181 = {ux_array_3, ux_array_2};
  assign T182 = T183 ? T166 : ux_array_2;
  assign T183 = io_ptw_resp_valid & T184;
  assign T184 = T176[2'h2:2'h2];
  assign T185 = T186 ? T166 : ux_array_3;
  assign T186 = io_ptw_resp_valid & T187;
  assign T187 = T176[2'h3:2'h3];
  assign T188 = T189;
  assign T189 = {T205, T190};
  assign T190 = {sx_array_1, sx_array_0};
  assign T191 = T198 ? T192 : sx_array_0;
  assign T192 = T194 & T193;
  assign T193 = io_ptw_resp_bits_error ^ 1'h1;
  assign T194 = T196 & T195;
  assign T195 = io_ptw_resp_bits_pte_typ[1'h1:1'h1];
  assign T196 = io_ptw_resp_bits_pte_v & T197;
  assign T197 = 4'h4 <= io_ptw_resp_bits_pte_typ;
  assign T198 = io_ptw_resp_valid & T199;
  assign T199 = T200[1'h0:1'h0];
  assign T200 = 1'h1 << T201;
  assign T201 = r_refill_waddr;
  assign T202 = T203 ? T192 : sx_array_1;
  assign T203 = io_ptw_resp_valid & T204;
  assign T204 = T200[1'h1:1'h1];
  assign T205 = {sx_array_3, sx_array_2};
  assign T206 = T207 ? T192 : sx_array_2;
  assign T207 = io_ptw_resp_valid & T208;
  assign T208 = T200[2'h2:2'h2];
  assign T209 = T210 ? T192 : sx_array_3;
  assign T210 = io_ptw_resp_valid & T211;
  assign T211 = T200[2'h3:2'h3];
  assign T212 = T213 | bad_va;
  assign T213 = T245 | T214;
  assign T214 = T215 ^ 1'h1;
  assign T215 = T216[2'h2:2'h2];
  assign T216 = T222 | T217;
  assign T217 = T219 ? T218 : 3'h0;
  assign T218 = 3'h3;
  assign T219 = T221 & T220;
  assign T220 = T365 < 33'h100000000;
  assign T365 = {1'h0, paddr};
  assign paddr = {io_resp_ppn, 12'h0};
  assign T221 = 32'h80000000 <= paddr;
  assign T222 = T228 | T223;
  assign T223 = T225 ? T224 : 3'h0;
  assign T224 = 3'h3;
  assign T225 = T227 & T226;
  assign T226 = paddr < 32'h40010200;
  assign T227 = 32'h40010000 <= paddr;
  assign T228 = T234 | T229;
  assign T229 = T231 ? T230 : 3'h0;
  assign T230 = 3'h3;
  assign T231 = T233 & T232;
  assign T232 = paddr < 32'h40010000;
  assign T233 = 32'h40008000 <= paddr;
  assign T234 = T240 | T235;
  assign T235 = T237 ? T236 : 3'h0;
  assign T236 = 3'h1;
  assign T237 = T239 & T238;
  assign T238 = paddr < 32'h40008000;
  assign T239 = 32'h40000000 <= paddr;
  assign T240 = T242 ? T241 : 3'h0;
  assign T241 = 3'h7;
  assign T242 = T244 & T243;
  assign T243 = paddr < 32'h40000000;
  assign T244 = 32'h0 <= paddr;
  assign T245 = addr_ok ^ 1'h1;
  assign addr_ok = T249 | T246;
  assign T246 = T248 & T247;
  assign T247 = T366 < 33'h100000000;
  assign T366 = {1'h0, paddr};
  assign T248 = 32'h80000000 <= paddr;
  assign T249 = T253 | T250;
  assign T250 = T252 & T251;
  assign T251 = paddr < 32'h40010200;
  assign T252 = 32'h40010000 <= paddr;
  assign T253 = T257 | T254;
  assign T254 = T256 & T255;
  assign T255 = paddr < 32'h40010000;
  assign T256 = 32'h40008000 <= paddr;
  assign T257 = T261 | T258;
  assign T258 = T260 & T259;
  assign T259 = paddr < 32'h40008000;
  assign T260 = 32'h40000000 <= paddr;
  assign T261 = T263 & T262;
  assign T262 = paddr < 32'h40000000;
  assign T263 = 32'h0 <= paddr;
  assign io_resp_xcpt_st = T264;
  assign T264 = T269 | T265;
  assign T265 = tlb_hit & T266;
  assign T266 = T267 ^ 1'h1;
  assign T267 = T268 != 4'h0;
  assign T268 = w_array & tag_cam_io_hits;
  assign T269 = T270 | bad_va;
  assign T270 = T273 | T271;
  assign T271 = T272 ^ 1'h1;
  assign T272 = T216[1'h1:1'h1];
  assign T273 = addr_ok ^ 1'h1;
  assign io_resp_xcpt_ld = T274;
  assign T274 = T325 | T275;
  assign T275 = tlb_hit & T276;
  assign T276 = T277 ^ 1'h1;
  assign T277 = T278 != 4'h0;
  assign T278 = r_array & tag_cam_io_hits;
  assign r_array = priv_s ? T303 : T279;
  assign T279 = T280;
  assign T280 = {T296, T281};
  assign T281 = {ur_array_1, ur_array_0};
  assign T282 = T289 ? T283 : ur_array_0;
  assign T283 = T285 & T284;
  assign T284 = io_ptw_resp_bits_error ^ 1'h1;
  assign T285 = T287 & T286;
  assign T286 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T287 = io_ptw_resp_bits_pte_v & T288;
  assign T288 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T289 = io_ptw_resp_valid & T290;
  assign T290 = T291[1'h0:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = r_refill_waddr;
  assign T293 = T294 ? T283 : ur_array_1;
  assign T294 = io_ptw_resp_valid & T295;
  assign T295 = T291[1'h1:1'h1];
  assign T296 = {ur_array_3, ur_array_2};
  assign T297 = T298 ? T283 : ur_array_2;
  assign T298 = io_ptw_resp_valid & T299;
  assign T299 = T291[2'h2:2'h2];
  assign T300 = T301 ? T283 : ur_array_3;
  assign T301 = io_ptw_resp_valid & T302;
  assign T302 = T291[2'h3:2'h3];
  assign T303 = T304;
  assign T304 = {T318, T305};
  assign T305 = {sr_array_1, sr_array_0};
  assign T306 = T311 ? T307 : sr_array_0;
  assign T307 = T309 & T308;
  assign T308 = io_ptw_resp_bits_error ^ 1'h1;
  assign T309 = io_ptw_resp_bits_pte_v & T310;
  assign T310 = 4'h2 <= io_ptw_resp_bits_pte_typ;
  assign T311 = io_ptw_resp_valid & T312;
  assign T312 = T313[1'h0:1'h0];
  assign T313 = 1'h1 << T314;
  assign T314 = r_refill_waddr;
  assign T315 = T316 ? T307 : sr_array_1;
  assign T316 = io_ptw_resp_valid & T317;
  assign T317 = T313[1'h1:1'h1];
  assign T318 = {sr_array_3, sr_array_2};
  assign T319 = T320 ? T307 : sr_array_2;
  assign T320 = io_ptw_resp_valid & T321;
  assign T321 = T313[2'h2:2'h2];
  assign T322 = T323 ? T307 : sr_array_3;
  assign T323 = io_ptw_resp_valid & T324;
  assign T324 = T313[2'h3:2'h3];
  assign T325 = T326 | bad_va;
  assign T326 = T329 | T327;
  assign T327 = T328 ^ 1'h1;
  assign T328 = T216[1'h0:1'h0];
  assign T329 = addr_ok ^ 1'h1;
  assign io_resp_ppn = T330;
  assign T330 = vm_enabled ? T332 : T331;
  assign T331 = io_req_bits_vpn[5'h13:1'h0];
  assign T332 = T337 | T333;
  assign T333 = T336 ? T334 : 20'h0;
  assign T334 = tag_ram[2'h3];
  assign T336 = tag_cam_io_hits[2'h3:2'h3];
  assign T337 = T341 | T338;
  assign T338 = T340 ? T339 : 20'h0;
  assign T339 = tag_ram[2'h2];
  assign T340 = tag_cam_io_hits[2'h2:2'h2];
  assign T341 = T345 | T342;
  assign T342 = T344 ? T343 : 20'h0;
  assign T343 = tag_ram[2'h1];
  assign T344 = tag_cam_io_hits[1'h1:1'h1];
  assign T345 = T347 ? T346 : 20'h0;
  assign T346 = tag_ram[2'h0];
  assign T347 = tag_cam_io_hits[1'h0:1'h0];
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T348;
  assign T348 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( T152 ),
       .io_clear_mask( T128 ),
       .io_tag( T363 ),
       //.io_hit(  )
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T114 ),
       .io_write_tag( T361 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T105) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T24) begin
      R9 <= T11;
    end
    if(T40) begin
      uw_array_0 <= T32;
    end
    if(T45) begin
      uw_array_1 <= T32;
    end
    if(T49) begin
      uw_array_2 <= T32;
    end
    if(T52) begin
      uw_array_3 <= T32;
    end
    if(T64) begin
      sw_array_0 <= T58;
    end
    if(T69) begin
      sw_array_1 <= T58;
    end
    if(T73) begin
      sw_array_2 <= T58;
    end
    if(T76) begin
      sw_array_3 <= T58;
    end
    if(T84) begin
      dirty_array_0 <= io_ptw_resp_bits_pte_d;
    end
    if(T89) begin
      dirty_array_1 <= io_ptw_resp_bits_pte_d;
    end
    if(T93) begin
      dirty_array_2 <= io_ptw_resp_bits_pte_d;
    end
    if(T96) begin
      dirty_array_3 <= io_ptw_resp_bits_pte_d;
    end
    if(T105) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T126) begin
      state <= 2'h3;
    end else if(T125) begin
      state <= 2'h3;
    end else if(T124) begin
      state <= 2'h2;
    end else if(T122) begin
      state <= 2'h0;
    end else if(T105) begin
      state <= 2'h1;
    end
    if(T138) begin
      valid_array_0 <= T137;
    end
    if(T143) begin
      valid_array_1 <= T137;
    end
    if(T147) begin
      valid_array_2 <= T137;
    end
    if(T150) begin
      valid_array_3 <= T137;
    end
    if(T105) begin
      r_req_instruction <= io_req_bits_instruction;
    end
    if(T105) begin
      r_req_store <= io_req_bits_store;
    end
    if(T174) begin
      ux_array_0 <= T166;
    end
    if(T179) begin
      ux_array_1 <= T166;
    end
    if(T183) begin
      ux_array_2 <= T166;
    end
    if(T186) begin
      ux_array_3 <= T166;
    end
    if(T198) begin
      sx_array_0 <= T192;
    end
    if(T203) begin
      sx_array_1 <= T192;
    end
    if(T207) begin
      sx_array_2 <= T192;
    end
    if(T210) begin
      sx_array_3 <= T192;
    end
    if(T289) begin
      ur_array_0 <= T283;
    end
    if(T294) begin
      ur_array_1 <= T283;
    end
    if(T298) begin
      ur_array_2 <= T283;
    end
    if(T301) begin
      ur_array_3 <= T283;
    end
    if(T311) begin
      sr_array_0 <= T307;
    end
    if(T316) begin
      sr_array_1 <= T307;
    end
    if(T320) begin
      sr_array_2 <= T307;
    end
    if(T323) begin
      sr_array_3 <= T307;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_pte_ppn;
  end
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [31:0] io_enq_bits_data,
    input [127:0] io_enq_bits_datablock,
    input  io_deq_ready,
    output io_deq_valid,
    output[31:0] io_deq_bits_data,
    output[127:0] io_deq_bits_datablock,
    output io_count
);

  wire T12;
  wire[1:0] T0;
  reg  full;
  wire T13;
  wire T1;
  wire do_enq;
  wire T2;
  wire do_deq;
  wire[127:0] T3;
  wire[159:0] T4;
  reg [159:0] ram [0:0];
  wire[159:0] T5;
  wire[159:0] T6;
  wire[159:0] T7;
  wire[31:0] T8;
  wire T9;
  wire empty;
  wire T10;
  wire T11;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T12;
  assign T12 = T0[1'h0:1'h0];
  assign T0 = {full, 1'h0};
  assign T13 = reset ? 1'h0 : T1;
  assign T1 = T2 ? do_enq : full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T2 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_datablock = T3;
  assign T3 = T4[7'h7f:1'h0];
  assign T4 = ram[1'h0];
  assign T6 = T7;
  assign T7 = {io_enq_bits_data, io_enq_bits_datablock};
  assign io_deq_bits_data = T8;
  assign T8 = T4[8'h9f:8'h80];
  assign io_deq_valid = T9;
  assign T9 = empty ^ 1'h1;
  assign empty = full ^ 1'h1;
  assign io_enq_ready = T10;
  assign T10 = T11 | io_deq_ready;
  assign T11 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      full <= 1'h0;
    end else if(T2) begin
      full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T6;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data_0,
    output io_cpu_resp_bits_mask,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output io_cpu_btb_resp_bits_mask,
    output io_cpu_btb_resp_bits_bridx,
    output[38:0] io_cpu_btb_resp_bits_target,
    output[2:0] io_cpu_btb_resp_bits_entry,
    output[3:0] io_cpu_btb_resp_bits_bht_history,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input  io_cpu_btb_update_bits_prediction_bits_mask,
    input  io_cpu_btb_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [2:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_btb_update_bits_pc,
    input [38:0] io_cpu_btb_update_bits_target,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isReturn,
    input [38:0] io_cpu_btb_update_bits_br_pc,
    input  io_cpu_bht_update_valid,
    input  io_cpu_bht_update_bits_prediction_valid,
    input  io_cpu_bht_update_bits_prediction_bits_taken,
    input  io_cpu_bht_update_bits_prediction_bits_mask,
    input  io_cpu_bht_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_bht_update_bits_prediction_bits_target,
    input [2:0] io_cpu_bht_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
    input [38:0] io_cpu_bht_update_bits_pc,
    input  io_cpu_bht_update_bits_taken,
    input  io_cpu_bht_update_bits_mispredict,
    input  io_cpu_ras_update_valid,
    input  io_cpu_ras_update_bits_isCall,
    input  io_cpu_ras_update_bits_isReturn,
    input [38:0] io_cpu_ras_update_bits_returnAddr,
    input  io_cpu_ras_update_bits_prediction_valid,
    input  io_cpu_ras_update_bits_prediction_bits_taken,
    input  io_cpu_ras_update_bits_prediction_bits_mask,
    input  io_cpu_ras_update_bits_prediction_bits_bridx,
    input [38:0] io_cpu_ras_update_bits_prediction_bits_target,
    input [2:0] io_cpu_ras_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
    input [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
    input  io_cpu_invalidate,
    output[39:0] io_cpu_npc,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data
);

  wire T0;
  wire T1;
  reg  s1_same_block;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire s0_same_block;
  wire T6;
  wire[39:0] T7;
  wire[39:0] s1_pc;
  wire[39:0] T8;
  wire[39:0] T9;
  reg [39:0] s1_pc_;
  wire[39:0] T10;
  wire[39:0] T11;
  wire[39:0] npc;
  wire[39:0] T12;
  wire[39:0] predicted_npc;
  wire[39:0] ntpc;
  wire[38:0] T13;
  wire[36:0] T14;
  wire[39:0] ntpc_0;
  wire T15;
  wire T16;
  wire T17;
  wire[39:0] btbTarget;
  wire T18;
  reg [39:0] s2_pc;
  wire[39:0] T71;
  wire[39:0] T19;
  wire T20;
  wire T21;
  wire icmiss;
  wire T22;
  wire s2_resp_valid;
  reg  s2_valid;
  wire T72;
  wire T23;
  wire T24;
  wire T25;
  wire[39:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire stall;
  wire T33;
  wire T34;
  wire[27:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[11:0] T73;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[38:0] T74;
  wire T50;
  wire T51;
  wire T52;
  wire[39:0] T53;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T54;
  wire T55;
  reg [3:0] s2_btb_resp_bits_bht_history;
  wire[3:0] T56;
  reg [2:0] s2_btb_resp_bits_entry;
  wire[2:0] T57;
  reg [38:0] s2_btb_resp_bits_target;
  wire[38:0] T58;
  reg  s2_btb_resp_bits_bridx;
  wire T59;
  reg  s2_btb_resp_bits_mask;
  wire T60;
  reg  s2_btb_resp_bits_taken;
  wire T61;
  reg  s2_btb_resp_valid;
  wire T75;
  wire T62;
  reg  s2_xcpt_if;
  wire T76;
  wire T63;
  wire T77;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T78;
  wire[31:0] T66;
  wire[127:0] fetch_data;
  wire[6:0] T67;
  wire[1:0] T68;
  wire[127:0] s2_resp_data;
  wire T69;
  wire T70;
  wire btb_io_resp_valid;
  wire btb_io_resp_bits_taken;
  wire btb_io_resp_bits_mask;
  wire btb_io_resp_bits_bridx;
  wire[38:0] btb_io_resp_bits_target;
  wire[2:0] btb_io_resp_bits_entry;
  wire[3:0] btb_io_resp_bits_bht_history;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire Queue_io_deq_valid;
  wire[127:0] Queue_io_deq_bits_datablock;
  wire icache_io_resp_valid;
  wire[127:0] icache_io_resp_bits_datablock;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire tlb_io_resp_miss;
  wire[19:0] tlb_io_resp_ppn;
  wire tlb_io_resp_xcpt_if;
  wire tlb_io_ptw_req_valid;
  wire[26:0] tlb_io_ptw_req_bits_addr;
  wire[1:0] tlb_io_ptw_req_bits_prv;
  wire tlb_io_ptw_req_bits_store;
  wire tlb_io_ptw_req_bits_fetch;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    s1_same_block = {1{$random}};
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_history = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_bridx = {1{$random}};
    s2_btb_resp_bits_mask = {1{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T34 & T1;
  assign T1 = s1_same_block ^ 1'h1;
  assign T2 = io_cpu_req_valid ? 1'h0 : T3;
  assign T3 = T32 ? T4 : s1_same_block;
  assign T4 = s0_same_block & T5;
  assign T5 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T27 & T6;
  assign T6 = T26 == T7;
  assign T7 = s1_pc & 40'h10;
  assign s1_pc = ~ T8;
  assign T8 = T9 | 40'h3;
  assign T9 = ~ s1_pc_;
  assign T10 = io_cpu_req_valid ? io_cpu_req_bits_pc : T11;
  assign T11 = T32 ? npc : s1_pc_;
  assign npc = T12;
  assign T12 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : ntpc;
  assign ntpc = {T15, T13};
  assign T13 = {T14, 2'h0};
  assign T14 = ntpc_0[6'h26:2'h2];
  assign ntpc_0 = s1_pc + 40'h4;
  assign T15 = T17 & T16;
  assign T16 = ntpc_0[6'h26:6'h26];
  assign T17 = s1_pc[6'h26:6'h26];
  assign btbTarget = {T18, btb_io_resp_bits_target};
  assign T18 = btb_io_resp_bits_target[6'h26:6'h26];
  assign T71 = reset ? 40'h200 : T19;
  assign T19 = T20 ? s1_pc : s2_pc;
  assign T20 = T32 & T21;
  assign T21 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T22;
  assign T22 = s2_resp_valid ^ 1'h1;
  assign s2_resp_valid = Queue_io_deq_valid;
  assign T72 = reset ? 1'h1 : T23;
  assign T23 = io_cpu_req_valid ? 1'h0 : T24;
  assign T24 = T32 ? T25 : s2_valid;
  assign T25 = icmiss ^ 1'h1;
  assign T26 = ntpc & 40'h10;
  assign T27 = T29 & T28;
  assign T28 = btb_io_resp_bits_taken ^ 1'h1;
  assign T29 = T31 & T30;
  assign T30 = io_cpu_req_valid ^ 1'h1;
  assign T31 = icmiss ^ 1'h1;
  assign T32 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T33;
  assign T33 = io_cpu_resp_ready ^ 1'h1;
  assign T34 = stall ^ 1'h1;
  assign T35 = s1_pc >> 4'hc;
  assign T36 = T38 & T37;
  assign T37 = icmiss ^ 1'h1;
  assign T38 = stall ^ 1'h1;
  assign T39 = T41 & T40;
  assign T40 = s1_same_block ^ 1'h1;
  assign T41 = stall ^ 1'h1;
  assign T42 = T43 | io_ptw_invalidate;
  assign T43 = T44 | icmiss;
  assign T44 = T45 | tlb_io_resp_xcpt_if;
  assign T45 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T73 = io_cpu_npc[4'hb:1'h0];
  assign T46 = T48 & T47;
  assign T47 = s0_same_block ^ 1'h1;
  assign T48 = stall ^ 1'h1;
  assign T49 = io_cpu_invalidate | io_ptw_invalidate;
  assign T74 = s1_pc[6'h26:1'h0];
  assign T50 = T52 & T51;
  assign T51 = icmiss ^ 1'h1;
  assign T52 = stall ^ 1'h1;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_npc = T53;
  assign T53 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T54 = T55 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T55 = T20 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign T56 = T55 ? btb_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T57 = T55 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T58 = T55 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign T59 = T55 ? btb_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign T60 = T55 ? btb_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T61 = T55 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T75 = reset ? 1'h0 : T62;
  assign T62 = T20 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T76 = reset ? 1'h0 : T63;
  assign T63 = T20 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_mask = T77;
  assign T77 = T64[1'h0:1'h0];
  assign T64 = s2_btb_resp_valid ? T65 : 2'h3;
  assign T65 = 2'h3 & T78;
  assign T78 = {1'h0, s2_btb_resp_bits_mask};
  assign io_cpu_resp_bits_data_0 = T66;
  assign T66 = fetch_data[5'h1f:1'h0];
  assign fetch_data = s2_resp_data >> T67;
  assign T67 = T68 << 3'h5;
  assign T68 = s2_pc[2'h3:2'h2];
  assign s2_resp_data = Queue_io_deq_bits_datablock;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_valid = T69;
  assign T69 = s2_valid & T70;
  assign T70 = s2_xcpt_if | s2_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req_valid( T50 ),
       .io_req_bits_addr( T74 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_mask( btb_io_resp_bits_mask ),
       .io_resp_bits_bridx( btb_io_resp_bits_bridx ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_history( btb_io_resp_bits_bht_history ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_btb_update_valid( io_cpu_btb_update_valid ),
       .io_btb_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_btb_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_btb_update_bits_prediction_bits_mask( io_cpu_btb_update_bits_prediction_bits_mask ),
       .io_btb_update_bits_prediction_bits_bridx( io_cpu_btb_update_bits_prediction_bits_bridx ),
       .io_btb_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_btb_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_btb_update_bits_prediction_bits_bht_history( io_cpu_btb_update_bits_prediction_bits_bht_history ),
       .io_btb_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_btb_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_btb_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_btb_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_btb_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_btb_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_btb_update_bits_br_pc( io_cpu_btb_update_bits_br_pc ),
       .io_bht_update_valid( io_cpu_bht_update_valid ),
       .io_bht_update_bits_prediction_valid( io_cpu_bht_update_bits_prediction_valid ),
       .io_bht_update_bits_prediction_bits_taken( io_cpu_bht_update_bits_prediction_bits_taken ),
       .io_bht_update_bits_prediction_bits_mask( io_cpu_bht_update_bits_prediction_bits_mask ),
       .io_bht_update_bits_prediction_bits_bridx( io_cpu_bht_update_bits_prediction_bits_bridx ),
       .io_bht_update_bits_prediction_bits_target( io_cpu_bht_update_bits_prediction_bits_target ),
       .io_bht_update_bits_prediction_bits_entry( io_cpu_bht_update_bits_prediction_bits_entry ),
       .io_bht_update_bits_prediction_bits_bht_history( io_cpu_bht_update_bits_prediction_bits_bht_history ),
       .io_bht_update_bits_prediction_bits_bht_value( io_cpu_bht_update_bits_prediction_bits_bht_value ),
       .io_bht_update_bits_pc( io_cpu_bht_update_bits_pc ),
       .io_bht_update_bits_taken( io_cpu_bht_update_bits_taken ),
       .io_bht_update_bits_mispredict( io_cpu_bht_update_bits_mispredict ),
       .io_ras_update_valid( io_cpu_ras_update_valid ),
       .io_ras_update_bits_isCall( io_cpu_ras_update_bits_isCall ),
       .io_ras_update_bits_isReturn( io_cpu_ras_update_bits_isReturn ),
       .io_ras_update_bits_returnAddr( io_cpu_ras_update_bits_returnAddr ),
       .io_ras_update_bits_prediction_valid( io_cpu_ras_update_bits_prediction_valid ),
       .io_ras_update_bits_prediction_bits_taken( io_cpu_ras_update_bits_prediction_bits_taken ),
       .io_ras_update_bits_prediction_bits_mask( io_cpu_ras_update_bits_prediction_bits_mask ),
       .io_ras_update_bits_prediction_bits_bridx( io_cpu_ras_update_bits_prediction_bits_bridx ),
       .io_ras_update_bits_prediction_bits_target( io_cpu_ras_update_bits_prediction_bits_target ),
       .io_ras_update_bits_prediction_bits_entry( io_cpu_ras_update_bits_prediction_bits_entry ),
       .io_ras_update_bits_prediction_bits_bht_history( io_cpu_ras_update_bits_prediction_bits_bht_history ),
       .io_ras_update_bits_prediction_bits_bht_value( io_cpu_ras_update_bits_prediction_bits_bht_value ),
       .io_invalidate( T49 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T46 ),
       .io_req_bits_idx( T73 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T42 ),
       .io_resp_ready( T39 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T36 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T35 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_req_bits_store( 1'h0 ),
       .io_resp_miss( tlb_io_resp_miss ),
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( tlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( tlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( tlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( tlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  Queue_8 Queue(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( icache_io_resp_valid ),
       //.io_enq_bits_data(  )
       .io_enq_bits_datablock( icache_io_resp_bits_datablock ),
       .io_deq_ready( T0 ),
       .io_deq_valid( Queue_io_deq_valid ),
       //.io_deq_bits_data(  )
       .io_deq_bits_datablock( Queue_io_deq_bits_datablock )
       //.io_count(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign Queue.io_enq_bits_data = {1{$random}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T32) begin
      s1_same_block <= T4;
    end
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T32) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 40'h200;
    end else if(T20) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T32) begin
      s2_valid <= T25;
    end
    if(T55) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T55) begin
      s2_btb_resp_bits_bht_history <= btb_io_resp_bits_bht_history;
    end
    if(T55) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T55) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T55) begin
      s2_btb_resp_bits_bridx <= btb_io_resp_bits_bridx;
    end
    if(T55) begin
      s2_btb_resp_bits_mask <= btb_io_resp_bits_mask;
    end
    if(T55) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T20) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T20) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [1:0] io_req_bits_addr_beat,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_client_xact_id,
    input  io_req_bits_voluntary,
    input [2:0] io_req_bits_r_type,
    input [127:0] io_req_bits_data,
    input  io_req_bits_way_en,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[1:0] io_release_bits_addr_beat,
    output[25:0] io_release_bits_addr_block,
    output[1:0] io_release_bits_client_xact_id,
    output io_release_bits_voluntary,
    output[2:0] io_release_bits_r_type,
    output[127:0] io_release_bits_data
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg  req_voluntary;
  wire T2;
  reg [1:0] req_client_xact_id;
  wire[1:0] T3;
  reg [25:0] req_addr_block;
  wire[25:0] T4;
  reg [1:0] beat_cnt;
  wire[1:0] T40;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  reg  r2_data_req_fired;
  wire T41;
  wire T9;
  wire T10;
  reg  r1_data_req_fired;
  wire T42;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  reg  active;
  wire T43;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [2:0] data_req_cnt;
  wire[2:0] T44;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire[2:0] T45;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire[11:0] T33;
  wire[7:0] T34;
  wire[1:0] T35;
  wire[5:0] req_idx;
  reg  req_way_en;
  wire T36;
  wire fire;
  wire T37;
  wire[19:0] T38;
  wire T39;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    req_voluntary = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr_block = {1{$random}};
    beat_cnt = {1{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    data_req_cnt = {1{$random}};
    req_way_en = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_release_bits_data = io_data_resp;
  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_voluntary = req_voluntary;
  assign T2 = T1 ? io_req_bits_voluntary : req_voluntary;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T3 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr_block = req_addr_block;
  assign T4 = T1 ? io_req_bits_addr_block : req_addr_block;
  assign io_release_bits_addr_beat = beat_cnt;
  assign T40 = reset ? 2'h0 : T5;
  assign T5 = T7 ? T6 : beat_cnt;
  assign T6 = beat_cnt + 2'h1;
  assign T7 = io_release_ready & io_release_valid;
  assign io_release_valid = T8;
  assign T8 = active & r2_data_req_fired;
  assign T41 = reset ? 1'h0 : T9;
  assign T9 = T18 ? 1'h0 : T10;
  assign T10 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T42 = reset ? 1'h0 : T11;
  assign T11 = T18 ? 1'h0 : T12;
  assign T12 = T14 ? 1'h1 : T13;
  assign T13 = active ? 1'h0 : r1_data_req_fired;
  assign T14 = active & T15;
  assign T15 = T17 & T16;
  assign T16 = io_meta_read_ready & io_meta_read_valid;
  assign T17 = io_data_req_ready & io_data_req_valid;
  assign T18 = T8 & T19;
  assign T19 = io_release_ready ^ 1'h1;
  assign T43 = reset ? 1'h0 : T20;
  assign T20 = T1 ? 1'h1 : T21;
  assign T21 = T31 ? T22 : active;
  assign T22 = T24 | T23;
  assign T23 = io_release_ready ^ 1'h1;
  assign T24 = data_req_cnt < 3'h4;
  assign T44 = reset ? 3'h0 : T25;
  assign T25 = T1 ? 3'h0 : T26;
  assign T26 = T18 ? T29 : T27;
  assign T27 = T14 ? T28 : data_req_cnt;
  assign T28 = data_req_cnt + 3'h1;
  assign T29 = data_req_cnt - T45;
  assign T45 = {1'h0, T30};
  assign T30 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign T31 = T8 & T32;
  assign T32 = r1_data_req_fired ^ 1'h1;
  assign io_data_req_bits_addr = T33;
  assign T33 = T34 << 3'h4;
  assign T34 = {req_idx, T35};
  assign T35 = data_req_cnt[1'h1:1'h0];
  assign req_idx = req_addr_block[3'h5:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T36 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T37;
  assign T37 = data_req_cnt < 3'h4;
  assign io_meta_read_bits_tag = T38;
  assign T38 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T39;
  assign T39 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T1) begin
      req_voluntary <= io_req_bits_voluntary;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_addr_block <= io_req_bits_addr_block;
    end
    if(reset) begin
      beat_cnt <= 2'h0;
    end else if(T7) begin
      beat_cnt <= T6;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(T18) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T18) begin
      r1_data_req_fired <= 1'h0;
    end else if(T14) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T31) begin
      active <= T22;
    end
    if(reset) begin
      data_req_cnt <= 3'h0;
    end else if(T1) begin
      data_req_cnt <= 3'h0;
    end else if(T18) begin
      data_req_cnt <= T29;
    end else if(T14) begin
      data_req_cnt <= T28;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr_block,
    input [1:0] io_req_bits_p_type,
    //input [1:0] io_req_bits_client_xact_id
    input  io_rep_ready,
    output io_rep_valid,
    output[1:0] io_rep_bits_addr_beat,
    output[25:0] io_rep_bits_addr_block,
    output[1:0] io_rep_bits_client_xact_id,
    output io_rep_bits_voluntary,
    output[2:0] io_rep_bits_r_type,
    output[127:0] io_rep_bits_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output io_wb_req_bits_way_en,
    input  io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_block_state_state
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg  way_en;
  wire T10;
  wire T11;
  reg [3:0] state;
  wire[3:0] T68;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire[3:0] T20;
  wire[3:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[3:0] T27;
  wire T28;
  wire T29;
  reg [1:0] old_coh_state;
  wire[1:0] T30;
  wire tag_matches;
  wire T31;
  wire[3:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire[127:0] reply_data;
  wire[2:0] reply_r_type;
  wire[2:0] T39;
  wire[2:0] T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] miss_coh_state;
  wire T45;
  reg [1:0] req_p_type;
  wire[1:0] T46;
  wire[2:0] T47;
  wire T48;
  wire T49;
  wire[2:0] T50;
  wire T51;
  wire T52;
  wire reply_voluntary;
  wire[1:0] reply_client_xact_id;
  wire[25:0] reply_addr_block;
  reg [25:0] req_addr_block;
  wire[25:0] T53;
  wire[1:0] reply_addr_beat;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[19:0] T62;
  wire[5:0] T69;
  wire T63;
  wire[19:0] T64;
  wire[5:0] T70;
  wire T65;
  wire T66;
  wire T67;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    way_en = {1{$random}};
    state = {1{$random}};
    old_coh_state = {1{$random}};
    req_p_type = {1{$random}};
    req_addr_block = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T9 | T3;
  assign T3 = T4 ^ 1'h1;
  assign T4 = T6 | T5;
  assign T5 = 3'h2 == io_rep_bits_r_type;
  assign T6 = T8 | T7;
  assign T7 = 3'h1 == io_rep_bits_r_type;
  assign T8 = 3'h0 == io_rep_bits_r_type;
  assign T9 = io_rep_valid ^ 1'h1;
  assign io_wb_req_bits_way_en = way_en;
  assign T10 = T11 ? io_way_en : way_en;
  assign T11 = state == 4'h3;
  assign T68 = reset ? 4'h0 : T12;
  assign T12 = T38 ? 4'h0 : T13;
  assign T13 = T36 ? 4'h8 : T14;
  assign T14 = T35 ? 4'h7 : T15;
  assign T15 = T33 ? T32 : T16;
  assign T16 = T31 ? T27 : T17;
  assign T17 = T25 ? 4'h1 : T18;
  assign T18 = T11 ? 4'h4 : T19;
  assign T19 = T24 ? 4'h3 : T20;
  assign T20 = T23 ? 4'h2 : T21;
  assign T21 = T22 ? 4'h1 : state;
  assign T22 = io_req_ready & io_req_valid;
  assign T23 = io_meta_read_ready & io_meta_read_valid;
  assign T24 = state == 4'h2;
  assign T25 = T11 & T26;
  assign T26 = io_mshr_rdy ^ 1'h1;
  assign T27 = T28 ? 4'h6 : 4'h5;
  assign T28 = tag_matches & T29;
  assign T29 = 2'h3 == old_coh_state;
  assign T30 = T11 ? io_block_state_state : old_coh_state;
  assign tag_matches = way_en != 1'h0;
  assign T31 = state == 4'h4;
  assign T32 = tag_matches ? 4'h8 : 4'h0;
  assign T33 = T34 & io_rep_ready;
  assign T34 = state == 4'h5;
  assign T35 = io_wb_req_ready & io_wb_req_valid;
  assign T36 = T37 & io_wb_req_ready;
  assign T37 = state == 4'h7;
  assign T38 = io_meta_write_ready & io_meta_write_valid;
  assign io_wb_req_bits_data = reply_data;
  assign reply_data = 128'h0;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign reply_r_type = T39;
  assign T39 = T52 ? T50 : T40;
  assign T40 = T49 ? T47 : T41;
  assign T41 = T45 ? T42 : 3'h3;
  assign T42 = T43 ? 3'h2 : 3'h5;
  assign T43 = 2'h3 == T44;
  assign T44 = tag_matches ? old_coh_state : miss_coh_state;
  assign miss_coh_state = 2'h0;
  assign T45 = req_p_type == 2'h2;
  assign T46 = T22 ? io_req_bits_p_type : req_p_type;
  assign T47 = T48 ? 3'h1 : 3'h4;
  assign T48 = 2'h3 == T44;
  assign T49 = req_p_type == 2'h1;
  assign T50 = T51 ? 3'h0 : 3'h3;
  assign T51 = 2'h3 == T44;
  assign T52 = req_p_type == 2'h0;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign reply_voluntary = 1'h0;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign reply_client_xact_id = 2'h0;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign reply_addr_block = req_addr_block;
  assign T53 = T22 ? io_req_bits_addr_block : req_addr_block;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign reply_addr_beat = 2'h0;
  assign io_wb_req_valid = T54;
  assign T54 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T55;
  assign T55 = T56;
  assign T56 = T61 ? 2'h0 : T57;
  assign T57 = T60 ? 2'h1 : T58;
  assign T58 = T59 ? old_coh_state : old_coh_state;
  assign T59 = req_p_type == 2'h2;
  assign T60 = req_p_type == 2'h1;
  assign T61 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T62;
  assign T62 = req_addr_block >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T69;
  assign T69 = req_addr_block[3'h5:1'h0];
  assign io_meta_write_valid = T63;
  assign T63 = state == 4'h8;
  assign io_meta_read_bits_tag = T64;
  assign T64 = req_addr_block >> 3'h6;
  assign io_meta_read_bits_idx = T70;
  assign T70 = req_addr_block[3'h5:1'h0];
  assign io_meta_read_valid = T65;
  assign T65 = state == 4'h1;
  assign io_rep_bits_data = reply_data;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_valid = T66;
  assign T66 = state == 4'h5;
  assign io_req_ready = T67;
  assign T67 = state == 4'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "ProbeUnit should not send releases with data");
    $finish;
  end
// synthesis translate_on
`endif
    if(T11) begin
      way_en <= io_way_en;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T38) begin
      state <= 4'h0;
    end else if(T36) begin
      state <= 4'h8;
    end else if(T35) begin
      state <= 4'h7;
    end else if(T33) begin
      state <= T32;
    end else if(T31) begin
      state <= T27;
    end else if(T25) begin
      state <= 4'h1;
    end else if(T11) begin
      state <= 4'h4;
    end else if(T24) begin
      state <= 4'h3;
    end else if(T23) begin
      state <= 4'h2;
    end else if(T22) begin
      state <= 4'h1;
    end
    if(T11) begin
      old_coh_state <= io_block_state_state;
    end
    if(T22) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(T22) begin
      req_addr_block <= io_req_bits_addr_block;
    end
  end
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[19:0] T0;
  wire T1;
  wire[5:0] T2;
  wire T3;
  wire T4;
  wire T5;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T0;
  assign T0 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T1 = chosen;
  assign io_out_bits_idx = T2;
  assign T2 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T3;
  assign T3 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T4;
  assign T4 = T5 & io_out_ready;
  assign T5 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[1:0] T0;
  wire T1;
  wire[19:0] T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T0;
  assign T0 = T1 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T1 = chosen;
  assign io_out_bits_data_tag = T2;
  assign T2 = T1 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T3;
  assign T3 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T4;
  assign T4 = T1 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module LockingArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [25:0] io_in_2_bits_addr_block,
    input [1:0] io_in_2_bits_client_xact_id,
    input [1:0] io_in_2_bits_addr_beat,
    input  io_in_2_bits_is_builtin_type,
    input [2:0] io_in_2_bits_a_type,
    input [16:0] io_in_2_bits_union,
    input [127:0] io_in_2_bits_data,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input [1:0] io_in_1_bits_addr_beat,
    input  io_in_1_bits_is_builtin_type,
    input [2:0] io_in_1_bits_a_type,
    input [16:0] io_in_1_bits_union,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input [1:0] io_in_0_bits_addr_beat,
    input  io_in_0_bits_is_builtin_type,
    input [2:0] io_in_0_bits_a_type,
    input [16:0] io_in_0_bits_union,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output[1:0] io_out_bits_addr_beat,
    output io_out_bits_is_builtin_type,
    output[2:0] io_out_bits_a_type,
    output[16:0] io_out_bits_union,
    output[127:0] io_out_bits_data,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  reg [1:0] lockIdx;
  wire[1:0] T65;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T66;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T67;
  wire[1:0] T19;
  wire[127:0] T20;
  wire[127:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire T27;
  wire T28;
  wire[2:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  wire[25:0] T45;
  wire[25:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid ? 2'h0 : T1;
  assign T1 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T65 = reset ? 2'h2 : T2;
  assign T2 = T7 ? T3 : lockIdx;
  assign T3 = T6 ? 2'h0 : T4;
  assign T4 = T5 ? 2'h1 : 2'h2;
  assign T5 = io_in_1_ready & io_in_1_valid;
  assign T6 = io_in_0_ready & io_in_0_valid;
  assign T7 = T9 & T8;
  assign T8 = locked ^ 1'h1;
  assign T9 = T12 & T10;
  assign T10 = io_out_bits_is_builtin_type & T11;
  assign T11 = 3'h3 == io_out_bits_a_type;
  assign T12 = io_out_ready & io_out_valid;
  assign T66 = reset ? 1'h0 : T13;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = T7 ? 1'h1 : locked;
  assign T15 = T12 & T16;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T67 = reset ? 2'h0 : T19;
  assign T19 = T9 ? T17 : R18;
  assign io_out_bits_data = T20;
  assign T20 = T24 ? io_in_2_bits_data : T21;
  assign T21 = T22 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T22 = T23[1'h0:1'h0];
  assign T23 = chosen;
  assign T24 = T23[1'h1:1'h1];
  assign io_out_bits_union = T25;
  assign T25 = T28 ? io_in_2_bits_union : T26;
  assign T26 = T27 ? io_in_1_bits_union : io_in_0_bits_union;
  assign T27 = T23[1'h0:1'h0];
  assign T28 = T23[1'h1:1'h1];
  assign io_out_bits_a_type = T29;
  assign T29 = T32 ? io_in_2_bits_a_type : T30;
  assign T30 = T31 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign T31 = T23[1'h0:1'h0];
  assign T32 = T23[1'h1:1'h1];
  assign io_out_bits_is_builtin_type = T33;
  assign T33 = T36 ? io_in_2_bits_is_builtin_type : T34;
  assign T34 = T35 ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign T35 = T23[1'h0:1'h0];
  assign T36 = T23[1'h1:1'h1];
  assign io_out_bits_addr_beat = T37;
  assign T37 = T40 ? io_in_2_bits_addr_beat : T38;
  assign T38 = T39 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign T39 = T23[1'h0:1'h0];
  assign T40 = T23[1'h1:1'h1];
  assign io_out_bits_client_xact_id = T41;
  assign T41 = T44 ? io_in_2_bits_client_xact_id : T42;
  assign T42 = T43 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign T43 = T23[1'h0:1'h0];
  assign T44 = T23[1'h1:1'h1];
  assign io_out_bits_addr_block = T45;
  assign T45 = T48 ? io_in_2_bits_addr_block : T46;
  assign T46 = T47 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign T47 = T23[1'h0:1'h0];
  assign T48 = T23[1'h1:1'h1];
  assign io_out_valid = T49;
  assign T49 = T52 ? io_in_2_valid : T50;
  assign T50 = T51 ? io_in_1_valid : io_in_0_valid;
  assign T51 = T23[1'h0:1'h0];
  assign T52 = T23[1'h1:1'h1];
  assign io_in_0_ready = T53;
  assign T53 = T54 & io_out_ready;
  assign T54 = locked ? T55 : 1'h1;
  assign T55 = lockIdx == 2'h0;
  assign io_in_1_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = locked ? T59 : T58;
  assign T58 = io_in_0_valid ^ 1'h1;
  assign T59 = lockIdx == 2'h1;
  assign io_in_2_ready = T60;
  assign T60 = T61 & io_out_ready;
  assign T61 = locked ? T64 : T62;
  assign T62 = T63 ^ 1'h1;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign T64 = lockIdx == 2'h2;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 2'h2;
    end else if(T7) begin
      lockIdx <= T3;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h0;
    end else if(T7) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T9) begin
      R18 <= T17;
    end
  end
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_voluntary,
    input [2:0] io_in_1_bits_r_type,
    input [127:0] io_in_1_bits_data,
    input  io_in_1_bits_way_en,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_voluntary,
    input [2:0] io_in_0_bits_r_type,
    input [127:0] io_in_0_bits_data,
    input  io_in_0_bits_way_en,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output io_out_bits_voluntary,
    output[2:0] io_out_bits_r_type,
    output[127:0] io_out_bits_data,
    output io_out_bits_way_en,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire[127:0] T2;
  wire[2:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[25:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_way_en = T0;
  assign T0 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T1 = chosen;
  assign io_out_bits_data = T2;
  assign T2 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_r_type = T3;
  assign T3 = T1 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_voluntary = T4;
  assign T4 = T1 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T1 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T6;
  assign T6 = T1 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T7;
  assign T7 = T1 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_7(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [39:0] io_in_1_bits_addr,
    input [8:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_kill,
    input  io_in_1_bits_phys,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_kill,
    input  io_in_0_bits_phys,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output io_out_bits_kill,
    output io_out_bits_phys,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[4:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire[2:0] T4;
  wire[4:0] T5;
  wire[8:0] T6;
  wire[39:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T0;
  assign T0 = T1 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T1 = chosen;
  assign io_out_bits_phys = T2;
  assign T2 = T1 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_kill = T3;
  assign T3 = T1 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_bits_typ = T4;
  assign T4 = T1 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_cmd = T5;
  assign T5 = T1 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T6;
  assign T6 = T1 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_addr = T7;
  assign T7 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_8(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits = T0;
  assign T0 = T1 ? io_in_1_bits : io_in_0_bits;
  assign T1 = chosen;
  assign io_out_valid = T2;
  assign T2 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T3;
  assign T3 = T4 & io_out_ready;
  assign T4 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [39:0] io_enq_bits_addr,
    input [8:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_kill,
    input  io_enq_bits_phys,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[39:0] io_deq_bits_addr,
    output[8:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_kill,
    output io_deq_bits_phys,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T29;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T30;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T31;
  wire T8;
  wire T9;
  wire[4:0] T10;
  wire[63:0] T11;
  reg [63:0] ram [15:0];
  wire[63:0] T12;
  wire[63:0] T13;
  wire[63:0] T14;
  wire[9:0] T15;
  wire[5:0] T16;
  wire[3:0] T17;
  wire[53:0] T18;
  wire[13:0] T19;
  wire T20;
  wire T21;
  wire[2:0] T22;
  wire[4:0] T23;
  wire[8:0] T24;
  wire[39:0] T25;
  wire T26;
  wire empty;
  wire T27;
  wire T28;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T29 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T30 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T31 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T10;
  assign T10 = T11[3'h4:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {io_enq_bits_phys, io_enq_bits_sdq_id};
  assign T17 = {io_enq_bits_typ, io_enq_bits_kill};
  assign T18 = {io_enq_bits_addr, T19};
  assign T19 = {io_enq_bits_tag, io_enq_bits_cmd};
  assign io_deq_bits_phys = T20;
  assign T20 = T11[3'h5:3'h5];
  assign io_deq_bits_kill = T21;
  assign T21 = T11[3'h6:3'h6];
  assign io_deq_bits_typ = T22;
  assign T22 = T11[4'h9:3'h7];
  assign io_deq_bits_cmd = T23;
  assign T23 = T11[4'he:4'ha];
  assign io_deq_bits_tag = T24;
  assign T24 = T11[5'h17:4'hf];
  assign io_deq_bits_addr = T25;
  assign T25 = T11[6'h3f:5'h18];
  assign io_deq_valid = T26;
  assign T26 = empty ^ 1'h1;
  assign empty = ptr_match & T27;
  assign T27 = maybe_full ^ 1'h1;
  assign io_enq_ready = T28;
  assign T28 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  req_way_en;
  wire T133;
  wire[127:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire T139;
  wire[1:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_voluntary = T139;
  assign T139 = 1'h1;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 2'h0;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3:2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 2'h0;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_15 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [4:0] io_req_bits_sdq_id,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output io_wb_req_bits_way_en,
    output io_probe_rdy
);

  wire T0;
  wire T1;
  wire T2;
  reg [3:0] state;
  wire[3:0] T216;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  wire refill_count_done;
  wire T22;
  reg [1:0] refill_cnt;
  wire[1:0] T217;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire gnt_multi_data;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire sec_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire cmd_requires_second_acquire;
  wire T80;
  wire T81;
  wire T82;
  reg [4:0] req_cmd;
  wire[4:0] T83;
  wire[4:0] T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire idx_match;
  wire[5:0] T115;
  wire[5:0] req_idx;
  reg [39:0] req_addr;
  wire[39:0] T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  reg [1:0] meta_hazard;
  wire[1:0] T218;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  req_way_en;
  wire T133;
  wire[127:0] T134;
  wire[2:0] T135;
  wire[2:0] T136;
  wire T137;
  reg [1:0] req_old_meta_coh_state;
  wire[1:0] T138;
  wire T139;
  wire[1:0] T140;
  wire[25:0] T141;
  wire[25:0] T142;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T143;
  wire[1:0] T144;
  wire T145;
  wire[4:0] T146;
  wire[39:0] T219;
  wire[31:0] T147;
  wire[31:0] T148;
  wire[11:0] T149;
  wire[5:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  reg [1:0] new_coh_state_state;
  wire[1:0] T154;
  wire[1:0] T220;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[1:0] coh_on_grant_state;
  wire[1:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[1:0] coh_on_hit_state;
  wire[1:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[11:0] T187;
  wire[7:0] T188;
  wire[127:0] T189;
  wire[16:0] T190;
  wire[16:0] T221;
  wire[5:0] T191;
  wire[2:0] T192;
  wire[2:0] T222;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire[25:0] T207;
  wire[25:0] T208;
  wire[25:0] T209;
  wire T210;
  wire[19:0] T223;
  wire[27:0] T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire rpq_io_enq_ready;
  wire rpq_io_deq_valid;
  wire[39:0] rpq_io_deq_bits_addr;
  wire[8:0] rpq_io_deq_bits_tag;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire[4:0] rpq_io_deq_bits_sdq_id;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_cnt = {1{$random}};
    req_cmd = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_coh_state = {1{$random}};
    req_old_meta_tag = {1{$random}};
    new_coh_state_state = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T69 ? 1'h0 : T1;
  assign T1 = T67 | T2;
  assign T2 = state == 4'h0;
  assign T216 = reset ? 4'h0 : T3;
  assign T3 = T65 ? T63 : T4;
  assign T4 = T61 ? 4'h4 : T5;
  assign T5 = T38 ? 4'h6 : T6;
  assign T6 = T37 ? 4'h2 : T7;
  assign T7 = T35 ? 4'h3 : T8;
  assign T8 = T33 ? 4'h4 : T9;
  assign T9 = T32 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T31 & refill_done;
  assign refill_done = io_mem_grant_valid & T21;
  assign T21 = T30 | refill_count_done;
  assign refill_count_done = T25 & T22;
  assign T22 = refill_cnt == 2'h3;
  assign T217 = reset ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_cnt;
  assign T24 = refill_cnt + 2'h1;
  assign T25 = io_mem_grant_valid & gnt_multi_data;
  assign gnt_multi_data = io_mem_grant_bits_is_builtin_type ? T29 : T26;
  assign T26 = T28 | T27;
  assign T27 = 4'h1 == io_mem_grant_bits_g_type;
  assign T28 = 4'h0 == io_mem_grant_bits_g_type;
  assign T29 = 4'h5 == io_mem_grant_bits_g_type;
  assign T30 = gnt_multi_data ^ 1'h1;
  assign T31 = state == 4'h5;
  assign T32 = io_mem_req_ready & io_mem_req_valid;
  assign T33 = T34 & io_meta_write_ready;
  assign T34 = state == 4'h3;
  assign T35 = T36 & io_mem_grant_valid;
  assign T36 = state == 4'h2;
  assign T37 = io_wb_req_ready & io_wb_req_valid;
  assign T38 = T59 & T39;
  assign T39 = T48 ? T45 : T40;
  assign T40 = T42 | T41;
  assign T41 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T42 = T44 | T43;
  assign T43 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T44 = 2'h1 == io_req_bits_old_meta_coh_state;
  assign T45 = T47 | T46;
  assign T46 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T47 = 2'h2 == io_req_bits_old_meta_coh_state;
  assign T48 = T50 | T49;
  assign T49 = io_req_bits_cmd == 5'h6;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h3;
  assign T52 = T56 | T53;
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h4;
  assign T55 = io_req_bits_cmd[2'h3:2'h3];
  assign T56 = T58 | T57;
  assign T57 = io_req_bits_cmd == 5'h7;
  assign T58 = io_req_bits_cmd == 5'h1;
  assign T59 = T60 & io_req_bits_tag_match;
  assign T60 = io_req_pri_val & io_req_pri_rdy;
  assign T61 = T59 & T62;
  assign T62 = T39 ^ 1'h1;
  assign T63 = T64 ? 4'h1 : 4'h3;
  assign T64 = 2'h3 == io_req_bits_old_meta_coh_state;
  assign T65 = T60 & T66;
  assign T66 = io_req_bits_tag_match ^ 1'h1;
  assign T67 = io_replay_ready & T68;
  assign T68 = state == 4'h8;
  assign T69 = io_meta_read_ready ^ 1'h1;
  assign T70 = T75 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T74 | T73;
  assign T73 = io_req_bits_cmd == 5'h3;
  assign T74 = io_req_bits_cmd == 5'h2;
  assign T75 = T117 | T76;
  assign T76 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T77;
  assign T77 = T110 | T78;
  assign T78 = T107 & T79;
  assign T79 = cmd_requires_second_acquire ^ 1'h1;
  assign cmd_requires_second_acquire = T96 & T80;
  assign T80 = T81 ^ 1'h1;
  assign T81 = T87 | T82;
  assign T82 = req_cmd == 5'h6;
  assign T83 = T60 ? io_req_bits_cmd : T84;
  assign T84 = T85 ? io_req_bits_cmd : req_cmd;
  assign T85 = T86 & cmd_requires_second_acquire;
  assign T86 = io_req_sec_val & io_req_sec_rdy;
  assign T87 = T89 | T88;
  assign T88 = req_cmd == 5'h3;
  assign T89 = T93 | T90;
  assign T90 = T92 | T91;
  assign T91 = req_cmd == 5'h4;
  assign T92 = req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = req_cmd == 5'h7;
  assign T95 = req_cmd == 5'h1;
  assign T96 = T98 | T97;
  assign T97 = io_req_bits_cmd == 5'h6;
  assign T98 = T100 | T99;
  assign T99 = io_req_bits_cmd == 5'h3;
  assign T100 = T104 | T101;
  assign T101 = T103 | T102;
  assign T102 = io_req_bits_cmd == 5'h4;
  assign T103 = io_req_bits_cmd[2'h3:2'h3];
  assign T104 = T106 | T105;
  assign T105 = io_req_bits_cmd == 5'h7;
  assign T106 = io_req_bits_cmd == 5'h1;
  assign T107 = T109 | T108;
  assign T108 = 4'h5 == state;
  assign T109 = 4'h4 == state;
  assign T110 = T112 | T111;
  assign T111 = 4'h3 == state;
  assign T112 = T114 | T113;
  assign T113 = 4'h2 == state;
  assign T114 = 4'h1 == state;
  assign idx_match = req_idx == T115;
  assign T115 = io_req_bits_addr[4'hb:3'h6];
  assign req_idx = req_addr[4'hb:3'h6];
  assign T116 = T60 ? io_req_bits_addr : req_addr;
  assign T117 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T118;
  assign T118 = T132 | T119;
  assign T119 = T126 & T120;
  assign T120 = meta_hazard == 2'h0;
  assign T218 = reset ? 2'h0 : T121;
  assign T121 = T125 ? 2'h1 : T122;
  assign T122 = T124 ? T123 : meta_hazard;
  assign T123 = meta_hazard + 2'h1;
  assign T124 = meta_hazard != 2'h0;
  assign T125 = io_meta_write_ready & io_meta_write_valid;
  assign T126 = T127 ^ 1'h1;
  assign T127 = T129 | T128;
  assign T128 = 4'h3 == state;
  assign T129 = T131 | T130;
  assign T130 = 4'h2 == state;
  assign T131 = 4'h1 == state;
  assign T132 = idx_match ^ 1'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T133 = T60 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_data = T134;
  assign T134 = 128'h0;
  assign io_wb_req_bits_r_type = T135;
  assign T135 = T136;
  assign T136 = T137 ? 3'h0 : 3'h3;
  assign T137 = 2'h3 == req_old_meta_coh_state;
  assign T138 = T60 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign io_wb_req_bits_voluntary = T139;
  assign T139 = 1'h1;
  assign io_wb_req_bits_client_xact_id = T140;
  assign T140 = 2'h1;
  assign io_wb_req_bits_addr_block = T141;
  assign T141 = T142;
  assign T142 = {req_old_meta_tag, req_idx};
  assign T143 = T60 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_bits_addr_beat = T144;
  assign T144 = 2'h0;
  assign io_wb_req_valid = T145;
  assign T145 = state == 4'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_cmd = T146;
  assign T146 = T69 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_addr = T219;
  assign T219 = {8'h0, T147};
  assign T147 = T148;
  assign T148 = {io_tag, T149};
  assign T149 = {req_idx, T150};
  assign T150 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_valid = T151;
  assign T151 = T152 & rpq_io_deq_valid;
  assign T152 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T153;
  assign T153 = T182 ? T181 : new_coh_state_state;
  assign T154 = 2'h0;
  assign T220 = reset ? T154 : T155;
  assign T155 = T38 ? coh_on_hit_state : T156;
  assign T156 = T172 ? coh_on_grant_state : new_coh_state_state;
  assign coh_on_grant_state = T157;
  assign T157 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T158;
  assign T158 = T171 ? 2'h1 : T159;
  assign T159 = T170 ? T162 : T160;
  assign T160 = T161 ? 2'h3 : 2'h0;
  assign T161 = io_mem_grant_bits_g_type == 4'h2;
  assign T162 = T163 ? 2'h3 : 2'h2;
  assign T163 = T167 | T164;
  assign T164 = T166 | T165;
  assign T165 = req_cmd == 5'h4;
  assign T166 = req_cmd[2'h3:2'h3];
  assign T167 = T169 | T168;
  assign T168 = req_cmd == 5'h7;
  assign T169 = req_cmd == 5'h1;
  assign T170 = io_mem_grant_bits_g_type == 4'h1;
  assign T171 = io_mem_grant_bits_g_type == 4'h0;
  assign T172 = T31 & io_mem_grant_valid;
  assign coh_on_hit_state = T173;
  assign T173 = T174 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T174 = T178 | T175;
  assign T175 = T177 | T176;
  assign T176 = io_req_bits_cmd == 5'h4;
  assign T177 = io_req_bits_cmd[2'h3:2'h3];
  assign T178 = T180 | T179;
  assign T179 = io_req_bits_cmd == 5'h7;
  assign T180 = io_req_bits_cmd == 5'h1;
  assign T181 = 2'h0;
  assign T182 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_valid = T183;
  assign T183 = T185 | T184;
  assign T184 = state == 4'h3;
  assign T185 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = T186;
  assign T186 = state == 4'h8;
  assign io_refill_addr = T187;
  assign T187 = T188 << 3'h4;
  assign T188 = {req_idx, refill_cnt};
  assign io_refill_way_en = req_way_en;
  assign io_mem_req_bits_data = T189;
  assign T189 = 128'h0;
  assign io_mem_req_bits_union = T190;
  assign T190 = T221;
  assign T221 = {11'h0, T191};
  assign T191 = {req_cmd, 1'h1};
  assign io_mem_req_bits_a_type = T192;
  assign T192 = T222;
  assign T222 = {2'h0, T193};
  assign T193 = T195 | T194;
  assign T194 = req_cmd == 5'h6;
  assign T195 = T197 | T196;
  assign T196 = req_cmd == 5'h3;
  assign T197 = T201 | T198;
  assign T198 = T200 | T199;
  assign T199 = req_cmd == 5'h4;
  assign T200 = req_cmd[2'h3:2'h3];
  assign T201 = T203 | T202;
  assign T202 = req_cmd == 5'h7;
  assign T203 = req_cmd == 5'h1;
  assign io_mem_req_bits_is_builtin_type = T204;
  assign T204 = 1'h0;
  assign io_mem_req_bits_addr_beat = T205;
  assign T205 = 2'h0;
  assign io_mem_req_bits_client_xact_id = T206;
  assign T206 = 2'h1;
  assign io_mem_req_bits_addr_block = T207;
  assign T207 = T208;
  assign T208 = T209;
  assign T209 = {io_tag, req_idx};
  assign io_mem_req_valid = T210;
  assign T210 = state == 4'h4;
  assign io_tag = T223;
  assign T223 = T211[5'h13:1'h0];
  assign T211 = req_addr >> 4'hc;
  assign io_idx_match = T212;
  assign T212 = T213 & idx_match;
  assign T213 = state != 4'h0;
  assign io_req_sec_rdy = T214;
  assign T214 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T215;
  assign T215 = state == 4'h0;
  Queue_15 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T70 ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_sdq_id( io_req_bits_sdq_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T65) begin
      state <= T63;
    end else if(T61) begin
      state <= 4'h4;
    end else if(T38) begin
      state <= 4'h6;
    end else if(T37) begin
      state <= 4'h2;
    end else if(T35) begin
      state <= 4'h3;
    end else if(T33) begin
      state <= 4'h4;
    end else if(T32) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(reset) begin
      refill_cnt <= 2'h0;
    end else if(T25) begin
      refill_cnt <= T24;
    end
    if(T60) begin
      req_cmd <= io_req_bits_cmd;
    end else if(T85) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T60) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T125) begin
      meta_hazard <= 2'h1;
    end else if(T124) begin
      meta_hazard <= T123;
    end
    if(T60) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T60) begin
      req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
    end
    if(T60) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(reset) begin
      new_coh_state_state <= T154;
    end else if(T38) begin
      new_coh_state_state <= coh_on_hit_state;
    end else if(T172) begin
      new_coh_state_state <= coh_on_grant_state;
    end
  end
endmodule

module Arbiter_9(
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits = io_in_0_bits;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module Arbiter_10(
    output io_in_0_ready,
    input  io_in_0_valid,
    input [39:0] io_in_0_bits_addr,
    input [8:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [2:0] io_in_0_bits_typ,
    input [63:0] io_in_0_bits_data,
    input  io_in_0_bits_nack,
    input  io_in_0_bits_replay,
    input  io_in_0_bits_has_data,
    input [63:0] io_in_0_bits_data_word_bypass,
    input [63:0] io_in_0_bits_store_data,
    input  io_out_ready,
    output io_out_valid,
    output[39:0] io_out_bits_addr,
    output[8:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[2:0] io_out_bits_typ,
    output[63:0] io_out_bits_data,
    output io_out_bits_nack,
    output io_out_bits_replay,
    output io_out_bits_has_data,
    output[63:0] io_out_bits_data_word_bypass,
    output[63:0] io_out_bits_store_data,
    output io_chosen
);

  wire chosen;


  assign io_chosen = chosen;
  assign chosen = 1'h0;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_nack = io_in_0_bits_nack;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_valid = io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
endmodule

module IOMSHR(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_acquire_ready,
    output io_acquire_valid,
    output[25:0] io_acquire_bits_addr_block,
    output[1:0] io_acquire_bits_client_xact_id,
    output[1:0] io_acquire_bits_addr_beat,
    output io_acquire_bits_is_builtin_type,
    output[2:0] io_acquire_bits_a_type,
    output[16:0] io_acquire_bits_union,
    output[127:0] io_acquire_bits_data,
    input  io_grant_valid,
    input [1:0] io_grant_bits_addr_beat,
    input [1:0] io_grant_bits_client_xact_id,
    input [2:0] io_grant_bits_manager_xact_id,
    input  io_grant_bits_is_builtin_type,
    input [3:0] io_grant_bits_g_type,
    input [127:0] io_grant_bits_data,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[8:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    //output[63:0] io_resp_bits_data_word_bypass
    output[63:0] io_resp_bits_store_data
);

  reg [63:0] req_data;
  wire[63:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg [4:0] req_cmd;
  wire[4:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[63:0] T12;
  wire[63:0] T141;
  wire req_cmd_sc;
  wire[63:0] T13;
  wire[7:0] T14;
  wire[7:0] T15;
  wire[7:0] T16;
  wire[63:0] T17;
  wire[15:0] T18;
  wire[15:0] T19;
  wire[63:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  reg [63:0] grant_word;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[127:0] T25;
  wire[6:0] T26;
  wire T27;
  reg [39:0] req_addr;
  wire[39:0] T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  reg [1:0] state;
  wire[1:0] T142;
  wire[1:0] T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T143;
  wire T55;
  wire T56;
  wire T57;
  wire[2:0] T58;
  reg [2:0] req_typ;
  wire[2:0] T59;
  wire T60;
  wire[1:0] T61;
  wire[15:0] T62;
  wire T63;
  wire[47:0] T64;
  wire[47:0] T65;
  wire[47:0] T66;
  wire[47:0] T144;
  wire T67;
  wire T68;
  wire T69;
  wire[7:0] T70;
  wire T71;
  wire[55:0] T72;
  wire[55:0] T73;
  wire[55:0] T74;
  wire[55:0] T145;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  reg [8:0] req_tag;
  wire[8:0] T79;
  wire T80;
  wire[127:0] T81;
  wire[127:0] put_acquire_data;
  wire[127:0] beat_data;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[31:0] T86;
  wire T87;
  wire[1:0] T88;
  wire[63:0] T89;
  wire[31:0] T90;
  wire[15:0] T91;
  wire T92;
  wire[63:0] T93;
  wire[31:0] T94;
  wire[15:0] T95;
  wire[7:0] T96;
  wire T97;
  wire[127:0] get_acquire_data;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire[16:0] T107;
  wire[16:0] put_acquire_union;
  wire[16:0] T146;
  wire[23:0] T108;
  wire[22:0] beat_mask;
  wire[3:0] T109;
  wire beat_offset;
  wire[7:0] T110;
  wire[3:0] T111;
  wire[3:0] T112;
  wire[1:0] T113;
  wire[1:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire[1:0] T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire T129;
  wire[3:0] T130;
  wire T131;
  wire[16:0] get_acquire_union;
  wire[16:0] T147;
  wire[12:0] T132;
  wire[6:0] T133;
  wire[3:0] addr_byte;
  wire[2:0] T134;
  wire[2:0] put_acquire_a_type;
  wire[2:0] get_acquire_a_type;
  wire T135;
  wire put_acquire_is_builtin_type;
  wire get_acquire_is_builtin_type;
  wire[1:0] T136;
  wire[1:0] put_acquire_addr_beat;
  wire[1:0] addr_beat;
  wire[1:0] get_acquire_addr_beat;
  wire[1:0] T137;
  wire[1:0] put_acquire_client_xact_id;
  wire[1:0] get_acquire_client_xact_id;
  wire[25:0] T138;
  wire[25:0] put_acquire_addr_block;
  wire[25:0] addr_block;
  wire[25:0] get_acquire_addr_block;
  wire T139;
  wire T140;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    req_data = {2{$random}};
    req_cmd = {1{$random}};
    grant_word = {2{$random}};
    req_addr = {2{$random}};
    state = {1{$random}};
    req_typ = {1{$random}};
    req_tag = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_resp_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  assign io_resp_bits_store_data = req_data;
  assign T0 = T1 ? io_req_bits_data : req_data;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_has_data = T2;
  assign T2 = T7 | T3;
  assign T3 = T6 | T4;
  assign T4 = req_cmd == 5'h4;
  assign T5 = T1 ? io_req_bits_cmd : req_cmd;
  assign T6 = req_cmd[2'h3:2'h3];
  assign T7 = T9 | T8;
  assign T8 = req_cmd == 5'h7;
  assign T9 = T11 | T10;
  assign T10 = req_cmd == 5'h6;
  assign T11 = req_cmd == 5'h0;
  assign io_resp_bits_replay = io_resp_valid;
  assign io_resp_bits_nack = 1'h0;
  assign io_resp_bits_data = T12;
  assign T12 = T13 | T141;
  assign T141 = {63'h0, req_cmd_sc};
  assign req_cmd_sc = req_cmd == 5'h7;
  assign T13 = {T72, T14};
  assign T14 = req_cmd_sc ? 8'h0 : T15;
  assign T15 = T71 ? T70 : T16;
  assign T16 = T17[3'h7:1'h0];
  assign T17 = {T64, T18};
  assign T18 = T63 ? T62 : T19;
  assign T19 = T20[4'hf:1'h0];
  assign T20 = {T52, T21};
  assign T21 = T51 ? T50 : T22;
  assign T22 = grant_word[5'h1f:1'h0];
  assign T23 = T29 ? T24 : grant_word;
  assign T24 = T25[6'h3f:1'h0];
  assign T25 = io_grant_bits_data >> T26;
  assign T26 = {T27, 6'h0};
  assign T27 = req_addr[2'h3:2'h3];
  assign T28 = T1 ? io_req_bits_addr : req_addr;
  assign T29 = T39 & T30;
  assign T30 = T34 | T31;
  assign T31 = T33 | T32;
  assign T32 = req_cmd == 5'h4;
  assign T33 = req_cmd[2'h3:2'h3];
  assign T34 = T36 | T35;
  assign T35 = req_cmd == 5'h7;
  assign T36 = T38 | T37;
  assign T37 = req_cmd == 5'h6;
  assign T38 = req_cmd == 5'h0;
  assign T39 = T40 & io_grant_valid;
  assign T40 = state == 2'h2;
  assign T142 = reset ? 2'h0 : T41;
  assign T41 = T49 ? 2'h0 : T42;
  assign T42 = T47 ? 2'h0 : T43;
  assign T43 = T29 ? 2'h3 : T44;
  assign T44 = T46 ? 2'h2 : T45;
  assign T45 = T1 ? 2'h1 : state;
  assign T46 = io_acquire_ready & io_acquire_valid;
  assign T47 = T39 & T48;
  assign T48 = T30 ^ 1'h1;
  assign T49 = io_resp_ready & io_resp_valid;
  assign T50 = grant_word[6'h3f:6'h20];
  assign T51 = req_addr[2'h2:2'h2];
  assign T52 = T60 ? T54 : T53;
  assign T53 = grant_word[6'h3f:6'h20];
  assign T54 = 32'h0 - T143;
  assign T143 = {31'h0, T55};
  assign T55 = T57 & T56;
  assign T56 = T21[5'h1f:5'h1f];
  assign T57 = $signed(1'h0) <= $signed(T58);
  assign T58 = req_typ;
  assign T59 = T1 ? io_req_bits_typ : req_typ;
  assign T60 = T61 == 2'h2;
  assign T61 = req_typ[1'h1:1'h0];
  assign T62 = T20[5'h1f:5'h10];
  assign T63 = req_addr[1'h1:1'h1];
  assign T64 = T69 ? T66 : T65;
  assign T65 = T20[6'h3f:5'h10];
  assign T66 = 48'h0 - T144;
  assign T144 = {47'h0, T67};
  assign T67 = T57 & T68;
  assign T68 = T18[4'hf:4'hf];
  assign T69 = T61 == 2'h1;
  assign T70 = T17[4'hf:4'h8];
  assign T71 = req_addr[1'h0:1'h0];
  assign T72 = T77 ? T74 : T73;
  assign T73 = T17[6'h3f:4'h8];
  assign T74 = 56'h0 - T145;
  assign T145 = {55'h0, T75};
  assign T75 = T57 & T76;
  assign T76 = T14[3'h7:3'h7];
  assign T77 = T78 | req_cmd_sc;
  assign T78 = T61 == 2'h0;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_tag = req_tag;
  assign T79 = T1 ? io_req_bits_tag : req_tag;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_valid = T80;
  assign T80 = state == 2'h3;
  assign io_acquire_bits_data = T81;
  assign T81 = T98 ? get_acquire_data : put_acquire_data;
  assign put_acquire_data = beat_data;
  assign beat_data = {T82, T82};
  assign T82 = T97 ? T93 : T83;
  assign T83 = T92 ? T89 : T84;
  assign T84 = T87 ? T85 : req_data;
  assign T85 = {T86, T86};
  assign T86 = req_data[5'h1f:1'h0];
  assign T87 = T88 == 2'h2;
  assign T88 = req_typ[1'h1:1'h0];
  assign T89 = {T90, T90};
  assign T90 = {T91, T91};
  assign T91 = req_data[4'hf:1'h0];
  assign T92 = T88 == 2'h1;
  assign T93 = {T94, T94};
  assign T94 = {T95, T95};
  assign T95 = {T96, T96};
  assign T96 = req_data[3'h7:1'h0];
  assign T97 = T88 == 2'h0;
  assign get_acquire_data = 128'h0;
  assign T98 = T102 | T99;
  assign T99 = T101 | T100;
  assign T100 = req_cmd == 5'h4;
  assign T101 = req_cmd[2'h3:2'h3];
  assign T102 = T104 | T103;
  assign T103 = req_cmd == 5'h7;
  assign T104 = T106 | T105;
  assign T105 = req_cmd == 5'h6;
  assign T106 = req_cmd == 5'h0;
  assign io_acquire_bits_union = T107;
  assign T107 = T98 ? get_acquire_union : put_acquire_union;
  assign put_acquire_union = T146;
  assign T146 = T108[5'h10:1'h0];
  assign T108 = {beat_mask, 1'h0};
  assign beat_mask = T110 << T109;
  assign T109 = {beat_offset, 3'h0};
  assign beat_offset = req_addr[2'h3:2'h3];
  assign T110 = {T127, T111};
  assign T111 = T126 ? 4'h0 : T112;
  assign T112 = {T121, T113};
  assign T113 = T120 ? 2'h0 : T114;
  assign T114 = {T117, T115};
  assign T115 = T116 == 1'h0;
  assign T116 = req_addr[1'h0:1'h0];
  assign T117 = T119 | T118;
  assign T118 = 2'h1 <= T88;
  assign T119 = req_addr[1'h0:1'h0];
  assign T120 = req_addr[1'h1:1'h1];
  assign T121 = T124 | T122;
  assign T122 = T123 ? 2'h3 : 2'h0;
  assign T123 = 2'h2 <= T88;
  assign T124 = T125 ? T114 : 2'h0;
  assign T125 = req_addr[1'h1:1'h1];
  assign T126 = req_addr[2'h2:2'h2];
  assign T127 = T130 | T128;
  assign T128 = T129 ? 4'hf : 4'h0;
  assign T129 = 2'h3 <= T88;
  assign T130 = T131 ? T112 : 4'h0;
  assign T131 = req_addr[2'h2:2'h2];
  assign get_acquire_union = T147;
  assign T147 = {4'h0, T132};
  assign T132 = {T133, 6'h0};
  assign T133 = {addr_byte, req_typ};
  assign addr_byte = req_addr[2'h3:1'h0];
  assign io_acquire_bits_a_type = T134;
  assign T134 = T98 ? get_acquire_a_type : put_acquire_a_type;
  assign put_acquire_a_type = 3'h2;
  assign get_acquire_a_type = 3'h0;
  assign io_acquire_bits_is_builtin_type = T135;
  assign T135 = T98 ? get_acquire_is_builtin_type : put_acquire_is_builtin_type;
  assign put_acquire_is_builtin_type = 1'h1;
  assign get_acquire_is_builtin_type = 1'h1;
  assign io_acquire_bits_addr_beat = T136;
  assign T136 = T98 ? get_acquire_addr_beat : put_acquire_addr_beat;
  assign put_acquire_addr_beat = addr_beat;
  assign addr_beat = req_addr[3'h5:3'h4];
  assign get_acquire_addr_beat = addr_beat;
  assign io_acquire_bits_client_xact_id = T137;
  assign T137 = T98 ? get_acquire_client_xact_id : put_acquire_client_xact_id;
  assign put_acquire_client_xact_id = 2'h2;
  assign get_acquire_client_xact_id = 2'h2;
  assign io_acquire_bits_addr_block = T138;
  assign T138 = T98 ? get_acquire_addr_block : put_acquire_addr_block;
  assign put_acquire_addr_block = addr_block;
  assign addr_block = req_addr[5'h1f:3'h6];
  assign get_acquire_addr_block = addr_block;
  assign io_acquire_valid = T139;
  assign T139 = state == 2'h1;
  assign io_req_ready = T140;
  assign T140 = state == 2'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_data <= io_req_bits_data;
    end
    if(T1) begin
      req_cmd <= io_req_bits_cmd;
    end
    if(T29) begin
      grant_word <= T24;
    end
    if(T1) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T49) begin
      state <= 2'h0;
    end else if(T47) begin
      state <= 2'h0;
    end else if(T29) begin
      state <= 2'h3;
    end else if(T46) begin
      state <= 2'h2;
    end else if(T1) begin
      state <= 2'h1;
    end
    if(T1) begin
      req_typ <= io_req_bits_typ;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [39:0] io_req_bits_addr,
    input [8:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_kill,
    input  io_req_bits_phys,
    input [63:0] io_req_bits_data,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input  io_resp_ready,
    output io_resp_valid,
    output[39:0] io_resp_bits_addr,
    output[8:0] io_resp_bits_tag,
    output[4:0] io_resp_bits_cmd,
    output[2:0] io_resp_bits_typ,
    output[63:0] io_resp_bits_data,
    output io_resp_bits_nack,
    output io_resp_bits_replay,
    output io_resp_bits_has_data,
    output[63:0] io_resp_bits_data_word_bypass,
    output[63:0] io_resp_bits_store_data,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr_block,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[1:0] io_mem_req_bits_addr_beat,
    output io_mem_req_bits_is_builtin_type,
    output[2:0] io_mem_req_bits_a_type,
    output[16:0] io_mem_req_bits_union,
    output[127:0] io_mem_req_bits_data,
    output io_refill_way_en,
    output[11:0] io_refill_addr,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output[39:0] io_replay_bits_addr,
    output[8:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_kill,
    output io_replay_bits_phys,
    output[63:0] io_replay_bits_data,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[1:0] io_wb_req_bits_addr_beat,
    output[25:0] io_wb_req_bits_addr_block,
    output[1:0] io_wb_req_bits_client_xact_id,
    output io_wb_req_bits_voluntary,
    output[2:0] io_wb_req_bits_r_type,
    output[127:0] io_wb_req_bits_data,
    output io_wb_req_bits_way_en,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire cacheable;
  wire T4;
  wire T5;
  wire[4:0] T111;
  wire[4:0] T112;
  wire[4:0] T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire[4:0] T116;
  wire[4:0] T117;
  wire[4:0] T118;
  wire[4:0] T119;
  wire[4:0] T120;
  wire[4:0] T121;
  wire[4:0] T122;
  wire[4:0] T123;
  wire[4:0] T124;
  wire[4:0] T125;
  wire[4:0] T126;
  wire T127;
  wire[16:0] T6;
  wire[16:0] T7;
  reg [16:0] sdq_val;
  wire[16:0] T128;
  wire[31:0] T129;
  wire[31:0] T8;
  wire[31:0] T130;
  wire[31:0] T9;
  wire[31:0] T131;
  wire[16:0] T10;
  wire[16:0] T11;
  wire[16:0] T132;
  wire sdq_enq;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[16:0] T21;
  wire[16:0] T22;
  wire[16:0] T23;
  wire[16:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire[16:0] T28;
  wire[16:0] T29;
  wire[16:0] T30;
  wire[16:0] T31;
  wire[16:0] T32;
  wire[16:0] T33;
  wire[16:0] T34;
  wire[16:0] T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire[31:0] T57;
  wire[31:0] T58;
  wire[31:0] T59;
  wire[31:0] T133;
  wire[16:0] T60;
  wire[16:0] T134;
  wire free_sdq;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire[31:0] T69;
  wire[31:0] T135;
  wire T70;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T71;
  wire tag_match;
  wire[27:0] T72;
  wire[27:0] T151;
  wire[19:0] T73;
  wire[19:0] T74;
  wire[19:0] tagList_1;
  wire idxMatch_1;
  wire[19:0] T75;
  wire[19:0] tagList_0;
  wire idxMatch_0;
  wire T76;
  wire sdq_rdy;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire idx_match;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[63:0] T96;
  reg [63:0] sdq [16:0];
  wire[63:0] T97;
  wire T98;
  wire T99;
  wire[4:0] T100;
  reg [4:0] R101;
  wire[4:0] T102;
  wire[11:0] T103;
  wire[11:0] refillMux_0_addr;
  wire[11:0] refillMux_1_addr;
  wire T104;
  wire T152;
  wire T105;
  wire refillMux_0_way_en;
  wire refillMux_1_way_en;
  wire T106;
  wire T107;
  wire T108;
  wire pri_rdy;
  wire T109;
  wire sec_rdy;
  wire T110;
  wire meta_read_arb_io_in_1_ready;
  wire meta_read_arb_io_in_0_ready;
  wire meta_read_arb_io_out_valid;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire meta_write_arb_io_in_1_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_write_arb_io_out_valid;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire meta_write_arb_io_out_bits_way_en;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire mem_req_arb_io_in_2_ready;
  wire mem_req_arb_io_in_1_ready;
  wire mem_req_arb_io_in_0_ready;
  wire mem_req_arb_io_out_valid;
  wire[25:0] mem_req_arb_io_out_bits_addr_block;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[1:0] mem_req_arb_io_out_bits_addr_beat;
  wire mem_req_arb_io_out_bits_is_builtin_type;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[16:0] mem_req_arb_io_out_bits_union;
  wire[127:0] mem_req_arb_io_out_bits_data;
  wire wb_req_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire wb_req_arb_io_out_valid;
  wire[1:0] wb_req_arb_io_out_bits_addr_beat;
  wire[25:0] wb_req_arb_io_out_bits_addr_block;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire wb_req_arb_io_out_bits_voluntary;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire[127:0] wb_req_arb_io_out_bits_data;
  wire wb_req_arb_io_out_bits_way_en;
  wire replay_arb_io_in_1_ready;
  wire replay_arb_io_in_0_ready;
  wire replay_arb_io_out_valid;
  wire[39:0] replay_arb_io_out_bits_addr;
  wire[8:0] replay_arb_io_out_bits_tag;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_bits_phys;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire alloc_arb_io_in_1_ready;
  wire alloc_arb_io_in_0_ready;
  wire mmio_alloc_arb_io_in_0_ready;
  wire resp_arb_io_in_0_ready;
  wire resp_arb_io_out_valid;
  wire[39:0] resp_arb_io_out_bits_addr;
  wire[8:0] resp_arb_io_out_bits_tag;
  wire[4:0] resp_arb_io_out_bits_cmd;
  wire[2:0] resp_arb_io_out_bits_typ;
  wire[63:0] resp_arb_io_out_bits_data;
  wire resp_arb_io_out_bits_nack;
  wire resp_arb_io_out_bits_replay;
  wire resp_arb_io_out_bits_has_data;
  wire[63:0] resp_arb_io_out_bits_data_word_bypass;
  wire[63:0] resp_arb_io_out_bits_store_data;
  wire IOMSHR_io_req_ready;
  wire IOMSHR_io_acquire_valid;
  wire[25:0] IOMSHR_io_acquire_bits_addr_block;
  wire[1:0] IOMSHR_io_acquire_bits_client_xact_id;
  wire[1:0] IOMSHR_io_acquire_bits_addr_beat;
  wire IOMSHR_io_acquire_bits_is_builtin_type;
  wire[2:0] IOMSHR_io_acquire_bits_a_type;
  wire[16:0] IOMSHR_io_acquire_bits_union;
  wire[127:0] IOMSHR_io_acquire_bits_data;
  wire IOMSHR_io_resp_valid;
  wire[39:0] IOMSHR_io_resp_bits_addr;
  wire[8:0] IOMSHR_io_resp_bits_tag;
  wire[4:0] IOMSHR_io_resp_bits_cmd;
  wire[2:0] IOMSHR_io_resp_bits_typ;
  wire[63:0] IOMSHR_io_resp_bits_data;
  wire IOMSHR_io_resp_bits_nack;
  wire IOMSHR_io_resp_bits_replay;
  wire IOMSHR_io_resp_bits_has_data;
  wire[63:0] IOMSHR_io_resp_bits_store_data;
  wire MSHR_io_req_pri_rdy;
  wire MSHR_io_req_sec_rdy;
  wire MSHR_io_idx_match;
  wire[19:0] MSHR_io_tag;
  wire MSHR_io_mem_req_valid;
  wire[25:0] MSHR_io_mem_req_bits_addr_block;
  wire[1:0] MSHR_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_io_mem_req_bits_addr_beat;
  wire MSHR_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_io_mem_req_bits_a_type;
  wire[16:0] MSHR_io_mem_req_bits_union;
  wire[127:0] MSHR_io_mem_req_bits_data;
  wire MSHR_io_refill_way_en;
  wire[11:0] MSHR_io_refill_addr;
  wire MSHR_io_meta_read_valid;
  wire[5:0] MSHR_io_meta_read_bits_idx;
  wire[19:0] MSHR_io_meta_read_bits_tag;
  wire MSHR_io_meta_write_valid;
  wire[5:0] MSHR_io_meta_write_bits_idx;
  wire MSHR_io_meta_write_bits_way_en;
  wire[19:0] MSHR_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_io_meta_write_bits_data_coh_state;
  wire MSHR_io_replay_valid;
  wire[39:0] MSHR_io_replay_bits_addr;
  wire[8:0] MSHR_io_replay_bits_tag;
  wire[4:0] MSHR_io_replay_bits_cmd;
  wire[2:0] MSHR_io_replay_bits_typ;
  wire MSHR_io_replay_bits_kill;
  wire MSHR_io_replay_bits_phys;
  wire[4:0] MSHR_io_replay_bits_sdq_id;
  wire MSHR_io_wb_req_valid;
  wire[1:0] MSHR_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_io_wb_req_bits_addr_block;
  wire[1:0] MSHR_io_wb_req_bits_client_xact_id;
  wire MSHR_io_wb_req_bits_voluntary;
  wire[2:0] MSHR_io_wb_req_bits_r_type;
  wire[127:0] MSHR_io_wb_req_bits_data;
  wire MSHR_io_wb_req_bits_way_en;
  wire MSHR_io_probe_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_1_io_idx_match;
  wire[19:0] MSHR_1_io_tag;
  wire MSHR_1_io_mem_req_valid;
  wire[25:0] MSHR_1_io_mem_req_bits_addr_block;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[1:0] MSHR_1_io_mem_req_bits_addr_beat;
  wire MSHR_1_io_mem_req_bits_is_builtin_type;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[16:0] MSHR_1_io_mem_req_bits_union;
  wire[127:0] MSHR_1_io_mem_req_bits_data;
  wire MSHR_1_io_refill_way_en;
  wire[11:0] MSHR_1_io_refill_addr;
  wire MSHR_1_io_meta_read_valid;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire MSHR_1_io_meta_write_valid;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire MSHR_1_io_meta_write_bits_way_en;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire MSHR_1_io_replay_valid;
  wire[39:0] MSHR_1_io_replay_bits_addr;
  wire[8:0] MSHR_1_io_replay_bits_tag;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_bits_phys;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire MSHR_1_io_wb_req_valid;
  wire[1:0] MSHR_1_io_wb_req_bits_addr_beat;
  wire[25:0] MSHR_1_io_wb_req_bits_addr_block;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire MSHR_1_io_wb_req_bits_voluntary;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire[127:0] MSHR_1_io_wb_req_bits_data;
  wire MSHR_1_io_wb_req_bits_way_en;
  wire MSHR_1_io_probe_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R101 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_mem_grant_valid & T1;
  assign T1 = io_mem_grant_bits_client_xact_id == 2'h2;
  assign T2 = io_req_valid & T3;
  assign T3 = cacheable ^ 1'h1;
  assign cacheable = io_req_bits_addr < 40'h40000000;
  assign T4 = io_mem_grant_valid & T5;
  assign T5 = io_mem_grant_bits_client_xact_id == 2'h1;
  assign T111 = T150 ? 1'h0 : T112;
  assign T112 = T149 ? 1'h1 : T113;
  assign T113 = T148 ? 2'h2 : T114;
  assign T114 = T147 ? 2'h3 : T115;
  assign T115 = T146 ? 3'h4 : T116;
  assign T116 = T145 ? 3'h5 : T117;
  assign T117 = T144 ? 3'h6 : T118;
  assign T118 = T143 ? 3'h7 : T119;
  assign T119 = T142 ? 4'h8 : T120;
  assign T120 = T141 ? 4'h9 : T121;
  assign T121 = T140 ? 4'ha : T122;
  assign T122 = T139 ? 4'hb : T123;
  assign T123 = T138 ? 4'hc : T124;
  assign T124 = T137 ? 4'hd : T125;
  assign T125 = T136 ? 4'he : T126;
  assign T126 = T127 ? 4'hf : 5'h10;
  assign T127 = T6[4'hf:4'hf];
  assign T6 = ~ T7;
  assign T7 = sdq_val[5'h10:1'h0];
  assign T128 = T129[5'h10:1'h0];
  assign T129 = reset ? 32'h0 : T8;
  assign T8 = T70 ? T9 : T130;
  assign T130 = {15'h0, sdq_val};
  assign T9 = T57 | T131;
  assign T131 = {15'h0, T10};
  assign T10 = T21 & T11;
  assign T11 = 17'h0 - T132;
  assign T132 = {16'h0, sdq_enq};
  assign sdq_enq = T19 & T12;
  assign T12 = T16 | T13;
  assign T13 = T15 | T14;
  assign T14 = io_req_bits_cmd == 5'h4;
  assign T15 = io_req_bits_cmd[2'h3:2'h3];
  assign T16 = T18 | T17;
  assign T17 = io_req_bits_cmd == 5'h7;
  assign T18 = io_req_bits_cmd == 5'h1;
  assign T19 = T20 & cacheable;
  assign T20 = io_req_valid & io_req_ready;
  assign T21 = T56 ? 17'h1 : T22;
  assign T22 = T55 ? 17'h2 : T23;
  assign T23 = T54 ? 17'h4 : T24;
  assign T24 = T53 ? 17'h8 : T25;
  assign T25 = T52 ? 17'h10 : T26;
  assign T26 = T51 ? 17'h20 : T27;
  assign T27 = T50 ? 17'h40 : T28;
  assign T28 = T49 ? 17'h80 : T29;
  assign T29 = T48 ? 17'h100 : T30;
  assign T30 = T47 ? 17'h200 : T31;
  assign T31 = T46 ? 17'h400 : T32;
  assign T32 = T45 ? 17'h800 : T33;
  assign T33 = T44 ? 17'h1000 : T34;
  assign T34 = T43 ? 17'h2000 : T35;
  assign T35 = T42 ? 17'h4000 : T36;
  assign T36 = T41 ? 17'h8000 : T37;
  assign T37 = T38 ? 17'h10000 : 17'h0;
  assign T38 = T39[5'h10:5'h10];
  assign T39 = ~ T40;
  assign T40 = sdq_val[5'h10:1'h0];
  assign T41 = T39[4'hf:4'hf];
  assign T42 = T39[4'he:4'he];
  assign T43 = T39[4'hd:4'hd];
  assign T44 = T39[4'hc:4'hc];
  assign T45 = T39[4'hb:4'hb];
  assign T46 = T39[4'ha:4'ha];
  assign T47 = T39[4'h9:4'h9];
  assign T48 = T39[4'h8:4'h8];
  assign T49 = T39[3'h7:3'h7];
  assign T50 = T39[3'h6:3'h6];
  assign T51 = T39[3'h5:3'h5];
  assign T52 = T39[3'h4:3'h4];
  assign T53 = T39[2'h3:2'h3];
  assign T54 = T39[2'h2:2'h2];
  assign T55 = T39[1'h1:1'h1];
  assign T56 = T39[1'h0:1'h0];
  assign T57 = T135 & T58;
  assign T58 = ~ T59;
  assign T59 = T69 & T133;
  assign T133 = {15'h0, T60};
  assign T60 = 17'h0 - T134;
  assign T134 = {16'h0, free_sdq};
  assign free_sdq = T68 & T61;
  assign T61 = T65 | T62;
  assign T62 = T64 | T63;
  assign T63 = io_replay_bits_cmd == 5'h4;
  assign T64 = io_replay_bits_cmd[2'h3:2'h3];
  assign T65 = T67 | T66;
  assign T66 = io_replay_bits_cmd == 5'h7;
  assign T67 = io_replay_bits_cmd == 5'h1;
  assign T68 = io_replay_ready & io_replay_valid;
  assign T69 = 1'h1 << replay_arb_io_out_bits_sdq_id;
  assign T135 = {15'h0, sdq_val};
  assign T70 = io_replay_valid | sdq_enq;
  assign T136 = T6[4'he:4'he];
  assign T137 = T6[4'hd:4'hd];
  assign T138 = T6[4'hc:4'hc];
  assign T139 = T6[4'hb:4'hb];
  assign T140 = T6[4'ha:4'ha];
  assign T141 = T6[4'h9:4'h9];
  assign T142 = T6[4'h8:4'h8];
  assign T143 = T6[3'h7:3'h7];
  assign T144 = T6[3'h6:3'h6];
  assign T145 = T6[3'h5:3'h5];
  assign T146 = T6[3'h4:3'h4];
  assign T147 = T6[2'h3:2'h3];
  assign T148 = T6[2'h2:2'h2];
  assign T149 = T6[1'h1:1'h1];
  assign T150 = T6[1'h0:1'h0];
  assign T71 = T76 & tag_match;
  assign tag_match = T151 == T72;
  assign T72 = io_req_bits_addr >> 4'hc;
  assign T151 = {8'h0, T73};
  assign T73 = T75 | T74;
  assign T74 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T75 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_io_tag;
  assign idxMatch_0 = MSHR_io_idx_match;
  assign T76 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T77 ^ 1'h1;
  assign T77 = sdq_val == 17'h1ffff;
  assign T78 = io_mem_grant_valid & T79;
  assign T79 = io_mem_grant_bits_client_xact_id == 2'h0;
  assign T80 = T81 & tag_match;
  assign T81 = io_req_valid & sdq_rdy;
  assign T82 = T84 & T83;
  assign T83 = idx_match ^ 1'h1;
  assign idx_match = MSHR_io_idx_match | MSHR_1_io_idx_match;
  assign T84 = T85 & cacheable;
  assign T85 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T86;
  assign T86 = T91 ? 1'h0 : T87;
  assign T87 = T90 ? 1'h0 : T88;
  assign T88 = T89 == 1'h0;
  assign T89 = MSHR_io_req_pri_rdy ^ 1'h1;
  assign T90 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign T91 = IOMSHR_io_req_ready ^ 1'h1;
  assign io_probe_rdy = T92;
  assign T92 = T95 ? 1'h0 : T93;
  assign T93 = T94 == 1'h0;
  assign T94 = MSHR_io_probe_rdy ^ 1'h1;
  assign T95 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_replay_bits_data = T96;
  assign T96 = sdq[R101];
  assign T98 = sdq_enq & T99;
  assign T99 = T100 < 5'h11;
  assign T100 = T111[3'h4:1'h0];
  assign T102 = free_sdq ? replay_arb_io_out_bits_sdq_id : R101;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_refill_addr = T103;
  assign T103 = T104 ? refillMux_1_addr : refillMux_0_addr;
  assign refillMux_0_addr = MSHR_io_refill_addr;
  assign refillMux_1_addr = MSHR_1_io_refill_addr;
  assign T104 = T152;
  assign T152 = io_mem_grant_bits_client_xact_id[1'h0:1'h0];
  assign io_refill_way_en = T105;
  assign T105 = T104 ? refillMux_1_way_en : refillMux_0_way_en;
  assign refillMux_0_way_en = MSHR_io_refill_way_en;
  assign refillMux_1_way_en = MSHR_1_io_refill_way_en;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_nack = resp_arb_io_out_bits_nack;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_req_ready = T106;
  assign T106 = T110 ? IOMSHR_io_req_ready : T107;
  assign T107 = T108 & sdq_rdy;
  assign T108 = idx_match ? T109 : pri_rdy;
  assign pri_rdy = MSHR_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T109 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  assign T110 = cacheable ^ 1'h1;
  Arbiter_6 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  LockingArbiter_1 mem_req_arb(.clk(clk), .reset(reset),
       .io_in_2_ready( mem_req_arb_io_in_2_ready ),
       .io_in_2_valid( IOMSHR_io_acquire_valid ),
       .io_in_2_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_in_2_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_in_2_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_in_2_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_in_2_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_in_2_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_in_2_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_in_1_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_in_1_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_in_1_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_in_1_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_mem_req_valid ),
       .io_in_0_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_in_0_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_in_0_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_in_0_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_in_0_bits_union( MSHR_io_mem_req_bits_union ),
       .io_in_0_bits_data( MSHR_io_mem_req_bits_data ),
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr_block( mem_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_addr_beat( mem_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_is_builtin_type( mem_req_arb_io_out_bits_is_builtin_type ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_union( mem_req_arb_io_out_bits_union ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_1_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_in_0_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_in_0_bits_data( MSHR_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_addr_beat( wb_req_arb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wb_req_arb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( wb_req_arb_io_out_bits_voluntary ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type ),
       .io_out_bits_data( wb_req_arb_io_out_bits_data ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en )
       //.io_chosen(  )
  );
  Arbiter_7 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_replay_valid ),
       .io_in_0_bits_addr( MSHR_io_replay_bits_addr ),
       .io_in_0_bits_tag( MSHR_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_in_0_bits_typ( MSHR_io_replay_bits_typ ),
       .io_in_0_bits_kill( MSHR_io_replay_bits_kill ),
       .io_in_0_bits_phys( MSHR_io_replay_bits_phys ),
       .io_in_0_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_8 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T82 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  MSHR_0 MSHR(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_io_req_pri_rdy ),
       .io_req_sec_val( T80 ),
       .io_req_sec_rdy( MSHR_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T111 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_io_idx_match ),
       .io_tag( MSHR_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_io_refill_way_en ),
       .io_refill_addr( MSHR_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_io_replay_valid ),
       .io_replay_bits_addr( MSHR_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T78 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( MSHR_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( MSHR_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( MSHR_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_io_probe_rdy )
  );
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T71 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_sdq_id( T111 ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( MSHR_1_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( MSHR_1_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( MSHR_1_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( MSHR_1_io_mem_req_bits_union ),
       .io_mem_req_bits_data( MSHR_1_io_mem_req_bits_data ),
       .io_refill_way_en( MSHR_1_io_refill_way_en ),
       .io_refill_addr( MSHR_1_io_refill_addr ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( T4 ),
       .io_mem_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_mem_grant_bits_data ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( MSHR_1_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( MSHR_1_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( MSHR_1_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( MSHR_1_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  Arbiter_9 mmio_alloc_arb(
       .io_in_0_ready( mmio_alloc_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_req_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T2 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign mmio_alloc_arb.io_in_0_bits = {1{$random}};
// synthesis translate_on
`endif
  Arbiter_10 resp_arb(
       .io_in_0_ready( resp_arb_io_in_0_ready ),
       .io_in_0_valid( IOMSHR_io_resp_valid ),
       .io_in_0_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_in_0_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_in_0_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_in_0_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_in_0_bits_data( IOMSHR_io_resp_bits_data ),
       .io_in_0_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_in_0_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_in_0_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_in_0_bits_data_word_bypass(  )
       .io_in_0_bits_store_data( IOMSHR_io_resp_bits_store_data ),
       .io_out_ready( io_resp_ready ),
       .io_out_valid( resp_arb_io_out_valid ),
       .io_out_bits_addr( resp_arb_io_out_bits_addr ),
       .io_out_bits_tag( resp_arb_io_out_bits_tag ),
       .io_out_bits_cmd( resp_arb_io_out_bits_cmd ),
       .io_out_bits_typ( resp_arb_io_out_bits_typ ),
       .io_out_bits_data( resp_arb_io_out_bits_data ),
       .io_out_bits_nack( resp_arb_io_out_bits_nack ),
       .io_out_bits_replay( resp_arb_io_out_bits_replay ),
       .io_out_bits_has_data( resp_arb_io_out_bits_has_data ),
       .io_out_bits_data_word_bypass( resp_arb_io_out_bits_data_word_bypass ),
       .io_out_bits_store_data( resp_arb_io_out_bits_store_data )
       //.io_chosen(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign resp_arb.io_in_0_bits_data_word_bypass = {2{$random}};
// synthesis translate_on
`endif
  IOMSHR IOMSHR(.clk(clk), .reset(reset),
       .io_req_ready( IOMSHR_io_req_ready ),
       .io_req_valid( mmio_alloc_arb_io_in_0_ready ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_data( io_req_bits_data ),
       .io_acquire_ready( mem_req_arb_io_in_2_ready ),
       .io_acquire_valid( IOMSHR_io_acquire_valid ),
       .io_acquire_bits_addr_block( IOMSHR_io_acquire_bits_addr_block ),
       .io_acquire_bits_client_xact_id( IOMSHR_io_acquire_bits_client_xact_id ),
       .io_acquire_bits_addr_beat( IOMSHR_io_acquire_bits_addr_beat ),
       .io_acquire_bits_is_builtin_type( IOMSHR_io_acquire_bits_is_builtin_type ),
       .io_acquire_bits_a_type( IOMSHR_io_acquire_bits_a_type ),
       .io_acquire_bits_union( IOMSHR_io_acquire_bits_union ),
       .io_acquire_bits_data( IOMSHR_io_acquire_bits_data ),
       .io_grant_valid( T0 ),
       .io_grant_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_grant_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_grant_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_grant_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_grant_bits_g_type( io_mem_grant_bits_g_type ),
       .io_grant_bits_data( io_mem_grant_bits_data ),
       .io_resp_ready( resp_arb_io_in_0_ready ),
       .io_resp_valid( IOMSHR_io_resp_valid ),
       .io_resp_bits_addr( IOMSHR_io_resp_bits_addr ),
       .io_resp_bits_tag( IOMSHR_io_resp_bits_tag ),
       .io_resp_bits_cmd( IOMSHR_io_resp_bits_cmd ),
       .io_resp_bits_typ( IOMSHR_io_resp_bits_typ ),
       .io_resp_bits_data( IOMSHR_io_resp_bits_data ),
       .io_resp_bits_nack( IOMSHR_io_resp_bits_nack ),
       .io_resp_bits_replay( IOMSHR_io_resp_bits_replay ),
       .io_resp_bits_has_data( IOMSHR_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( IOMSHR_io_resp_bits_store_data )
  );

  always @(posedge clk) begin
    sdq_val <= T128;
    if (T98)
      sdq[T111] <= io_req_bits_data;
    if(free_sdq) begin
      R101 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input  io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[21:0] tags;
  wire[21:0] T1;
  wire[21:0] T2;
  wire[21:0] T3;
  wire[21:0] T4;
  wire[21:0] T5;
  wire[21:0] T24;
  wire T6;
  wire T7;
  wire T8;
  wire rst;
  reg [6:0] rst_cnt;
  wire[6:0] T25;
  wire[6:0] T9;
  wire[6:0] T10;
  wire[21:0] T11;
  wire[21:0] wdata;
  wire[21:0] T12;
  wire[1:0] T13;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T14;
  wire[19:0] T15;
  wire[19:0] rstVal_tag;
  wire T16;
  wire[5:0] T26;
  wire[6:0] waddr;
  wire[6:0] T27;
  reg [5:0] R17;
  wire[5:0] T18;
  wire[19:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R17 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = tags[1'h1:1'h0];
  assign tags = T1;
  assign T1 = T2[5'h15:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T26),
    .W0E(T16),
    .W0I(T11),
    .W0M(T4),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(T2)
  );
  assign T4 = T5;
  assign T5 = 22'h0 - T24;
  assign T24 = {21'h0, T6};
  assign T6 = T7;
  assign T7 = rst ? 1'h1 : T8;
  assign T8 = io_write_bits_way_en;
  assign rst = rst_cnt < 7'h40;
  assign T25 = reset ? 7'h0 : T9;
  assign T9 = rst ? T10 : rst_cnt;
  assign T10 = rst_cnt + 7'h1;
  assign T11 = wdata;
  assign wdata = T12;
  assign T12 = {T15, T13};
  assign T13 = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T14;
  assign T14 = 2'h0;
  assign T15 = rst ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T16 = rst | io_write_valid;
  assign T26 = waddr[3'h5:1'h0];
  assign waddr = rst ? rst_cnt : T27;
  assign T27 = {1'h0, io_write_bits_idx};
  assign T18 = io_read_valid ? io_read_bits_idx : R17;
  assign io_resp_0_tag = T19;
  assign T19 = tags[5'h15:2'h2];
  assign io_write_ready = T20;
  assign T20 = rst ^ 1'h1;
  assign io_read_ready = T21;
  assign T21 = T23 & T22;
  assign T22 = io_write_valid ^ 1'h1;
  assign T23 = rst ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(rst) begin
      rst_cnt <= T10;
    end
    if(io_read_valid) begin
      R17 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_0(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] chosen;
  wire[2:0] choose;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire[5:0] T5;
  wire T6;
  wire[2:0] T7;
  wire[5:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 3'h0 : T0;
  assign T0 = io_in_1_valid ? 3'h1 : T1;
  assign T1 = io_in_2_valid ? 3'h2 : T2;
  assign T2 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T3;
  assign T3 = T11 ? io_in_4_bits_idx : T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = chosen;
  assign T8 = T9 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign T11 = T7[2'h2:2'h2];
  assign io_out_valid = T12;
  assign T12 = T19 ? io_in_4_valid : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? io_in_1_valid : io_in_0_valid;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T17 ? io_in_3_valid : io_in_2_valid;
  assign T17 = T7[1'h0:1'h0];
  assign T18 = T7[1'h1:1'h1];
  assign T19 = T7[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = T28 | io_in_2_valid;
  assign T28 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T32 | io_in_3_valid;
  assign T32 = T33 | io_in_2_valid;
  assign T33 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input  io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire[127:0] T1;
  wire[63:0] T2;
  wire[127:0] T3;
  wire T19;
  wire[7:0] raddr;
  wire[127:0] T5;
  wire[127:0] T6;
  wire[127:0] T7;
  wire[63:0] T8;
  wire[63:0] T21;
  wire T9;
  wire[63:0] T10;
  wire[63:0] T22;
  wire T11;
  wire[127:0] T12;
  wire[127:0] T13;
  wire[63:0] T14;
  wire[63:0] T15;
  wire T16;
  wire[7:0] waddr;
  reg [7:0] R17;
  wire[7:0] T18;
  wire[63:0] T20;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_resp_0 = T0;
  assign T0 = T1;
  assign T1 = {T20, T2};
  assign T2 = T3[6'h3f:1'h0];
  assign T19 = io_read_bits_way_en & io_read_valid;
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T4 T4 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T16),
    .W0I(T12),
    .W0M(T6),
    .R1A(raddr),
    .R1E(T19),
    .R1O(T3)
  );
  assign T6 = T7;
  assign T7 = {T10, T8};
  assign T8 = 64'h0 - T21;
  assign T21 = {63'h0, T9};
  assign T9 = io_write_bits_wmask[1'h0:1'h0];
  assign T10 = 64'h0 - T22;
  assign T22 = {63'h0, T11};
  assign T11 = io_write_bits_wmask[1'h1:1'h1];
  assign T12 = T13;
  assign T13 = {T15, T14};
  assign T14 = io_write_bits_data[6'h3f:1'h0];
  assign T15 = io_write_bits_data[7'h7f:7'h40];
  assign T16 = io_write_bits_way_en & io_write_valid;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T18 = T19 ? raddr : R17;
  assign T20 = T3[7'h7f:7'h40];
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T19) begin
      R17 <= raddr;
    end
  end
endmodule

module Arbiter_2(
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] chosen;
  wire[1:0] choose;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[11:0] T2;
  wire[11:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[11:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid ? 2'h0 : T0;
  assign T0 = io_in_1_valid ? 2'h1 : T1;
  assign T1 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = chosen;
  assign T6 = T7 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T7 = T5[1'h0:1'h0];
  assign T8 = T5[1'h1:1'h1];
  assign io_out_bits_way_en = T9;
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T11 = T5[1'h0:1'h0];
  assign T12 = T13 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T13 = T5[1'h0:1'h0];
  assign T14 = T5[1'h1:1'h1];
  assign io_out_valid = T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T5[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T5[1'h0:1'h0];
  assign T20 = T5[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T25 ^ 1'h1;
  assign T25 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T26;
  assign T26 = T27 & io_out_ready;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T29 | io_in_2_valid;
  assign T29 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire[127:0] T0;
  wire T1;
  wire[1:0] T2;
  wire[11:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T0;
  assign T0 = T1 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T1 = chosen;
  assign io_out_bits_wmask = T2;
  assign T2 = T1 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T3;
  assign T3 = T1 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T4;
  assign T4 = T1 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T5;
  assign T5 = T1 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [4:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] wmask;
  wire[63:0] T3;
  wire[31:0] T4;
  wire[15:0] T5;
  wire[7:0] T6;
  wire[7:0] T119;
  wire T7;
  wire[7:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire T28;
  wire[3:0] T29;
  wire T30;
  wire[7:0] T31;
  wire[7:0] T120;
  wire T32;
  wire[15:0] T33;
  wire[7:0] T34;
  wire[7:0] T121;
  wire T35;
  wire[7:0] T36;
  wire[7:0] T122;
  wire T37;
  wire[31:0] T38;
  wire[15:0] T39;
  wire[7:0] T40;
  wire[7:0] T123;
  wire T41;
  wire[7:0] T42;
  wire[7:0] T124;
  wire T43;
  wire[15:0] T44;
  wire[7:0] T45;
  wire[7:0] T125;
  wire T46;
  wire[7:0] T47;
  wire[7:0] T126;
  wire T48;
  wire[63:0] T49;
  wire[63:0] out;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] T55;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[31:0] T58;
  wire T59;
  wire[63:0] T60;
  wire[31:0] T61;
  wire[15:0] T62;
  wire T63;
  wire[63:0] T64;
  wire[31:0] T65;
  wire[15:0] T66;
  wire[7:0] T67;
  wire T68;
  wire T69;
  wire max;
  wire T70;
  wire T71;
  wire min;
  wire T72;
  wire T73;
  wire less;
  wire T74;
  wire cmp_rhs;
  wire T75;
  wire[63:0] rhs;
  wire[63:0] T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire word;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire cmp_lhs;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire sgned;
  wire T94;
  wire T95;
  wire lt;
  wire T96;
  wire T97;
  wire lt_lo;
  wire[31:0] T98;
  wire[31:0] T99;
  wire eq_hi;
  wire[31:0] T100;
  wire[31:0] T101;
  wire lt_hi;
  wire[31:0] T102;
  wire[31:0] T103;
  wire T104;
  wire T105;
  wire T106;
  wire[63:0] T107;
  wire T108;
  wire[63:0] T109;
  wire T110;
  wire[63:0] T111;
  wire T112;
  wire[63:0] adder_out;
  wire[63:0] T113;
  wire[63:0] mask;
  wire[63:0] T127;
  wire[31:0] T114;
  wire T115;
  wire[63:0] T116;
  wire[63:0] T117;
  wire T118;


  assign io_out = T0;
  assign T0 = T49 | T1;
  assign T1 = T2 & io_lhs;
  assign T2 = ~ wmask;
  assign wmask = T3;
  assign T3 = {T38, T4};
  assign T4 = {T33, T5};
  assign T5 = {T31, T6};
  assign T6 = 8'h0 - T119;
  assign T119 = {7'h0, T7};
  assign T7 = T8[1'h0:1'h0];
  assign T8 = {T26, T9};
  assign T9 = T25 ? 4'h0 : T10;
  assign T10 = {T20, T11};
  assign T11 = T19 ? 2'h0 : T12;
  assign T12 = {T15, T13};
  assign T13 = T14 == 1'h0;
  assign T14 = io_addr[1'h0:1'h0];
  assign T15 = T18 | T16;
  assign T16 = 2'h1 <= T17;
  assign T17 = io_typ[1'h1:1'h0];
  assign T18 = io_addr[1'h0:1'h0];
  assign T19 = io_addr[1'h1:1'h1];
  assign T20 = T23 | T21;
  assign T21 = T22 ? 2'h3 : 2'h0;
  assign T22 = 2'h2 <= T17;
  assign T23 = T24 ? T12 : 2'h0;
  assign T24 = io_addr[1'h1:1'h1];
  assign T25 = io_addr[2'h2:2'h2];
  assign T26 = T29 | T27;
  assign T27 = T28 ? 4'hf : 4'h0;
  assign T28 = 2'h3 <= T17;
  assign T29 = T30 ? T10 : 4'h0;
  assign T30 = io_addr[2'h2:2'h2];
  assign T31 = 8'h0 - T120;
  assign T120 = {7'h0, T32};
  assign T32 = T8[1'h1:1'h1];
  assign T33 = {T36, T34};
  assign T34 = 8'h0 - T121;
  assign T121 = {7'h0, T35};
  assign T35 = T8[2'h2:2'h2];
  assign T36 = 8'h0 - T122;
  assign T122 = {7'h0, T37};
  assign T37 = T8[2'h3:2'h3];
  assign T38 = {T44, T39};
  assign T39 = {T42, T40};
  assign T40 = 8'h0 - T123;
  assign T123 = {7'h0, T41};
  assign T41 = T8[3'h4:3'h4];
  assign T42 = 8'h0 - T124;
  assign T124 = {7'h0, T43};
  assign T43 = T8[3'h5:3'h5];
  assign T44 = {T47, T45};
  assign T45 = 8'h0 - T125;
  assign T125 = {7'h0, T46};
  assign T46 = T8[3'h6:3'h6];
  assign T47 = 8'h0 - T126;
  assign T126 = {7'h0, T48};
  assign T48 = T8[3'h7:3'h7];
  assign T49 = wmask & out;
  assign out = T118 ? adder_out : T50;
  assign T50 = T112 ? T111 : T51;
  assign T51 = T110 ? T109 : T52;
  assign T52 = T108 ? T107 : T53;
  assign T53 = T69 ? io_lhs : T54;
  assign T54 = T68 ? T64 : T55;
  assign T55 = T63 ? T60 : T56;
  assign T56 = T59 ? T57 : io_rhs;
  assign T57 = {T58, T58};
  assign T58 = io_rhs[5'h1f:1'h0];
  assign T59 = T17 == 2'h2;
  assign T60 = {T61, T61};
  assign T61 = {T62, T62};
  assign T62 = io_rhs[4'hf:1'h0];
  assign T63 = T17 == 2'h1;
  assign T64 = {T65, T65};
  assign T65 = {T66, T66};
  assign T66 = {T67, T67};
  assign T67 = io_rhs[3'h7:1'h0];
  assign T68 = T17 == 2'h0;
  assign T69 = less ? min : max;
  assign max = T71 | T70;
  assign T70 = io_cmd == 5'hf;
  assign T71 = io_cmd == 5'hd;
  assign min = T73 | T72;
  assign T72 = io_cmd == 5'he;
  assign T73 = io_cmd == 5'hc;
  assign less = T106 ? lt : T74;
  assign T74 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T80 ? T79 : T75;
  assign T75 = rhs[6'h3f:6'h3f];
  assign rhs = T78 ? T76 : io_rhs;
  assign T76 = {T77, T77};
  assign T77 = io_rhs[5'h1f:1'h0];
  assign T78 = T17 == 2'h2;
  assign T79 = rhs[5'h1f:5'h1f];
  assign T80 = word & T81;
  assign T81 = T82 ^ 1'h1;
  assign T82 = io_addr[2'h2:2'h2];
  assign word = T84 | T83;
  assign T83 = io_typ == 3'h4;
  assign T84 = T86 | T85;
  assign T85 = io_typ == 3'h0;
  assign T86 = T88 | T87;
  assign T87 = io_typ == 3'h6;
  assign T88 = io_typ == 3'h2;
  assign cmp_lhs = T91 ? T90 : T89;
  assign T89 = io_lhs[6'h3f:6'h3f];
  assign T90 = io_lhs[5'h1f:5'h1f];
  assign T91 = word & T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = io_addr[2'h2:2'h2];
  assign sgned = T95 | T94;
  assign T94 = io_cmd == 5'hd;
  assign T95 = io_cmd == 5'hc;
  assign lt = word ? T104 : T96;
  assign T96 = lt_hi | T97;
  assign T97 = eq_hi & lt_lo;
  assign lt_lo = T99 < T98;
  assign T98 = rhs[5'h1f:1'h0];
  assign T99 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T101 == T100;
  assign T100 = rhs[6'h3f:6'h20];
  assign T101 = io_lhs[6'h3f:6'h20];
  assign lt_hi = T103 < T102;
  assign T102 = rhs[6'h3f:6'h20];
  assign T103 = io_lhs[6'h3f:6'h20];
  assign T104 = T105 ? lt_hi : lt_lo;
  assign T105 = io_addr[2'h2:2'h2];
  assign T106 = cmp_lhs == cmp_rhs;
  assign T107 = io_lhs ^ rhs;
  assign T108 = io_cmd == 5'h9;
  assign T109 = io_lhs | rhs;
  assign T110 = io_cmd == 5'ha;
  assign T111 = io_lhs & rhs;
  assign T112 = io_cmd == 5'hb;
  assign adder_out = T116 + T113;
  assign T113 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T127;
  assign T127 = {32'h0, T114};
  assign T114 = T115 << 5'h1f;
  assign T115 = io_addr[2'h2:2'h2];
  assign T116 = T117;
  assign T117 = io_lhs & mask;
  assign T118 = io_cmd == 5'h8;
endmodule

module LockingArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_addr_beat,
    input [25:0] io_in_1_bits_addr_block,
    input [1:0] io_in_1_bits_client_xact_id,
    input  io_in_1_bits_voluntary,
    input [2:0] io_in_1_bits_r_type,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_addr_beat,
    input [25:0] io_in_0_bits_addr_block,
    input [1:0] io_in_0_bits_client_xact_id,
    input  io_in_0_bits_voluntary,
    input [2:0] io_in_0_bits_r_type,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_addr_beat,
    output[25:0] io_out_bits_addr_block,
    output[1:0] io_out_bits_client_xact_id,
    output io_out_bits_voluntary,
    output[2:0] io_out_bits_r_type,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire chosen;
  wire T0;
  wire choose;
  reg  lockIdx;
  wire T35;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg  locked;
  wire T36;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire[1:0] T17;
  reg [1:0] R18;
  wire[1:0] T37;
  wire[1:0] T19;
  wire[127:0] T20;
  wire T21;
  wire[2:0] T22;
  wire T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lockIdx = {1{$random}};
    locked = {1{$random}};
    R18 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = T0;
  assign T0 = locked ? lockIdx : choose;
  assign choose = io_in_0_valid == 1'h0;
  assign T35 = reset ? 1'h1 : T1;
  assign T1 = T4 ? T2 : lockIdx;
  assign T2 = T3 == 1'h0;
  assign T3 = io_in_0_ready & io_in_0_valid;
  assign T4 = T6 & T5;
  assign T5 = locked ^ 1'h1;
  assign T6 = T12 & T7;
  assign T7 = T9 | T8;
  assign T8 = 3'h2 == io_out_bits_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h1 == io_out_bits_r_type;
  assign T11 = 3'h0 == io_out_bits_r_type;
  assign T12 = io_out_ready & io_out_valid;
  assign T36 = reset ? 1'h0 : T13;
  assign T13 = T15 ? 1'h0 : T14;
  assign T14 = T4 ? 1'h1 : locked;
  assign T15 = T12 & T16;
  assign T16 = T17 == 2'h0;
  assign T17 = R18 + 2'h1;
  assign T37 = reset ? 2'h0 : T19;
  assign T19 = T6 ? T17 : R18;
  assign io_out_bits_data = T20;
  assign T20 = T21 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T21 = chosen;
  assign io_out_bits_r_type = T22;
  assign T22 = T21 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign io_out_bits_voluntary = T23;
  assign T23 = T21 ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign io_out_bits_client_xact_id = T24;
  assign T24 = T21 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr_block = T25;
  assign T25 = T21 ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign io_out_bits_addr_beat = T26;
  assign T26 = T21 ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign io_out_valid = T27;
  assign T27 = T21 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = locked ? T30 : 1'h1;
  assign T30 = lockIdx == 1'h0;
  assign io_in_1_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = locked ? T34 : T33;
  assign T33 = io_in_0_valid ^ 1'h1;
  assign T34 = lockIdx == 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      lockIdx <= 1'h1;
    end else if(T4) begin
      lockIdx <= T2;
    end
    if(reset) begin
      locked <= 1'h0;
    end else if(T15) begin
      locked <= 1'h0;
    end else if(T4) begin
      locked <= 1'h1;
    end
    if(reset) begin
      R18 <= 2'h0;
    end else if(T6) begin
      R18 <= T17;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input [39:0] io_cpu_req_bits_addr,
    input [8:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_kill,
    input  io_cpu_req_bits_phys,
    input [63:0] io_cpu_req_bits_data,
    output io_cpu_resp_valid,
    output[39:0] io_cpu_resp_bits_addr,
    output[8:0] io_cpu_resp_bits_tag,
    output[4:0] io_cpu_resp_bits_cmd,
    output[2:0] io_cpu_resp_bits_typ,
    output[63:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data_word_bypass,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[8:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_invalidate_lr,
    output io_cpu_ordered,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[26:0] io_ptw_req_bits_addr,
    output[1:0] io_ptw_req_bits_prv,
    output io_ptw_req_bits_store,
    output io_ptw_req_bits_fetch,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [19:0] io_ptw_resp_bits_pte_ppn,
    input [2:0] io_ptw_resp_bits_pte_reserved_for_software,
    input  io_ptw_resp_bits_pte_d,
    input  io_ptw_resp_bits_pte_r,
    input [3:0] io_ptw_resp_bits_pte_typ,
    input  io_ptw_resp_bits_pte_v,
    input  io_ptw_status_sd,
    input [30:0] io_ptw_status_zero2,
    input  io_ptw_status_sd_rv32,
    input [8:0] io_ptw_status_zero1,
    input [4:0] io_ptw_status_vm,
    input  io_ptw_status_mprv,
    input [1:0] io_ptw_status_xs,
    input [1:0] io_ptw_status_fs,
    input [1:0] io_ptw_status_prv3,
    input  io_ptw_status_ie3,
    input [1:0] io_ptw_status_prv2,
    input  io_ptw_status_ie2,
    input [1:0] io_ptw_status_prv1,
    input  io_ptw_status_ie1,
    input [1:0] io_ptw_status_prv,
    input  io_ptw_status_ie,
    input  io_ptw_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[25:0] io_mem_acquire_bits_addr_block,
    output[1:0] io_mem_acquire_bits_client_xact_id,
    output[1:0] io_mem_acquire_bits_addr_beat,
    output io_mem_acquire_bits_is_builtin_type,
    output[2:0] io_mem_acquire_bits_a_type,
    output[16:0] io_mem_acquire_bits_union,
    output[127:0] io_mem_acquire_bits_data,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_addr_beat,
    input [1:0] io_mem_grant_bits_client_xact_id,
    input [2:0] io_mem_grant_bits_manager_xact_id,
    input  io_mem_grant_bits_is_builtin_type,
    input [3:0] io_mem_grant_bits_g_type,
    input [127:0] io_mem_grant_bits_data,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [25:0] io_mem_probe_bits_addr_block,
    input [1:0] io_mem_probe_bits_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_addr_beat,
    output[25:0] io_mem_release_bits_addr_block,
    output[1:0] io_mem_release_bits_client_xact_id,
    output io_mem_release_bits_voluntary,
    output[2:0] io_mem_release_bits_r_type,
    output[127:0] io_mem_release_bits_data
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  reg  R4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg [63:0] s2_req_data;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg  s1_replay;
  wire T416;
  wire T20;
  wire T21;
  wire s1_write;
  wire T22;
  wire T23;
  reg [4:0] s1_req_cmd;
  wire[4:0] T24;
  wire[4:0] T25;
  wire[4:0] T26;
  reg [4:0] s2_req_cmd;
  wire[4:0] T27;
  wire s2_recycle;
  wire T28;
  reg  s2_recycle_next;
  wire T417;
  wire T29;
  wire T30;
  reg  s1_valid;
  wire T418;
  wire T31;
  wire s2_recycle_ecc;
  wire s2_data_correctable;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire s2_word_idx;
  reg [39:0] s2_req_addr;
  wire[39:0] T36;
  wire[39:0] T419;
  wire[31:0] s1_addr;
  wire[11:0] T37;
  reg [39:0] s1_req_addr;
  wire[39:0] T38;
  wire[39:0] T39;
  wire[39:0] T40;
  wire[39:0] T41;
  wire[39:0] T42;
  wire[39:0] T420;
  wire[31:0] T43;
  wire[25:0] T44;
  wire[39:0] T421;
  wire[31:0] T45;
  wire[25:0] T46;
  wire T47;
  wire[1:0] T48;
  wire T49;
  wire s2_hit;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  reg [1:0] s2_hit_state_state;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire s2_tag_match;
  reg  s2_tag_match_way;
  wire T82;
  wire s1_tag_match_way;
  wire T83;
  wire T84;
  wire T85;
  wire s1_tag_eq_way;
  wire T86;
  wire[19:0] T87;
  wire T88;
  wire s2_replay;
  wire T89;
  reg  R90;
  wire T422;
  reg  s2_valid;
  wire T423;
  wire s1_valid_masked;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  reg  s1_clk_en;
  reg [63:0] s1_req_data;
  wire[63:0] T96;
  wire[63:0] T97;
  wire[63:0] T98;
  wire T99;
  reg  s1_recycled;
  wire T424;
  wire T100;
  wire[63:0] T425;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[6:0] T101;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T102;
  wire[63:0] T103;
  wire[127:0] s2_data_0;
  wire[127:0] T104;
  wire[127:0] T105;
  reg [63:0] R106;
  wire[63:0] T426;
  wire[127:0] T107;
  wire[127:0] T427;
  wire[127:0] T108;
  wire T109;
  wire T110;
  reg [63:0] R111;
  wire[63:0] T112;
  wire[63:0] T113;
  wire[63:0] T114;
  wire[127:0] T428;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T115;
  wire[63:0] T116;
  wire[63:0] T117;
  reg [63:0] s4_req_data;
  wire[63:0] T118;
  wire T119;
  reg  s3_valid;
  wire T429;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire s2_sc_fail;
  wire T130;
  wire s2_lrsc_addr_match;
  wire T131;
  wire[33:0] T132;
  reg [33:0] lrsc_addr;
  wire[33:0] T133;
  wire[33:0] T134;
  wire T135;
  wire s2_lr;
  wire T136;
  wire T137;
  wire s2_valid_masked;
  wire T138;
  wire T139;
  wire s2_nack;
  wire s2_nack_miss;
  wire T140;
  wire T141;
  wire T142;
  wire s2_nack_victim;
  reg  s2_nack_hit;
  wire T143;
  wire s1_nack;
  wire T144;
  wire T145;
  wire T146;
  wire[5:0] T147;
  wire T148;
  wire T149;
  wire lrsc_valid;
  reg [4:0] lrsc_count;
  wire[4:0] T430;
  wire[4:0] T150;
  wire[4:0] T151;
  wire[4:0] T152;
  wire[4:0] T153;
  wire[4:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire s2_sc;
  wire T158;
  wire T159;
  reg [63:0] s3_req_data;
  wire[63:0] T431;
  wire[127:0] T160;
  wire[127:0] T432;
  wire[63:0] T161;
  wire[127:0] T162;
  wire[127:0] T433;
  wire[127:0] s2_data_corrected;
  wire[127:0] T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  reg [4:0] s3_req_cmd;
  wire[4:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[36:0] T185;
  reg [39:0] s3_req_addr;
  wire[39:0] T186;
  wire[36:0] T434;
  wire[28:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[36:0] T198;
  wire[36:0] T435;
  wire[28:0] T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  reg [4:0] s4_req_cmd;
  wire[4:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire[36:0] T216;
  reg [39:0] s4_req_addr;
  wire[39:0] T217;
  wire[36:0] T436;
  wire[28:0] T218;
  reg  s4_valid;
  wire T437;
  wire T219;
  reg  s2_store_bypass;
  wire T220;
  wire T221;
  reg [2:0] s2_req_typ;
  wire[2:0] T222;
  reg [2:0] s1_req_typ;
  wire[2:0] T223;
  wire[2:0] T224;
  wire[2:0] T225;
  wire[5:0] T438;
  wire[127:0] T226;
  wire[1:0] rowWMask;
  wire rowIdx;
  wire T227;
  wire[11:0] T439;
  reg  s3_way;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[11:0] T440;
  wire[11:0] T441;
  wire[11:0] T442;
  wire[127:0] T241;
  wire[127:0] T242;
  wire[63:0] wdata_encoded_0;
  wire[63:0] wdata_encoded_1;
  wire[5:0] T443;
  wire[33:0] T243;
  wire[5:0] T444;
  wire[33:0] T244;
  reg  s1_req_phys;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  reg  s2_req_phys;
  wire T250;
  wire[27:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire s1_readwrite;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire s1_read;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire cache_pass;
  wire T269;
  reg  s2_killed;
  wire T270;
  wire T445;
  wire[1:0] T271;
  wire[1:0] s2_replaced_way_en;
  reg  R272;
  wire T273;
  wire[1:0] T446;
  wire[1:0] T274;
  reg [1:0] s2_repl_meta_coh_state;
  wire[1:0] T275;
  wire[1:0] T276;
  wire[19:0] T277;
  reg [19:0] s2_repl_meta_tag;
  wire[19:0] T278;
  wire[19:0] T279;
  reg  s2_req_kill;
  wire T280;
  reg  s1_req_kill;
  wire T281;
  wire T282;
  wire T283;
  reg [8:0] s2_req_tag;
  wire[8:0] T284;
  reg [8:0] s1_req_tag;
  wire[8:0] T285;
  wire[8:0] T286;
  wire[8:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire misaligned;
  wire[39:0] T324;
  wire[39:0] T447;
  wire[2:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[1:0] T328;
  wire T329;
  wire T330;
  wire[63:0] T331;
  wire[63:0] uncache_resp_bits_store_data;
  wire[63:0] cache_resp_bits_store_data;
  wire[63:0] T332;
  wire[31:0] T333;
  wire[31:0] T334;
  wire[31:0] T335;
  wire T336;
  wire[31:0] T337;
  wire[31:0] T338;
  wire[31:0] T339;
  wire[31:0] T448;
  wire T340;
  wire T341;
  wire T342;
  wire[2:0] T343;
  wire T344;
  wire[1:0] T345;
  wire T346;
  wire uncache_resp_bits_has_data;
  wire cache_resp_bits_has_data;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire uncache_resp_bits_replay;
  wire cache_resp_bits_replay;
  wire T357;
  wire uncache_resp_bits_nack;
  wire cache_resp_bits_nack;
  wire T358;
  wire[63:0] T359;
  wire[63:0] uncache_resp_bits_data;
  wire[63:0] cache_resp_bits_data;
  wire[63:0] T360;
  wire[63:0] T449;
  wire[63:0] T361;
  wire[7:0] T362;
  wire[7:0] T363;
  wire[7:0] T364;
  wire[63:0] T365;
  wire[15:0] T366;
  wire[15:0] T367;
  wire[63:0] T368;
  wire[31:0] T369;
  wire[31:0] T370;
  wire[31:0] T371;
  wire T372;
  wire[31:0] T373;
  wire[31:0] T374;
  wire[31:0] T375;
  wire[31:0] T450;
  wire T376;
  wire T377;
  wire T378;
  wire[15:0] T379;
  wire T380;
  wire[47:0] T381;
  wire[47:0] T382;
  wire[47:0] T383;
  wire[47:0] T451;
  wire T384;
  wire T385;
  wire T386;
  wire[7:0] T387;
  wire T388;
  wire[55:0] T389;
  wire[55:0] T390;
  wire[55:0] T391;
  wire[55:0] T452;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[2:0] T396;
  wire[2:0] uncache_resp_bits_typ;
  wire[2:0] cache_resp_bits_typ;
  wire[4:0] T397;
  wire[4:0] uncache_resp_bits_cmd;
  wire[4:0] cache_resp_bits_cmd;
  wire[8:0] T398;
  wire[8:0] uncache_resp_bits_tag;
  wire[8:0] cache_resp_bits_tag;
  wire[39:0] T399;
  wire[39:0] uncache_resp_bits_addr;
  wire[39:0] cache_resp_bits_addr;
  wire T400;
  wire uncache_resp_valid;
  wire cache_resp_valid;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  reg  block_miss;
  wire T453;
  wire T414;
  wire T415;
  wire wb_io_req_ready;
  wire wb_io_meta_read_valid;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_data_req_valid;
  wire wb_io_data_req_bits_way_en;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_release_valid;
  wire[1:0] wb_io_release_bits_addr_beat;
  wire[25:0] wb_io_release_bits_addr_block;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire wb_io_release_bits_voluntary;
  wire[2:0] wb_io_release_bits_r_type;
  wire[127:0] wb_io_release_bits_data;
  wire prober_io_req_ready;
  wire prober_io_rep_valid;
  wire[1:0] prober_io_rep_bits_addr_beat;
  wire[25:0] prober_io_rep_bits_addr_block;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire prober_io_rep_bits_voluntary;
  wire[2:0] prober_io_rep_bits_r_type;
  wire[127:0] prober_io_rep_bits_data;
  wire prober_io_meta_read_valid;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_write_valid;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire prober_io_meta_write_bits_way_en;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire prober_io_wb_req_valid;
  wire[1:0] prober_io_wb_req_bits_addr_beat;
  wire[25:0] prober_io_wb_req_bits_addr_block;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire prober_io_wb_req_bits_voluntary;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire[127:0] prober_io_wb_req_bits_data;
  wire prober_io_wb_req_bits_way_en;
  wire meta_io_read_ready;
  wire meta_io_write_ready;
  wire[19:0] meta_io_resp_0_tag;
  wire[1:0] meta_io_resp_0_coh_state;
  wire metaReadArb_io_in_4_ready;
  wire metaReadArb_io_in_3_ready;
  wire metaReadArb_io_in_2_ready;
  wire metaReadArb_io_in_1_ready;
  wire metaReadArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  wire metaWriteArb_io_in_1_ready;
  wire metaWriteArb_io_in_0_ready;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire metaWriteArb_io_out_bits_way_en;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire data_io_write_ready;
  wire[127:0] data_io_resp_0;
  wire readArb_io_in_3_ready;
  wire readArb_io_in_2_ready;
  wire readArb_io_in_1_ready;
  wire readArb_io_out_valid;
  wire readArb_io_out_bits_way_en;
  wire[11:0] readArb_io_out_bits_addr;
  wire writeArb_io_in_1_ready;
  wire writeArb_io_out_valid;
  wire writeArb_io_out_bits_way_en;
  wire[11:0] writeArb_io_out_bits_addr;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] amoalu_io_out;
  wire releaseArb_io_in_1_ready;
  wire releaseArb_io_in_0_ready;
  wire releaseArb_io_out_valid;
  wire[1:0] releaseArb_io_out_bits_addr_beat;
  wire[25:0] releaseArb_io_out_bits_addr_block;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire releaseArb_io_out_bits_voluntary;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire[127:0] releaseArb_io_out_bits_data;
  wire FlowThroughSerializer_io_in_ready;
  wire FlowThroughSerializer_io_out_valid;
  wire[1:0] FlowThroughSerializer_io_out_bits_addr_beat;
  wire[1:0] FlowThroughSerializer_io_out_bits_client_xact_id;
  wire[2:0] FlowThroughSerializer_io_out_bits_manager_xact_id;
  wire FlowThroughSerializer_io_out_bits_is_builtin_type;
  wire[3:0] FlowThroughSerializer_io_out_bits_g_type;
  wire[127:0] FlowThroughSerializer_io_out_bits_data;
  wire wbArb_io_in_1_ready;
  wire wbArb_io_in_0_ready;
  wire wbArb_io_out_valid;
  wire[1:0] wbArb_io_out_bits_addr_beat;
  wire[25:0] wbArb_io_out_bits_addr_block;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire wbArb_io_out_bits_voluntary;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire[127:0] wbArb_io_out_bits_data;
  wire wbArb_io_out_bits_way_en;
  wire dtlb_io_req_ready;
  wire dtlb_io_resp_miss;
  wire[19:0] dtlb_io_resp_ppn;
  wire dtlb_io_resp_xcpt_ld;
  wire dtlb_io_resp_xcpt_st;
  wire dtlb_io_ptw_req_valid;
  wire[26:0] dtlb_io_ptw_req_bits_addr;
  wire[1:0] dtlb_io_ptw_req_bits_prv;
  wire dtlb_io_ptw_req_bits_store;
  wire dtlb_io_ptw_req_bits_fetch;
  wire mshrs_io_req_ready;
  wire mshrs_io_resp_valid;
  wire[39:0] mshrs_io_resp_bits_addr;
  wire[8:0] mshrs_io_resp_bits_tag;
  wire[4:0] mshrs_io_resp_bits_cmd;
  wire[2:0] mshrs_io_resp_bits_typ;
  wire[63:0] mshrs_io_resp_bits_data;
  wire mshrs_io_resp_bits_nack;
  wire mshrs_io_resp_bits_replay;
  wire mshrs_io_resp_bits_has_data;
  wire[63:0] mshrs_io_resp_bits_store_data;
  wire mshrs_io_secondary_miss;
  wire mshrs_io_mem_req_valid;
  wire[25:0] mshrs_io_mem_req_bits_addr_block;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[1:0] mshrs_io_mem_req_bits_addr_beat;
  wire mshrs_io_mem_req_bits_is_builtin_type;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[16:0] mshrs_io_mem_req_bits_union;
  wire[127:0] mshrs_io_mem_req_bits_data;
  wire mshrs_io_refill_way_en;
  wire[11:0] mshrs_io_refill_addr;
  wire mshrs_io_meta_read_valid;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire mshrs_io_meta_write_bits_way_en;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire mshrs_io_replay_valid;
  wire[39:0] mshrs_io_replay_bits_addr;
  wire[8:0] mshrs_io_replay_bits_tag;
  wire[4:0] mshrs_io_replay_bits_cmd;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire mshrs_io_replay_bits_kill;
  wire mshrs_io_replay_bits_phys;
  wire[63:0] mshrs_io_replay_bits_data;
  wire mshrs_io_wb_req_valid;
  wire[1:0] mshrs_io_wb_req_bits_addr_beat;
  wire[25:0] mshrs_io_wb_req_bits_addr_block;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire mshrs_io_wb_req_bits_voluntary;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire[127:0] mshrs_io_wb_req_bits_data;
  wire mshrs_io_wb_req_bits_way_en;
  wire mshrs_io_probe_rdy;
  wire mshrs_io_fence_rdy;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    R4 = {1{$random}};
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s2_recycle_next = {1{$random}};
    s1_valid = {1{$random}};
    s2_req_addr = {2{$random}};
    s1_req_addr = {2{$random}};
    s2_hit_state_state = {1{$random}};
    s2_tag_match_way = {1{$random}};
    R90 = {1{$random}};
    s2_valid = {1{$random}};
    s1_clk_en = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R106 = {2{$random}};
    R111 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_data = {2{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    s2_killed = {1{$random}};
    R272 = {1{$random}};
    s2_repl_meta_coh_state = {1{$random}};
    s2_repl_meta_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    block_miss = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = T3 ^ 1'h1;
  assign T3 = R4 & io_cpu_resp_valid;
  assign T5 = T6 | io_cpu_xcpt_pf_st;
  assign T6 = T7 | io_cpu_xcpt_pf_ld;
  assign T7 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T8 = writeArb_io_in_1_ready | T9;
  assign T9 = T10 ^ 1'h1;
  assign T10 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T14 : T11;
  assign T11 = T13 | T12;
  assign T12 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T13 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T14 = T16 | T15;
  assign T15 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T16 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T17 = T99 ? s1_req_data : T18;
  assign T18 = T21 ? T19 : s2_req_data;
  assign T19 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T416 = reset ? 1'h0 : T20;
  assign T20 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T21 = s1_clk_en & s1_write;
  assign s1_write = T93 | T22;
  assign T22 = T92 | T23;
  assign T23 = s1_req_cmd == 5'h4;
  assign T24 = s2_recycle ? s2_req_cmd : T25;
  assign T25 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T26;
  assign T26 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T27 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T28;
  assign T28 = s2_recycle_ecc | s2_recycle_next;
  assign T417 = reset ? 1'h0 : T29;
  assign T29 = T30 ? s2_recycle_ecc : s2_recycle_next;
  assign T30 = s1_valid | s1_replay;
  assign T418 = reset ? 1'h0 : T31;
  assign T31 = io_cpu_req_ready & io_cpu_req_valid;
  assign s2_recycle_ecc = T49 & s2_data_correctable;
  assign s2_data_correctable = T47 & T32;
  assign T32 = T33 - 1'h1;
  assign T33 = 1'h1 << T34;
  assign T34 = T35 + 1'h1;
  assign T35 = s2_word_idx - s2_word_idx;
  assign s2_word_idx = s2_req_addr[2'h3:2'h3];
  assign T36 = s1_clk_en ? T419 : s2_req_addr;
  assign T419 = {8'h0, s1_addr};
  assign s1_addr = {dtlb_io_resp_ppn, T37};
  assign T37 = s1_req_addr[4'hb:1'h0];
  assign T38 = s2_recycle ? s2_req_addr : T39;
  assign T39 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T40;
  assign T40 = prober_io_meta_read_valid ? T421 : T41;
  assign T41 = wb_io_meta_read_valid ? T420 : T42;
  assign T42 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T420 = {8'h0, T43};
  assign T43 = T44 << 3'h6;
  assign T44 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T421 = {8'h0, T45};
  assign T45 = T46 << 3'h6;
  assign T46 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T47 = T48 >> s2_word_idx;
  assign T48 = 2'h0;
  assign T49 = T88 & s2_hit;
  assign s2_hit = T61 & T50;
  assign T50 = s2_hit_state_state == T51;
  assign T51 = T52;
  assign T52 = T53 ? 2'h3 : s2_hit_state_state;
  assign T53 = T57 | T54;
  assign T54 = T56 | T55;
  assign T55 = s2_req_cmd == 5'h4;
  assign T56 = s2_req_cmd[2'h3:2'h3];
  assign T57 = T59 | T58;
  assign T58 = s2_req_cmd == 5'h7;
  assign T59 = s2_req_cmd == 5'h1;
  assign T60 = s1_clk_en ? meta_io_resp_0_coh_state : s2_hit_state_state;
  assign T61 = s2_tag_match & T62;
  assign T62 = T71 ? T68 : T63;
  assign T63 = T65 | T64;
  assign T64 = 2'h3 == s2_hit_state_state;
  assign T65 = T67 | T66;
  assign T66 = 2'h2 == s2_hit_state_state;
  assign T67 = 2'h1 == s2_hit_state_state;
  assign T68 = T70 | T69;
  assign T69 = 2'h3 == s2_hit_state_state;
  assign T70 = 2'h2 == s2_hit_state_state;
  assign T71 = T73 | T72;
  assign T72 = s2_req_cmd == 5'h6;
  assign T73 = T75 | T74;
  assign T74 = s2_req_cmd == 5'h3;
  assign T75 = T79 | T76;
  assign T76 = T78 | T77;
  assign T77 = s2_req_cmd == 5'h4;
  assign T78 = s2_req_cmd[2'h3:2'h3];
  assign T79 = T81 | T80;
  assign T80 = s2_req_cmd == 5'h7;
  assign T81 = s2_req_cmd == 5'h1;
  assign s2_tag_match = s2_tag_match_way != 1'h0;
  assign T82 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T83;
  assign T83 = T85 & T84;
  assign T84 = meta_io_resp_0_coh_state != 2'h0;
  assign T85 = s1_tag_eq_way;
  assign s1_tag_eq_way = T86;
  assign T86 = meta_io_resp_0_tag == T87;
  assign T87 = s1_addr >> 4'hc;
  assign T88 = s2_valid | s2_replay;
  assign s2_replay = R90 & T89;
  assign T89 = s2_req_cmd != 5'h5;
  assign T422 = reset ? 1'h0 : s1_replay;
  assign T423 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T91;
  assign T91 = io_cpu_req_bits_kill ^ 1'h1;
  assign T92 = s1_req_cmd[2'h3:2'h3];
  assign T93 = T95 | T94;
  assign T94 = s1_req_cmd == 5'h7;
  assign T95 = s1_req_cmd == 5'h1;
  assign T96 = s2_recycle ? s2_req_data : T97;
  assign T97 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T98;
  assign T98 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T99 = s1_clk_en & s1_recycled;
  assign T424 = reset ? 1'h0 : T100;
  assign T100 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T425 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T428 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> T101;
  assign T101 = {s2_word_idx, 6'h0};
  assign s2_data_uncorrected = T102;
  assign T102 = {T114, T103};
  assign T103 = s2_data_0[6'h3f:1'h0];
  assign s2_data_0 = T104;
  assign T104 = T105;
  assign T105 = {R111, R106};
  assign T426 = T107[6'h3f:1'h0];
  assign T107 = T109 ? T108 : T427;
  assign T427 = {64'h0, R106};
  assign T108 = data_io_resp_0 >> 1'h0;
  assign T109 = s1_clk_en & T110;
  assign T110 = s1_tag_eq_way;
  assign T112 = T109 ? T113 : R111;
  assign T113 = data_io_resp_0 >> 7'h40;
  assign T114 = s2_data_0[7'h7f:7'h40];
  assign T428 = {64'h0, s2_store_bypass_data};
  assign T115 = T203 ? T116 : s2_store_bypass_data;
  assign T116 = T188 ? amoalu_io_out : T117;
  assign T117 = T174 ? s3_req_data : s4_req_data;
  assign T118 = T119 ? s3_req_data : s4_req_data;
  assign T119 = s3_valid & metaReadArb_io_out_valid;
  assign T429 = reset ? 1'h0 : T120;
  assign T120 = T128 & T121;
  assign T121 = T125 | T122;
  assign T122 = T124 | T123;
  assign T123 = s2_req_cmd == 5'h4;
  assign T124 = s2_req_cmd[2'h3:2'h3];
  assign T125 = T127 | T126;
  assign T126 = s2_req_cmd == 5'h7;
  assign T127 = s2_req_cmd == 5'h1;
  assign T128 = T158 & T129;
  assign T129 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T130;
  assign T130 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = lrsc_valid & T131;
  assign T131 = lrsc_addr == T132;
  assign T132 = s2_req_addr >> 3'h6;
  assign T133 = T135 ? T134 : lrsc_addr;
  assign T134 = s2_req_addr >> 3'h6;
  assign T135 = T136 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T136 = T137 | s2_replay;
  assign T137 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T138;
  assign T138 = s2_valid & T139;
  assign T139 = s2_nack ^ 1'h1;
  assign s2_nack = T142 | s2_nack_miss;
  assign s2_nack_miss = T141 & T140;
  assign T140 = mshrs_io_req_ready ^ 1'h1;
  assign T141 = s2_hit ^ 1'h1;
  assign T142 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T143 = T149 ? s1_nack : s2_nack_hit;
  assign s1_nack = T148 | T144;
  assign T144 = T146 & T145;
  assign T145 = prober_io_req_ready ^ 1'h1;
  assign T146 = T147 == prober_io_meta_write_bits_idx;
  assign T147 = s1_req_addr[4'hb:3'h6];
  assign T148 = T252 & dtlb_io_resp_miss;
  assign T149 = s1_valid | s1_replay;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T430 = reset ? 5'h0 : T150;
  assign T150 = io_cpu_invalidate_lr ? 5'h0 : T151;
  assign T151 = T157 ? 5'h0 : T152;
  assign T152 = T155 ? 5'h1f : T153;
  assign T153 = lrsc_valid ? T154 : lrsc_count;
  assign T154 = lrsc_count - 5'h1;
  assign T155 = T135 & T156;
  assign T156 = lrsc_valid ^ 1'h1;
  assign T157 = T136 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T158 = T159 | s2_replay;
  assign T159 = s2_valid_masked & s2_hit;
  assign T431 = T160[6'h3f:1'h0];
  assign T160 = T164 ? T162 : T432;
  assign T432 = {64'h0, T161};
  assign T161 = T164 ? s2_req_data : s3_req_data;
  assign T162 = s2_data_correctable ? s2_data_corrected : T433;
  assign T433 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T163;
  assign T163 = {T114, T103};
  assign T164 = T173 & T165;
  assign T165 = T166 | s2_data_correctable;
  assign T166 = T170 | T167;
  assign T167 = T169 | T168;
  assign T168 = s2_req_cmd == 5'h4;
  assign T169 = s2_req_cmd[2'h3:2'h3];
  assign T170 = T172 | T171;
  assign T171 = s2_req_cmd == 5'h7;
  assign T172 = s2_req_cmd == 5'h1;
  assign T173 = s2_valid | s2_replay;
  assign T174 = T183 & T175;
  assign T175 = T180 | T176;
  assign T176 = T179 | T177;
  assign T177 = s3_req_cmd == 5'h4;
  assign T178 = T164 ? s2_req_cmd : s3_req_cmd;
  assign T179 = s3_req_cmd[2'h3:2'h3];
  assign T180 = T182 | T181;
  assign T181 = s3_req_cmd == 5'h7;
  assign T182 = s3_req_cmd == 5'h1;
  assign T183 = s3_valid & T184;
  assign T184 = T434 == T185;
  assign T185 = s3_req_addr >> 2'h3;
  assign T186 = T164 ? s2_req_addr : s3_req_addr;
  assign T434 = {8'h0, T187};
  assign T187 = s1_addr >> 2'h3;
  assign T188 = T196 & T189;
  assign T189 = T193 | T190;
  assign T190 = T192 | T191;
  assign T191 = s2_req_cmd == 5'h4;
  assign T192 = s2_req_cmd[2'h3:2'h3];
  assign T193 = T195 | T194;
  assign T194 = s2_req_cmd == 5'h7;
  assign T195 = s2_req_cmd == 5'h1;
  assign T196 = T200 & T197;
  assign T197 = T435 == T198;
  assign T198 = s2_req_addr >> 2'h3;
  assign T435 = {8'h0, T199};
  assign T199 = s1_addr >> 2'h3;
  assign T200 = T202 & T201;
  assign T201 = s2_sc_fail ^ 1'h1;
  assign T202 = s2_valid_masked | s2_replay;
  assign T203 = s1_clk_en & T204;
  assign T204 = T219 | T205;
  assign T205 = T214 & T206;
  assign T206 = T211 | T207;
  assign T207 = T210 | T208;
  assign T208 = s4_req_cmd == 5'h4;
  assign T209 = T119 ? s3_req_cmd : s4_req_cmd;
  assign T210 = s4_req_cmd[2'h3:2'h3];
  assign T211 = T213 | T212;
  assign T212 = s4_req_cmd == 5'h7;
  assign T213 = s4_req_cmd == 5'h1;
  assign T214 = s4_valid & T215;
  assign T215 = T436 == T216;
  assign T216 = s4_req_addr >> 2'h3;
  assign T217 = T119 ? s3_req_addr : s4_req_addr;
  assign T436 = {8'h0, T218};
  assign T218 = s1_addr >> 2'h3;
  assign T437 = reset ? 1'h0 : s3_valid;
  assign T219 = T188 | T174;
  assign T220 = T203 ? 1'h1 : T221;
  assign T221 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T222 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T223 = s2_recycle ? s2_req_typ : T224;
  assign T224 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T225;
  assign T225 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T438 = s2_req_addr[3'h5:1'h0];
  assign T226 = {s3_req_data, s3_req_data};
  assign rowWMask = 1'h1 << rowIdx;
  assign rowIdx = T227;
  assign T227 = s3_req_addr[2'h3:2'h3];
  assign T439 = s3_req_addr[4'hb:1'h0];
  assign T228 = T164 ? s2_tag_match_way : s3_way;
  assign T229 = T231 & T230;
  assign T230 = FlowThroughSerializer_io_out_bits_client_xact_id < 2'h2;
  assign T231 = FlowThroughSerializer_io_out_valid & T232;
  assign T232 = FlowThroughSerializer_io_out_bits_is_builtin_type ? T236 : T233;
  assign T233 = T235 | T234;
  assign T234 = 4'h1 == FlowThroughSerializer_io_out_bits_g_type;
  assign T235 = 4'h0 == FlowThroughSerializer_io_out_bits_g_type;
  assign T236 = T238 | T237;
  assign T237 = 4'h4 == FlowThroughSerializer_io_out_bits_g_type;
  assign T238 = 4'h5 == FlowThroughSerializer_io_out_bits_g_type;
  assign T239 = T240 | T8;
  assign T240 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T440 = s2_req_addr[4'hb:1'h0];
  assign T441 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T442 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T241 = T242;
  assign T242 = {wdata_encoded_1, wdata_encoded_0};
  assign wdata_encoded_0 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign wdata_encoded_1 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T443 = T243[3'h5:1'h0];
  assign T243 = s2_req_addr >> 3'h6;
  assign T444 = T244[3'h5:1'h0];
  assign T244 = io_cpu_req_bits_addr >> 3'h6;
  assign T245 = s2_recycle ? s2_req_phys : T246;
  assign T246 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T247;
  assign T247 = prober_io_meta_read_valid ? 1'h1 : T248;
  assign T248 = wb_io_meta_read_valid ? 1'h1 : T249;
  assign T249 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T250 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T251 = s1_req_addr >> 4'hc;
  assign T252 = T254 & T253;
  assign T253 = s1_req_phys ^ 1'h1;
  assign T254 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T258 | T255;
  assign T255 = T257 | T256;
  assign T256 = s1_req_cmd == 5'h3;
  assign T257 = s1_req_cmd == 5'h2;
  assign T258 = s1_read | s1_write;
  assign s1_read = T262 | T259;
  assign T259 = T261 | T260;
  assign T260 = s1_req_cmd == 5'h4;
  assign T261 = s1_req_cmd[2'h3:2'h3];
  assign T262 = T264 | T263;
  assign T263 = s1_req_cmd == 5'h7;
  assign T264 = T266 | T265;
  assign T265 = s1_req_cmd == 5'h6;
  assign T266 = s1_req_cmd == 5'h0;
  assign T267 = T8 & FlowThroughSerializer_io_out_valid;
  assign T268 = cache_pass ^ 1'h1;
  assign cache_pass = T269 | s2_replay;
  assign T269 = s2_valid | s2_killed;
  assign T270 = s1_valid & io_cpu_req_bits_kill;
  assign T445 = T271[1'h0:1'h0];
  assign T271 = s2_tag_match ? T446 : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R272;
  assign T273 = s1_clk_en ? 1'h0 : R272;
  assign T446 = {1'h0, s2_tag_match_way};
  assign T274 = s2_tag_match ? T276 : s2_repl_meta_coh_state;
  assign T275 = s1_clk_en ? meta_io_resp_0_coh_state : s2_repl_meta_coh_state;
  assign T276 = s2_hit_state_state;
  assign T277 = s2_tag_match ? T279 : s2_repl_meta_tag;
  assign T278 = s1_clk_en ? meta_io_resp_0_tag : s2_repl_meta_tag;
  assign T279 = s2_repl_meta_tag;
  assign T280 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T281 = s2_recycle ? s2_req_kill : T282;
  assign T282 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T283;
  assign T283 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T284 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T285 = s2_recycle ? s2_req_tag : T286;
  assign T286 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T287;
  assign T287 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T288 = s2_nack_hit ? 1'h0 : T289;
  assign T289 = T311 & T290;
  assign T290 = T298 | T291;
  assign T291 = T295 | T292;
  assign T292 = T294 | T293;
  assign T293 = s2_req_cmd == 5'h4;
  assign T294 = s2_req_cmd[2'h3:2'h3];
  assign T295 = T297 | T296;
  assign T296 = s2_req_cmd == 5'h7;
  assign T297 = s2_req_cmd == 5'h1;
  assign T298 = T308 | T299;
  assign T299 = T303 | T300;
  assign T300 = T302 | T301;
  assign T301 = s2_req_cmd == 5'h4;
  assign T302 = s2_req_cmd[2'h3:2'h3];
  assign T303 = T305 | T304;
  assign T304 = s2_req_cmd == 5'h7;
  assign T305 = T307 | T306;
  assign T306 = s2_req_cmd == 5'h6;
  assign T307 = s2_req_cmd == 5'h0;
  assign T308 = T310 | T309;
  assign T309 = s2_req_cmd == 5'h3;
  assign T310 = s2_req_cmd == 5'h2;
  assign T311 = s2_valid_masked & T312;
  assign T312 = s2_hit ^ 1'h1;
  assign T313 = io_mem_probe_valid & T314;
  assign T314 = lrsc_valid ^ 1'h1;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_probe_ready = T315;
  assign T315 = prober_io_req_ready & T316;
  assign T316 = lrsc_valid ^ 1'h1;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_ordered = T317;
  assign T317 = T319 & T318;
  assign T318 = s2_valid ^ 1'h1;
  assign T319 = mshrs_io_fence_rdy & T320;
  assign T320 = s1_valid ^ 1'h1;
  assign io_cpu_xcpt_pf_st = T321;
  assign T321 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T322;
  assign T322 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T323;
  assign T323 = s1_write & misaligned;
  assign misaligned = T324 != 40'h0;
  assign T324 = s1_req_addr & T447;
  assign T447 = {37'h0, T325};
  assign T325 = T326[2'h2:1'h0];
  assign T326 = T327 - 4'h1;
  assign T327 = 1'h1 << T328;
  assign T328 = s1_req_typ[1'h1:1'h0];
  assign io_cpu_xcpt_ma_ld = T329;
  assign T329 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T330;
  assign T330 = s1_replay & s1_read;
  assign io_cpu_resp_bits_store_data = T331;
  assign T331 = cache_pass ? cache_resp_bits_store_data : uncache_resp_bits_store_data;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign cache_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_data_word_bypass = T332;
  assign T332 = {T337, T333};
  assign T333 = T336 ? T335 : T334;
  assign T334 = s2_data_word[5'h1f:1'h0];
  assign T335 = s2_data_word[6'h3f:6'h20];
  assign T336 = s2_req_addr[2'h2:2'h2];
  assign T337 = T344 ? T339 : T338;
  assign T338 = s2_data_word[6'h3f:6'h20];
  assign T339 = 32'h0 - T448;
  assign T448 = {31'h0, T340};
  assign T340 = T342 & T341;
  assign T341 = T333[5'h1f:5'h1f];
  assign T342 = $signed(1'h0) <= $signed(T343);
  assign T343 = s2_req_typ;
  assign T344 = T345 == 2'h2;
  assign T345 = s2_req_typ[1'h1:1'h0];
  assign io_cpu_resp_bits_has_data = T346;
  assign T346 = cache_pass ? cache_resp_bits_has_data : uncache_resp_bits_has_data;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign cache_resp_bits_has_data = T347;
  assign T347 = T351 | T348;
  assign T348 = T350 | T349;
  assign T349 = s2_req_cmd == 5'h4;
  assign T350 = s2_req_cmd[2'h3:2'h3];
  assign T351 = T353 | T352;
  assign T352 = s2_req_cmd == 5'h7;
  assign T353 = T355 | T354;
  assign T354 = s2_req_cmd == 5'h6;
  assign T355 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_replay = T356;
  assign T356 = cache_pass ? cache_resp_bits_replay : uncache_resp_bits_replay;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign cache_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T357;
  assign T357 = cache_pass ? cache_resp_bits_nack : uncache_resp_bits_nack;
  assign uncache_resp_bits_nack = mshrs_io_resp_bits_nack;
  assign cache_resp_bits_nack = T358;
  assign T358 = s2_valid & s2_nack;
  assign io_cpu_resp_bits_data = T359;
  assign T359 = cache_pass ? cache_resp_bits_data : uncache_resp_bits_data;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign cache_resp_bits_data = T360;
  assign T360 = T361 | T449;
  assign T449 = {63'h0, s2_sc_fail};
  assign T361 = {T389, T362};
  assign T362 = s2_sc ? 8'h0 : T363;
  assign T363 = T388 ? T387 : T364;
  assign T364 = T365[3'h7:1'h0];
  assign T365 = {T381, T366};
  assign T366 = T380 ? T379 : T367;
  assign T367 = T368[4'hf:1'h0];
  assign T368 = {T373, T369};
  assign T369 = T372 ? T371 : T370;
  assign T370 = s2_data_word[5'h1f:1'h0];
  assign T371 = s2_data_word[6'h3f:6'h20];
  assign T372 = s2_req_addr[2'h2:2'h2];
  assign T373 = T378 ? T375 : T374;
  assign T374 = s2_data_word[6'h3f:6'h20];
  assign T375 = 32'h0 - T450;
  assign T450 = {31'h0, T376};
  assign T376 = T342 & T377;
  assign T377 = T369[5'h1f:5'h1f];
  assign T378 = T345 == 2'h2;
  assign T379 = T368[5'h1f:5'h10];
  assign T380 = s2_req_addr[1'h1:1'h1];
  assign T381 = T386 ? T383 : T382;
  assign T382 = T368[6'h3f:5'h10];
  assign T383 = 48'h0 - T451;
  assign T451 = {47'h0, T384};
  assign T384 = T342 & T385;
  assign T385 = T366[4'hf:4'hf];
  assign T386 = T345 == 2'h1;
  assign T387 = T365[4'hf:4'h8];
  assign T388 = s2_req_addr[1'h0:1'h0];
  assign T389 = T394 ? T391 : T390;
  assign T390 = T365[6'h3f:4'h8];
  assign T391 = 56'h0 - T452;
  assign T452 = {55'h0, T392};
  assign T392 = T342 & T393;
  assign T393 = T362[3'h7:3'h7];
  assign T394 = T395 | s2_sc;
  assign T395 = T345 == 2'h0;
  assign io_cpu_resp_bits_typ = T396;
  assign T396 = cache_pass ? cache_resp_bits_typ : uncache_resp_bits_typ;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign cache_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_cmd = T397;
  assign T397 = cache_pass ? cache_resp_bits_cmd : uncache_resp_bits_cmd;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_tag = T398;
  assign T398 = cache_pass ? cache_resp_bits_tag : uncache_resp_bits_tag;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign cache_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_addr = T399;
  assign T399 = cache_pass ? cache_resp_bits_addr : uncache_resp_bits_addr;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign cache_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_valid = T400;
  assign T400 = cache_pass ? cache_resp_valid : uncache_resp_valid;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign cache_resp_valid = T401;
  assign T401 = T403 & T402;
  assign T402 = s2_data_correctable ^ 1'h1;
  assign T403 = s2_replay | T404;
  assign T404 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T405;
  assign T405 = block_miss ? 1'h0 : T406;
  assign T406 = T413 ? 1'h0 : T407;
  assign T407 = T412 ? 1'h0 : T408;
  assign T408 = T409 == 1'h0;
  assign T409 = T411 & T410;
  assign T410 = io_cpu_req_bits_phys ^ 1'h1;
  assign T411 = dtlb_io_req_ready ^ 1'h1;
  assign T412 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T413 = readArb_io_in_3_ready ^ 1'h1;
  assign T453 = reset ? 1'h0 : T414;
  assign T414 = T415 & s2_nack_miss;
  assign T415 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_req_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_req_bits_data( wbArb_io_out_bits_data ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_release_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_release_bits_r_type( wb_io_release_bits_r_type ),
       .io_release_bits_data( wb_io_release_bits_data )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T313 ),
       .io_req_bits_addr_block( io_mem_probe_bits_addr_block ),
       .io_req_bits_p_type( io_mem_probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_rep_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( prober_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_block_state_state( s2_hit_state_state )
  );
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T288 ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag_match( s2_tag_match ),
       .io_req_bits_old_meta_tag( T277 ),
       .io_req_bits_old_meta_coh_state( T274 ),
       .io_req_bits_way_en( T445 ),
       .io_resp_ready( T268 ),
       .io_resp_valid( mshrs_io_resp_valid ),
       .io_resp_bits_addr( mshrs_io_resp_bits_addr ),
       .io_resp_bits_tag( mshrs_io_resp_bits_tag ),
       .io_resp_bits_cmd( mshrs_io_resp_bits_cmd ),
       .io_resp_bits_typ( mshrs_io_resp_bits_typ ),
       .io_resp_bits_data( mshrs_io_resp_bits_data ),
       .io_resp_bits_nack( mshrs_io_resp_bits_nack ),
       .io_resp_bits_replay( mshrs_io_resp_bits_replay ),
       .io_resp_bits_has_data( mshrs_io_resp_bits_has_data ),
       //.io_resp_bits_data_word_bypass(  )
       .io_resp_bits_store_data( mshrs_io_resp_bits_store_data ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( io_mem_acquire_ready ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr_block( mshrs_io_mem_req_bits_addr_block ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_addr_beat( mshrs_io_mem_req_bits_addr_beat ),
       .io_mem_req_bits_is_builtin_type( mshrs_io_mem_req_bits_is_builtin_type ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_union( mshrs_io_mem_req_bits_union ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_refill_way_en( mshrs_io_refill_way_en ),
       .io_refill_addr( mshrs_io_refill_addr ),
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_mem_grant_valid( T267 ),
       .io_mem_grant_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_mem_grant_bits_data( FlowThroughSerializer_io_out_bits_data ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_wb_req_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_wb_req_bits_data( mshrs_io_wb_req_bits_data ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T252 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T251 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_req_bits_store( s1_write ),
       .io_resp_miss( dtlb_io_resp_miss ),
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       //.io_resp_hit_idx(  )
       .io_ptw_req_ready( io_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dtlb_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dtlb_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dtlb_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dtlb_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( io_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_ptw_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( io_ptw_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( io_ptw_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( io_ptw_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( io_ptw_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( io_ptw_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( io_ptw_resp_bits_pte_v ),
       .io_ptw_status_sd( io_ptw_status_sd ),
       .io_ptw_status_zero2( io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( io_ptw_status_zero1 ),
       .io_ptw_status_vm( io_ptw_status_vm ),
       .io_ptw_status_mprv( io_ptw_status_mprv ),
       .io_ptw_status_xs( io_ptw_status_xs ),
       .io_ptw_status_fs( io_ptw_status_fs ),
       .io_ptw_status_prv3( io_ptw_status_prv3 ),
       .io_ptw_status_ie3( io_ptw_status_ie3 ),
       .io_ptw_status_prv2( io_ptw_status_prv2 ),
       .io_ptw_status_ie2( io_ptw_status_ie2 ),
       .io_ptw_status_prv1( io_ptw_status_prv1 ),
       .io_ptw_status_ie1( io_ptw_status_ie1 ),
       .io_ptw_status_prv( io_ptw_status_prv ),
       .io_ptw_status_ie( io_ptw_status_ie ),
       .io_ptw_invalidate( io_ptw_invalidate )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_0 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T444 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T443 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T241 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_2 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 1'h1 ),
       .io_in_3_bits_addr( T442 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 1'h1 ),
       .io_in_1_bits_addr( T441 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 1'h1 ),
       .io_in_0_bits_addr( T440 ),
       .io_out_ready( T239 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_3 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T229 ),
       .io_in_1_bits_way_en( mshrs_io_refill_way_en ),
       .io_in_1_bits_addr( mshrs_io_refill_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( FlowThroughSerializer_io_out_bits_data ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T439 ),
       .io_in_0_bits_wmask( rowWMask ),
       .io_in_0_bits_data( T226 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T438 ),
       .io_cmd( s2_req_cmd ),
       .io_typ( s2_req_typ ),
       .io_lhs( T425 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  LockingArbiter_0 releaseArb(.clk(clk), .reset(reset),
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr_beat( prober_io_rep_bits_addr_beat ),
       .io_in_1_bits_addr_block( prober_io_rep_bits_addr_block ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_voluntary( prober_io_rep_bits_voluntary ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr_beat( wb_io_release_bits_addr_beat ),
       .io_in_0_bits_addr_block( wb_io_release_bits_addr_block ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_voluntary( wb_io_release_bits_voluntary ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_out_ready( io_mem_release_ready ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr_beat( releaseArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( releaseArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( releaseArb_io_out_bits_voluntary ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type ),
       .io_out_bits_data( releaseArb_io_out_bits_data )
       //.io_chosen(  )
  );
  FlowThroughSerializer FlowThroughSerializer(
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_addr_beat( io_mem_grant_bits_addr_beat ),
       .io_in_bits_client_xact_id( io_mem_grant_bits_client_xact_id ),
       .io_in_bits_manager_xact_id( io_mem_grant_bits_manager_xact_id ),
       .io_in_bits_is_builtin_type( io_mem_grant_bits_is_builtin_type ),
       .io_in_bits_g_type( io_mem_grant_bits_g_type ),
       .io_in_bits_data( io_mem_grant_bits_data ),
       .io_out_ready( T8 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_addr_beat( FlowThroughSerializer_io_out_bits_addr_beat ),
       .io_out_bits_client_xact_id( FlowThroughSerializer_io_out_bits_client_xact_id ),
       .io_out_bits_manager_xact_id( FlowThroughSerializer_io_out_bits_manager_xact_id ),
       .io_out_bits_is_builtin_type( FlowThroughSerializer_io_out_bits_is_builtin_type ),
       .io_out_bits_g_type( FlowThroughSerializer_io_out_bits_g_type ),
       .io_out_bits_data( FlowThroughSerializer_io_out_bits_data )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_addr_beat( mshrs_io_wb_req_bits_addr_beat ),
       .io_in_1_bits_addr_block( mshrs_io_wb_req_bits_addr_block ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_voluntary( mshrs_io_wb_req_bits_voluntary ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_1_bits_data( mshrs_io_wb_req_bits_data ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_addr_beat( prober_io_wb_req_bits_addr_beat ),
       .io_in_0_bits_addr_block( prober_io_wb_req_bits_addr_block ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_voluntary( prober_io_wb_req_bits_voluntary ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_in_0_bits_data( prober_io_wb_req_bits_data ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_addr_beat( wbArb_io_out_bits_addr_beat ),
       .io_out_bits_addr_block( wbArb_io_out_bits_addr_block ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_voluntary( wbArb_io_out_bits_voluntary ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_out_bits_data( wbArb_io_out_bits_data ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "DCache exception occurred - cache response not killed.");
    $finish;
  end
// synthesis translate_on
`endif
    R4 <= T5;
    if(T99) begin
      s2_req_data <= s1_req_data;
    end else if(T21) begin
      s2_req_data <= T19;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T20;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T30) begin
      s2_recycle_next <= s2_recycle_ecc;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T31;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T419;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T421;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T420;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_hit_state_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(reset) begin
      R90 <= 1'h0;
    end else begin
      R90 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R106 <= T426;
    if(T109) begin
      R111 <= T113;
    end
    if(T203) begin
      s2_store_bypass_data <= T116;
    end
    if(T119) begin
      s4_req_data <= s3_req_data;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T120;
    end
    if(T135) begin
      lrsc_addr <= T134;
    end
    if(T149) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_invalidate_lr) begin
      lrsc_count <= 5'h0;
    end else if(T157) begin
      lrsc_count <= 5'h0;
    end else if(T155) begin
      lrsc_count <= 5'h1f;
    end else if(lrsc_valid) begin
      lrsc_count <= T154;
    end
    s3_req_data <= T431;
    if(T164) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T164) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T119) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T119) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T203) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T164) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    s2_killed <= T270;
    if(s1_clk_en) begin
      R272 <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_repl_meta_coh_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_repl_meta_tag <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T414;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [26:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_prv,
    input  io_in_1_bits_store,
    input  io_in_1_bits_fetch,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [26:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_prv,
    input  io_in_0_bits_store,
    input  io_in_0_bits_fetch,
    input  io_out_ready,
    output io_out_valid,
    output[26:0] io_out_bits_addr,
    output[1:0] io_out_bits_prv,
    output io_out_bits_store,
    output io_out_bits_fetch,
    output io_chosen
);

  wire chosen;
  wire choose;
  wire T0;
  wire T1;
  wire T2;
  reg  last_grant;
  wire T28;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire[26:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_chosen = chosen;
  assign chosen = choose;
  assign choose = T1 ? 1'h1 : T0;
  assign T0 = io_in_0_valid == 1'h0;
  assign T1 = io_in_1_valid & T2;
  assign T2 = last_grant < 1'h1;
  assign T28 = reset ? 1'h0 : T3;
  assign T3 = T4 ? chosen : last_grant;
  assign T4 = io_out_ready & io_out_valid;
  assign io_out_bits_fetch = T5;
  assign T5 = T6 ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T6 = chosen;
  assign io_out_bits_store = T7;
  assign T7 = T6 ? io_in_1_bits_store : io_in_0_bits_store;
  assign io_out_bits_prv = T8;
  assign T8 = T6 ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign io_out_bits_addr = T9;
  assign T9 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T6 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = T19 | T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = T17 | T15;
  assign T15 = io_in_1_valid & T16;
  assign T16 = last_grant < 1'h1;
  assign T17 = io_in_0_valid & T18;
  assign T18 = last_grant < 1'h0;
  assign T19 = last_grant < 1'h0;
  assign io_in_1_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T25 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T24 | io_in_0_valid;
  assign T24 = T17 | T15;
  assign T25 = T27 & T26;
  assign T26 = last_grant < 1'h1;
  assign T27 = T17 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 1'h0;
    end else if(T4) begin
      last_grant <= chosen;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [26:0] io_requestor_1_req_bits_addr,
    input [1:0] io_requestor_1_req_bits_prv,
    input  io_requestor_1_req_bits_store,
    input  io_requestor_1_req_bits_fetch,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[19:0] io_requestor_1_resp_bits_pte_ppn,
    output[2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
    output io_requestor_1_resp_bits_pte_d,
    output io_requestor_1_resp_bits_pte_r,
    output[3:0] io_requestor_1_resp_bits_pte_typ,
    output io_requestor_1_resp_bits_pte_v,
    output io_requestor_1_status_sd,
    output[30:0] io_requestor_1_status_zero2,
    output io_requestor_1_status_sd_rv32,
    output[8:0] io_requestor_1_status_zero1,
    output[4:0] io_requestor_1_status_vm,
    output io_requestor_1_status_mprv,
    output[1:0] io_requestor_1_status_xs,
    output[1:0] io_requestor_1_status_fs,
    output[1:0] io_requestor_1_status_prv3,
    output io_requestor_1_status_ie3,
    output[1:0] io_requestor_1_status_prv2,
    output io_requestor_1_status_ie2,
    output[1:0] io_requestor_1_status_prv1,
    output io_requestor_1_status_ie1,
    output[1:0] io_requestor_1_status_prv,
    output io_requestor_1_status_ie,
    output io_requestor_1_invalidate,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [26:0] io_requestor_0_req_bits_addr,
    input [1:0] io_requestor_0_req_bits_prv,
    input  io_requestor_0_req_bits_store,
    input  io_requestor_0_req_bits_fetch,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[19:0] io_requestor_0_resp_bits_pte_ppn,
    output[2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
    output io_requestor_0_resp_bits_pte_d,
    output io_requestor_0_resp_bits_pte_r,
    output[3:0] io_requestor_0_resp_bits_pte_typ,
    output io_requestor_0_resp_bits_pte_v,
    output io_requestor_0_status_sd,
    output[30:0] io_requestor_0_status_zero2,
    output io_requestor_0_status_sd_rv32,
    output[8:0] io_requestor_0_status_zero1,
    output[4:0] io_requestor_0_status_vm,
    output io_requestor_0_status_mprv,
    output[1:0] io_requestor_0_status_xs,
    output[1:0] io_requestor_0_status_fs,
    output[1:0] io_requestor_0_status_prv3,
    output io_requestor_0_status_ie3,
    output[1:0] io_requestor_0_status_prv2,
    output io_requestor_0_status_ie2,
    output[1:0] io_requestor_0_status_prv1,
    output io_requestor_0_status_ie1,
    output[1:0] io_requestor_0_status_prv,
    output io_requestor_0_status_ie,
    output io_requestor_0_invalidate,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    //output[8:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [8:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_status_sd,
    input [30:0] io_dpath_status_zero2,
    input  io_dpath_status_sd_rv32,
    input [8:0] io_dpath_status_zero1,
    input [4:0] io_dpath_status_vm,
    input  io_dpath_status_mprv,
    input [1:0] io_dpath_status_xs,
    input [1:0] io_dpath_status_fs,
    input [1:0] io_dpath_status_prv3,
    input  io_dpath_status_ie3,
    input [1:0] io_dpath_status_prv2,
    input  io_dpath_status_ie2,
    input [1:0] io_dpath_status_prv1,
    input  io_dpath_status_ie1,
    input [1:0] io_dpath_status_prv,
    input  io_dpath_status_ie
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T232;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  reg [1:0] count;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T22;
  wire pte_cache_hit;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[1:0] T26;
  reg  R27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire[1:0] T233;
  wire[1:0] T234;
  wire T235;
  wire[2:0] T36;
  wire T236;
  wire[1:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire T41;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  reg [2:0] R45;
  wire[2:0] T46;
  wire[2:0] T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire[5:0] T50;
  wire[1:0] T51;
  wire T52;
  wire[1:0] T237;
  wire T238;
  wire[1:0] T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire[2:0] T57;
  wire[2:0] T58;
  wire[2:0] T59;
  wire T60;
  wire T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[3:0] T70;
  wire T71;
  wire T72;
  reg  R73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  R78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[31:0] pte_addr;
  wire[28:0] T87;
  wire[28:0] T88;
  wire[8:0] vpn_idx;
  wire[8:0] T89;
  wire[8:0] T90;
  wire[8:0] T91;
  reg [26:0] r_req_addr;
  wire[26:0] T92;
  wire T93;
  wire[8:0] T94;
  wire[17:0] T95;
  wire T96;
  wire[1:0] T97;
  wire[8:0] T98;
  wire[26:0] T99;
  wire T100;
  reg [19:0] r_pte_ppn;
  wire[19:0] T101;
  wire[19:0] T102;
  wire[19:0] T103;
  wire[19:0] T104;
  wire[19:0] T105;
  wire T106;
  wire T107;
  wire set_dirty_bit;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  reg  r_req_store;
  wire T112;
  wire T113;
  wire T114;
  wire perm_ok;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  reg  r_req_fetch;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  reg [1:0] r_req_prv;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire[19:0] pte_cache_data;
  wire[19:0] T150;
  wire[19:0] T151;
  reg [19:0] T152 [2:0];
  wire[19:0] T153;
  wire T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire[19:0] T158;
  wire[19:0] T159;
  wire[19:0] T160;
  wire T161;
  wire[19:0] T162;
  wire[19:0] T163;
  wire T164;
  wire[31:0] T165;
  reg [31:0] T166 [2:0];
  wire[31:0] T167;
  wire T168;
  wire T169;
  wire[1:0] T170;
  wire T171;
  wire[31:0] T172;
  wire T173;
  wire[31:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire[2:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[63:0] T243;
  wire[29:0] T198;
  wire[29:0] T199;
  wire[5:0] T200;
  wire[4:0] T201;
  wire pte_wdata_v;
  wire[3:0] pte_wdata_typ;
  wire pte_wdata_r;
  wire[23:0] T202;
  wire[3:0] T203;
  wire pte_wdata_d;
  wire[2:0] pte_wdata_reserved_for_software;
  wire[19:0] pte_wdata_ppn;
  wire[4:0] T204;
  wire T205;
  wire[39:0] T244;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  reg  r_pte_v;
  wire T210;
  reg [3:0] r_pte_typ;
  wire[3:0] T211;
  reg  r_pte_r;
  wire T212;
  reg  r_pte_d;
  wire T213;
  reg [2:0] r_pte_reserved_for_software;
  wire[2:0] T214;
  wire[2:0] T215;
  wire[19:0] T245;
  wire[27:0] resp_ppn;
  wire[27:0] T216;
  wire[27:0] T217;
  wire[17:0] T218;
  wire[9:0] T219;
  wire[27:0] T220;
  wire[8:0] T221;
  wire[18:0] T222;
  wire T223;
  wire[1:0] T224;
  wire[27:0] r_resp_ppn;
  wire T225;
  wire resp_err;
  wire T226;
  wire T227;
  reg  r_req_dest;
  wire T228;
  wire resp_val;
  wire T229;
  wire[19:0] T246;
  wire T230;
  wire T231;
  wire arb_io_in_1_ready;
  wire arb_io_in_0_ready;
  wire arb_io_out_valid;
  wire[26:0] arb_io_out_bits_addr;
  wire[1:0] arb_io_out_bits_prv;
  wire arb_io_out_bits_store;
  wire arb_io_out_bits_fetch;
  wire arb_io_chosen;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    R27 = {1{$random}};
    R45 = {1{$random}};
    R73 = {1{$random}};
    R78 = {1{$random}};
    r_req_addr = {1{$random}};
    r_pte_ppn = {1{$random}};
    r_req_store = {1{$random}};
    r_req_fetch = {1{$random}};
    r_req_prv = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T152[initvar] = {1{$random}};
    for (initvar = 0; initvar < 3; initvar = initvar+1)
      T166[initvar] = {1{$random}};
    r_pte_v = {1{$random}};
    r_pte_typ = {1{$random}};
    r_pte_r = {1{$random}};
    r_pte_d = {1{$random}};
    r_pte_reserved_for_software = {1{$random}};
    r_req_dest = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
//  assign io_mem_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
  assign T0 = state == 3'h0;
  assign T232 = reset ? 3'h0 : T1;
  assign T1 = T197 ? 3'h0 : T2;
  assign T2 = T196 ? 3'h0 : T3;
  assign T3 = T195 ? 3'h1 : T4;
  assign T4 = T193 ? 3'h3 : T5;
  assign T5 = T191 ? 3'h4 : T6;
  assign T6 = T188 ? T187 : T7;
  assign T7 = T182 ? 3'h1 : T8;
  assign T8 = T181 ? 3'h6 : T9;
  assign T9 = T179 ? 3'h1 : T10;
  assign T10 = T176 ? 3'h2 : T11;
  assign T11 = T15 ? 3'h1 : T12;
  assign T12 = T13 ? 3'h1 : state;
  assign T13 = T14 & arb_io_out_valid;
  assign T14 = 3'h0 == state;
  assign T15 = T175 & T16;
  assign T16 = pte_cache_hit & T17;
  assign T17 = count < 2'h2;
  assign T18 = T182 ? T22 : T19;
  assign T19 = T15 ? T21 : T20;
  assign T20 = T14 ? 2'h0 : count;
  assign T21 = count + 2'h1;
  assign T22 = count + 2'h1;
  assign pte_cache_hit = T23 != 3'h0;
  assign T23 = T83 & T24;
  assign T24 = T25;
  assign T25 = {R78, T26};
  assign T26 = {R73, R27};
  assign T28 = T72 ? 1'h0 : T29;
  assign T29 = T30 ? 1'h1 : R27;
  assign T30 = T65 & T31;
  assign T31 = T32[1'h0:1'h0];
  assign T32 = 1'h1 << T33;
  assign T33 = T34;
  assign T34 = T64 ? T37 : T233;
  assign T233 = T236 ? 1'h0 : T234;
  assign T234 = T235 ? 1'h1 : 2'h2;
  assign T235 = T36[1'h1:1'h1];
  assign T36 = ~ T24;
  assign T236 = T36[1'h0:1'h0];
  assign T37 = T38[1'h1:1'h0];
  assign T38 = {T62, T39};
  assign T39 = T44 & T40;
  assign T40 = T41 - 1'h1;
  assign T41 = 1'h1 << T42;
  assign T42 = T43 + 2'h1;
  assign T43 = T62 - T62;
  assign T44 = R45 >> T62;
  assign T46 = T60 ? T47 : R45;
  assign T47 = T55 | T48;
  assign T48 = T54 ? 3'h0 : T49;
  assign T49 = T50[2'h2:1'h0];
  assign T50 = 3'h1 << T51;
  assign T51 = {1'h1, T52};
  assign T52 = T237[1'h1:1'h1];
  assign T237 = {T242, T238};
  assign T238 = T239[1'h1:1'h1];
  assign T239 = T241 | T240;
  assign T240 = T23[1'h1:1'h0];
  assign T241 = T23[2'h2:2'h2];
  assign T242 = T241 != 1'h0;
  assign T54 = T237[1'h0:1'h0];
  assign T55 = T57 & T56;
  assign T56 = ~ T49;
  assign T57 = T59 | T58;
  assign T58 = T52 ? 3'h0 : 3'h2;
  assign T59 = R45 & 3'h5;
  assign T60 = pte_cache_hit & T61;
  assign T61 = state == 3'h1;
  assign T62 = {1'h1, T63};
  assign T63 = R45[1'h1:1'h1];
  assign T64 = T24 == 3'h7;
  assign T65 = T67 & T66;
  assign T66 = pte_cache_hit ^ 1'h1;
  assign T67 = io_mem_resp_valid & T68;
  assign T68 = T71 & T69;
  assign T69 = T70 < 4'h2;
  assign T70 = io_mem_resp_bits_data[3'h4:1'h1];
  assign T71 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T72 = reset | io_dpath_invalidate;
  assign T74 = T72 ? 1'h0 : T75;
  assign T75 = T76 ? 1'h1 : R73;
  assign T76 = T65 & T77;
  assign T77 = T32[1'h1:1'h1];
  assign T79 = T72 ? 1'h0 : T80;
  assign T80 = T81 ? 1'h1 : R78;
  assign T81 = T65 & T82;
  assign T82 = T32[2'h2:2'h2];
  assign T83 = T84;
  assign T84 = {T173, T85};
  assign T85 = {T171, T86};
  assign T86 = T165 == pte_addr;
  assign pte_addr = T87 << 2'h3;
  assign T87 = T88;
  assign T88 = {r_pte_ppn, vpn_idx};
  assign vpn_idx = T100 ? T98 : T89;
  assign T89 = T96 ? T94 : T90;
  assign T90 = T91[4'h8:1'h0];
  assign T91 = r_req_addr >> 5'h12;
  assign T92 = T93 ? arb_io_out_bits_addr : r_req_addr;
  assign T93 = T0 & arb_io_out_valid;
  assign T94 = T95[4'h8:1'h0];
  assign T95 = r_req_addr >> 4'h9;
  assign T96 = T97[1'h0:1'h0];
  assign T97 = count;
  assign T98 = T99[4'h8:1'h0];
  assign T99 = r_req_addr >> 1'h0;
  assign T100 = T97[1'h1:1'h1];
  assign T101 = T15 ? pte_cache_data : T102;
  assign T102 = T106 ? T105 : T103;
  assign T103 = T93 ? T104 : r_pte_ppn;
  assign T104 = io_dpath_ptbr[5'h1f:4'hc];
  assign T105 = io_mem_resp_bits_data[5'h1d:4'ha];
  assign T106 = T148 & T107;
  assign T107 = set_dirty_bit ^ 1'h1;
  assign set_dirty_bit = perm_ok & T108;
  assign T108 = T113 | T109;
  assign T109 = r_req_store & T110;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_mem_resp_bits_data[3'h6:3'h6];
  assign T112 = T93 ? arb_io_out_bits_store : r_req_store;
  assign T113 = T114 ^ 1'h1;
  assign T114 = io_mem_resp_bits_data[3'h5:3'h5];
  assign perm_ok = T146 ? T134 : T115;
  assign T115 = r_req_fetch ? T127 : T116;
  assign T116 = r_req_store ? T121 : T117;
  assign T117 = T119 & T118;
  assign T118 = T70 < 4'h8;
  assign T119 = T71 & T120;
  assign T120 = 4'h2 <= T70;
  assign T121 = T123 & T122;
  assign T122 = T70[1'h0:1'h0];
  assign T123 = T125 & T124;
  assign T124 = T70 < 4'h8;
  assign T125 = T71 & T126;
  assign T126 = 4'h2 <= T70;
  assign T127 = T129 & T128;
  assign T128 = T70[1'h1:1'h1];
  assign T129 = T131 & T130;
  assign T130 = T70 < 4'h8;
  assign T131 = T71 & T132;
  assign T132 = 4'h2 <= T70;
  assign T133 = T93 ? arb_io_out_bits_fetch : r_req_fetch;
  assign T134 = r_req_fetch ? T142 : T135;
  assign T135 = r_req_store ? T138 : T136;
  assign T136 = T71 & T137;
  assign T137 = 4'h2 <= T70;
  assign T138 = T140 & T139;
  assign T139 = T70[1'h0:1'h0];
  assign T140 = T71 & T141;
  assign T141 = 4'h2 <= T70;
  assign T142 = T144 & T143;
  assign T143 = T70[1'h1:1'h1];
  assign T144 = T71 & T145;
  assign T145 = 4'h4 <= T70;
  assign T146 = r_req_prv[1'h0:1'h0];
  assign T147 = T93 ? arb_io_out_bits_prv : r_req_prv;
  assign T148 = io_mem_resp_valid & T149;
  assign T149 = state == 3'h2;
  assign pte_cache_data = T158 | T150;
  assign T150 = T157 ? T151 : 20'h0;
  assign T151 = T152[2'h2];
  assign T154 = T65 & T155;
  assign T155 = T156 < 2'h3;
  assign T156 = T34[1'h1:1'h0];
  assign T157 = T23[2'h2:2'h2];
  assign T158 = T162 | T159;
  assign T159 = T161 ? T160 : 20'h0;
  assign T160 = T152[2'h1];
  assign T161 = T23[1'h1:1'h1];
  assign T162 = T164 ? T163 : 20'h0;
  assign T163 = T152[2'h0];
  assign T164 = T23[1'h0:1'h0];
  assign T165 = T166[2'h0];
  assign T168 = T65 & T169;
  assign T169 = T170 < 2'h3;
  assign T170 = T34[1'h1:1'h0];
  assign T171 = T172 == pte_addr;
  assign T172 = T166[2'h1];
  assign T173 = T174 == pte_addr;
  assign T174 = T166[2'h2];
  assign T175 = 3'h1 == state;
  assign T176 = T175 & T177;
  assign T177 = T178 & io_mem_req_ready;
  assign T178 = T16 ^ 1'h1;
  assign T179 = T180 & io_mem_resp_bits_nack;
  assign T180 = 3'h2 == state;
  assign T181 = T180 & io_mem_resp_valid;
  assign T182 = T181 & T183;
  assign T183 = T185 & T184;
  assign T184 = count < 2'h2;
  assign T185 = T71 & T186;
  assign T186 = T70 < 4'h2;
  assign T187 = set_dirty_bit ? 3'h3 : 3'h5;
  assign T188 = T181 & T189;
  assign T189 = T71 & T190;
  assign T190 = 4'h2 <= T70;
  assign T191 = T192 & io_mem_req_ready;
  assign T192 = 3'h3 == state;
  assign T193 = T194 & io_mem_resp_bits_nack;
  assign T194 = 3'h4 == state;
  assign T195 = T194 & io_mem_resp_valid;
  assign T196 = 3'h5 == state;
  assign T197 = 3'h6 == state;
  assign io_mem_req_bits_data = T243;
  assign T243 = {34'h0, T198};
  assign T198 = T199;
  assign T199 = {T202, T200};
  assign T200 = {pte_wdata_r, T201};
  assign T201 = {pte_wdata_typ, pte_wdata_v};
  assign pte_wdata_v = 1'h0;
  assign pte_wdata_typ = 4'h0;
  assign pte_wdata_r = 1'h1;
  assign T202 = {pte_wdata_ppn, T203};
  assign T203 = {pte_wdata_reserved_for_software, pte_wdata_d};
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_reserved_for_software = 3'h0;
  assign pte_wdata_ppn = 20'h0;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_cmd = T204;
  assign T204 = T205 ? 5'ha : 5'h0;
  assign T205 = state == 3'h3;
  assign io_mem_req_bits_addr = T244;
  assign T244 = {8'h0, pte_addr};
  assign io_mem_req_valid = T206;
  assign T206 = T15 ? 1'h0 : T207;
  assign T207 = T209 | T208;
  assign T208 = state == 3'h3;
  assign T209 = state == 3'h1;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_ie = io_dpath_status_ie;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_0_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_0_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_0_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_0_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_0_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign T210 = T106 ? T71 : r_pte_v;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign T211 = T106 ? T70 : r_pte_typ;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign T212 = T106 ? T114 : r_pte_r;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign T213 = T106 ? T111 : r_pte_d;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign T214 = T106 ? T215 : r_pte_reserved_for_software;
  assign T215 = io_mem_resp_bits_data[4'h9:3'h7];
  assign io_requestor_0_resp_bits_pte_ppn = T245;
  assign T245 = resp_ppn[5'h13:1'h0];
  assign resp_ppn = T225 ? r_resp_ppn : T216;
  assign T216 = T223 ? T220 : T217;
  assign T217 = {T219, T218};
  assign T218 = r_req_addr[5'h11:1'h0];
  assign T219 = r_resp_ppn >> 5'h12;
  assign T220 = {T222, T221};
  assign T221 = r_req_addr[4'h8:1'h0];
  assign T222 = r_resp_ppn >> 4'h9;
  assign T223 = T224[1'h0:1'h0];
  assign T224 = count;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hc;
  assign T225 = T224[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = state == 3'h6;
  assign io_requestor_0_resp_valid = T226;
  assign T226 = resp_val & T227;
  assign T227 = r_req_dest == 1'h0;
  assign T228 = T93 ? arb_io_chosen : r_req_dest;
  assign resp_val = T229 | resp_err;
  assign T229 = state == 3'h5;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_ie = io_dpath_status_ie;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_ie1 = io_dpath_status_ie1;
  assign io_requestor_1_status_prv1 = io_dpath_status_prv1;
  assign io_requestor_1_status_ie2 = io_dpath_status_ie2;
  assign io_requestor_1_status_prv2 = io_dpath_status_prv2;
  assign io_requestor_1_status_ie3 = io_dpath_status_ie3;
  assign io_requestor_1_status_prv3 = io_dpath_status_prv3;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_ppn = T246;
  assign T246 = resp_ppn[5'h13:1'h0];
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T230;
  assign T230 = resp_val & T231;
  assign T231 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_2 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits_addr( io_requestor_1_req_bits_addr ),
       .io_in_1_bits_prv( io_requestor_1_req_bits_prv ),
       .io_in_1_bits_store( io_requestor_1_req_bits_store ),
       .io_in_1_bits_fetch( io_requestor_1_req_bits_fetch ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits_addr( io_requestor_0_req_bits_addr ),
       .io_in_0_bits_prv( io_requestor_0_req_bits_prv ),
       .io_in_0_bits_store( io_requestor_0_req_bits_store ),
       .io_in_0_bits_fetch( io_requestor_0_req_bits_fetch ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits_addr( arb_io_out_bits_addr ),
       .io_out_bits_prv( arb_io_out_bits_prv ),
       .io_out_bits_store( arb_io_out_bits_store ),
       .io_out_bits_fetch( arb_io_out_bits_fetch ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T197) begin
      state <= 3'h0;
    end else if(T196) begin
      state <= 3'h0;
    end else if(T195) begin
      state <= 3'h1;
    end else if(T193) begin
      state <= 3'h3;
    end else if(T191) begin
      state <= 3'h4;
    end else if(T188) begin
      state <= T187;
    end else if(T182) begin
      state <= 3'h1;
    end else if(T181) begin
      state <= 3'h6;
    end else if(T179) begin
      state <= 3'h1;
    end else if(T176) begin
      state <= 3'h2;
    end else if(T15) begin
      state <= 3'h1;
    end else if(T13) begin
      state <= 3'h1;
    end
    if(T182) begin
      count <= T22;
    end else if(T15) begin
      count <= T21;
    end else if(T14) begin
      count <= 2'h0;
    end
    if(T72) begin
      R27 <= 1'h0;
    end else if(T30) begin
      R27 <= 1'h1;
    end
    if(T60) begin
      R45 <= T47;
    end
    if(T72) begin
      R73 <= 1'h0;
    end else if(T76) begin
      R73 <= 1'h1;
    end
    if(T72) begin
      R78 <= 1'h0;
    end else if(T81) begin
      R78 <= 1'h1;
    end
    if(T93) begin
      r_req_addr <= arb_io_out_bits_addr;
    end
    if(T15) begin
      r_pte_ppn <= pte_cache_data;
    end else if(T106) begin
      r_pte_ppn <= T105;
    end else if(T93) begin
      r_pte_ppn <= T104;
    end
    if(T93) begin
      r_req_store <= arb_io_out_bits_store;
    end
    if(T93) begin
      r_req_fetch <= arb_io_out_bits_fetch;
    end
    if(T93) begin
      r_req_prv <= arb_io_out_bits_prv;
    end
    if (T154)
      T152[T34] <= T105;
    if (T168)
      T166[T34] <= pte_addr;
    if(T106) begin
      r_pte_v <= T71;
    end
    if(T106) begin
      r_pte_typ <= T70;
    end
    if(T106) begin
      r_pte_r <= T114;
    end
    if(T106) begin
      r_pte_d <= T111;
    end
    if(T106) begin
      r_pte_reserved_for_software <= T215;
    end
    if(T93) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [39:0] io_requestor_1_req_bits_addr,
    input [8:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_kill,
    input  io_requestor_1_req_bits_phys,
    input [63:0] io_requestor_1_req_bits_data,
    output io_requestor_1_resp_valid,
    output[39:0] io_requestor_1_resp_bits_addr,
    output[8:0] io_requestor_1_resp_bits_tag,
    output[4:0] io_requestor_1_resp_bits_cmd,
    output[2:0] io_requestor_1_resp_bits_typ,
    output[63:0] io_requestor_1_resp_bits_data,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data_word_bypass,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[8:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    input  io_requestor_1_invalidate_lr,
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [39:0] io_requestor_0_req_bits_addr,
    input [8:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_kill,
    input  io_requestor_0_req_bits_phys,
    input [63:0] io_requestor_0_req_bits_data,
    output io_requestor_0_resp_valid,
    output[39:0] io_requestor_0_resp_bits_addr,
    output[8:0] io_requestor_0_resp_bits_tag,
    output[4:0] io_requestor_0_resp_bits_cmd,
    output[2:0] io_requestor_0_resp_bits_typ,
    output[63:0] io_requestor_0_resp_bits_data,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data_word_bypass,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[8:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_invalidate_lr
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[39:0] io_mem_req_bits_addr,
    output[8:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_kill,
    output io_mem_req_bits_phys,
    output[63:0] io_mem_req_bits_data,
    input  io_mem_resp_valid,
    input [39:0] io_mem_resp_bits_addr,
    input [8:0] io_mem_resp_bits_tag,
    input [4:0] io_mem_resp_bits_cmd,
    input [2:0] io_mem_resp_bits_typ,
    input [63:0] io_mem_resp_bits_data,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data_word_bypass,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [8:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_invalidate_lr
    input  io_mem_ordered
);

  wire[63:0] T0;
  reg  r_valid_0;
  wire T1;
  wire T2;
  wire[2:0] T3;
  wire[4:0] T4;
  wire[8:0] T32;
  wire[9:0] T5;
  wire[9:0] T6;
  wire[9:0] T7;
  wire[39:0] T8;
  wire T9;
  wire[8:0] T33;
  wire[7:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[8:0] T34;
  wire[7:0] T18;
  wire T19;
  wire[8:0] T35;
  wire[7:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[8:0] T36;
  wire[7:0] T28;
  wire T29;
  wire T30;
  wire T31;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_invalidate_lr = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_req_bits_data = T0;
  assign T0 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_phys = T1;
  assign T1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_kill = T2;
  assign T2 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_bits_typ = T3;
  assign T3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_cmd = T4;
  assign T4 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T32;
  assign T32 = T5[4'h8:1'h0];
  assign T5 = io_requestor_0_req_valid ? T7 : T6;
  assign T6 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T7 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_addr = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_valid = T9;
  assign T9 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T33;
  assign T33 = {1'h0, T10};
  assign T10 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T11;
  assign T11 = io_mem_replay_next_valid & T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_replay = T14;
  assign T14 = io_mem_resp_bits_replay & T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T17;
  assign T17 = io_mem_resp_bits_nack & T15;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T34;
  assign T34 = {1'h0, T18};
  assign T18 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_valid = T19;
  assign T19 = io_mem_resp_valid & T15;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T35;
  assign T35 = {1'h0, T20};
  assign T20 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T21;
  assign T21 = io_mem_replay_next_valid & T22;
  assign T22 = T23 == 1'h1;
  assign T23 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_replay = T24;
  assign T24 = io_mem_resp_bits_replay & T25;
  assign T25 = T26 == 1'h1;
  assign T26 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T27;
  assign T27 = io_mem_resp_bits_nack & T25;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T36;
  assign T36 = {1'h0, T28};
  assign T28 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_valid = T29;
  assign T29 = io_mem_resp_valid & T25;
  assign io_requestor_1_req_ready = T30;
  assign T30 = io_requestor_0_req_ready & T31;
  assign T31 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RocketTile(input clk, input reset,
    input  io_cached_0_acquire_ready,
    output io_cached_0_acquire_valid,
    output[25:0] io_cached_0_acquire_bits_addr_block,
    output[1:0] io_cached_0_acquire_bits_client_xact_id,
    output[1:0] io_cached_0_acquire_bits_addr_beat,
    output io_cached_0_acquire_bits_is_builtin_type,
    output[2:0] io_cached_0_acquire_bits_a_type,
    output[16:0] io_cached_0_acquire_bits_union,
    output[127:0] io_cached_0_acquire_bits_data,
    output io_cached_0_grant_ready,
    input  io_cached_0_grant_valid,
    input [1:0] io_cached_0_grant_bits_addr_beat,
    input [1:0] io_cached_0_grant_bits_client_xact_id,
    input [2:0] io_cached_0_grant_bits_manager_xact_id,
    input  io_cached_0_grant_bits_is_builtin_type,
    input [3:0] io_cached_0_grant_bits_g_type,
    input [127:0] io_cached_0_grant_bits_data,
    output io_cached_0_probe_ready,
    input  io_cached_0_probe_valid,
    input [25:0] io_cached_0_probe_bits_addr_block,
    input [1:0] io_cached_0_probe_bits_p_type,
    input  io_cached_0_release_ready,
    output io_cached_0_release_valid,
    output[1:0] io_cached_0_release_bits_addr_beat,
    output[25:0] io_cached_0_release_bits_addr_block,
    output[1:0] io_cached_0_release_bits_client_xact_id,
    output io_cached_0_release_bits_voluntary,
    output[2:0] io_cached_0_release_bits_r_type,
    output[127:0] io_cached_0_release_bits_data,
    input  io_uncached_0_acquire_ready,
    output io_uncached_0_acquire_valid,
    output[25:0] io_uncached_0_acquire_bits_addr_block,
    output[1:0] io_uncached_0_acquire_bits_client_xact_id,
    output[1:0] io_uncached_0_acquire_bits_addr_beat,
    output io_uncached_0_acquire_bits_is_builtin_type,
    output[2:0] io_uncached_0_acquire_bits_a_type,
    output[16:0] io_uncached_0_acquire_bits_union,
    output[127:0] io_uncached_0_acquire_bits_data,
    output io_uncached_0_grant_ready,
    input  io_uncached_0_grant_valid,
    input [1:0] io_uncached_0_grant_bits_addr_beat,
    input [1:0] io_uncached_0_grant_bits_client_xact_id,
    input [2:0] io_uncached_0_grant_bits_manager_xact_id,
    input  io_uncached_0_grant_bits_is_builtin_type,
    input [3:0] io_uncached_0_grant_bits_g_type,
    input [127:0] io_uncached_0_grant_bits_data,
    input  io_host_reset,
    input  io_host_id,
    output io_host_csr_req_ready,
    input  io_host_csr_req_valid,
    input  io_host_csr_req_bits_rw,
    input [11:0] io_host_csr_req_bits_addr,
    input [63:0] io_host_csr_req_bits_data,
    input  io_host_csr_resp_ready,
    output io_host_csr_resp_valid,
    output[63:0] io_host_csr_resp_bits,
    output io_host_debug_stats_csr,
    //input  io_dma_req_ready
    output io_dma_req_valid,
    //output[1:0] io_dma_req_bits_client_xact_id
    //output[1:0] io_dma_req_bits_cmd
    //output[31:0] io_dma_req_bits_source
    //output[31:0] io_dma_req_bits_dest
    //output[31:0] io_dma_req_bits_length
    output io_dma_resp_ready
    //input  io_dma_resp_valid
    //input [1:0] io_dma_resp_bits_client_xact_id
    //input [1:0] io_dma_resp_bits_status
);

  wire dcArb_io_requestor_1_req_ready;
  wire dcArb_io_requestor_1_resp_valid;
  wire[39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[8:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[8:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_0_req_ready;
  wire dcArb_io_requestor_0_resp_valid;
  wire[39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[8:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_mem_req_valid;
  wire[39:0] dcArb_io_mem_req_bits_addr;
  wire[8:0] dcArb_io_mem_req_bits_tag;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_kill;
  wire dcArb_io_mem_req_bits_phys;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire core_io_host_csr_req_ready;
  wire core_io_host_csr_resp_valid;
  wire[63:0] core_io_host_csr_resp_bits;
  wire core_io_host_debug_stats_csr;
  wire core_io_imem_req_valid;
  wire[39:0] core_io_imem_req_bits_pc;
  wire core_io_imem_resp_ready;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_bits_mask;
  wire core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_btb_update_bits_pc;
  wire[38:0] core_io_imem_btb_update_bits_target;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_isReturn;
  wire[38:0] core_io_imem_btb_update_bits_br_pc;
  wire core_io_imem_bht_update_valid;
  wire core_io_imem_bht_update_bits_prediction_valid;
  wire core_io_imem_bht_update_bits_prediction_bits_taken;
  wire core_io_imem_bht_update_bits_prediction_bits_mask;
  wire core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire[38:0] core_io_imem_bht_update_bits_pc;
  wire core_io_imem_bht_update_bits_taken;
  wire core_io_imem_bht_update_bits_mispredict;
  wire core_io_imem_ras_update_valid;
  wire core_io_imem_ras_update_bits_isCall;
  wire core_io_imem_ras_update_bits_isReturn;
  wire[38:0] core_io_imem_ras_update_bits_returnAddr;
  wire core_io_imem_ras_update_bits_prediction_valid;
  wire core_io_imem_ras_update_bits_prediction_bits_taken;
  wire core_io_imem_ras_update_bits_prediction_bits_mask;
  wire core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire[38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire[2:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire[3:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire[1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire core_io_imem_invalidate;
  wire core_io_dmem_req_valid;
  wire[39:0] core_io_dmem_req_bits_addr;
  wire[8:0] core_io_dmem_req_bits_tag;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_bits_phys;
  wire[63:0] core_io_dmem_req_bits_data;
  wire core_io_dmem_invalidate_lr;
  wire[31:0] core_io_ptw_ptbr;
  wire core_io_ptw_invalidate;
  wire core_io_ptw_status_sd;
  wire[30:0] core_io_ptw_status_zero2;
  wire core_io_ptw_status_sd_rv32;
  wire[8:0] core_io_ptw_status_zero1;
  wire[4:0] core_io_ptw_status_vm;
  wire core_io_ptw_status_mprv;
  wire[1:0] core_io_ptw_status_xs;
  wire[1:0] core_io_ptw_status_fs;
  wire[1:0] core_io_ptw_status_prv3;
  wire core_io_ptw_status_ie3;
  wire[1:0] core_io_ptw_status_prv2;
  wire core_io_ptw_status_ie2;
  wire[1:0] core_io_ptw_status_prv1;
  wire core_io_ptw_status_ie1;
  wire[1:0] core_io_ptw_status_prv;
  wire core_io_ptw_status_ie;
  wire ptw_io_requestor_1_req_ready;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_resp_bits_error;
  wire[19:0] ptw_io_requestor_1_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_1_resp_bits_pte_d;
  wire ptw_io_requestor_1_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_1_resp_bits_pte_typ;
  wire ptw_io_requestor_1_resp_bits_pte_v;
  wire ptw_io_requestor_1_status_sd;
  wire[30:0] ptw_io_requestor_1_status_zero2;
  wire ptw_io_requestor_1_status_sd_rv32;
  wire[8:0] ptw_io_requestor_1_status_zero1;
  wire[4:0] ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_mprv;
  wire[1:0] ptw_io_requestor_1_status_xs;
  wire[1:0] ptw_io_requestor_1_status_fs;
  wire[1:0] ptw_io_requestor_1_status_prv3;
  wire ptw_io_requestor_1_status_ie3;
  wire[1:0] ptw_io_requestor_1_status_prv2;
  wire ptw_io_requestor_1_status_ie2;
  wire[1:0] ptw_io_requestor_1_status_prv1;
  wire ptw_io_requestor_1_status_ie1;
  wire[1:0] ptw_io_requestor_1_status_prv;
  wire ptw_io_requestor_1_status_ie;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_0_req_ready;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_resp_bits_error;
  wire[19:0] ptw_io_requestor_0_resp_bits_pte_ppn;
  wire[2:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire ptw_io_requestor_0_resp_bits_pte_d;
  wire ptw_io_requestor_0_resp_bits_pte_r;
  wire[3:0] ptw_io_requestor_0_resp_bits_pte_typ;
  wire ptw_io_requestor_0_resp_bits_pte_v;
  wire ptw_io_requestor_0_status_sd;
  wire[30:0] ptw_io_requestor_0_status_zero2;
  wire ptw_io_requestor_0_status_sd_rv32;
  wire[8:0] ptw_io_requestor_0_status_zero1;
  wire[4:0] ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_mprv;
  wire[1:0] ptw_io_requestor_0_status_xs;
  wire[1:0] ptw_io_requestor_0_status_fs;
  wire[1:0] ptw_io_requestor_0_status_prv3;
  wire ptw_io_requestor_0_status_ie3;
  wire[1:0] ptw_io_requestor_0_status_prv2;
  wire ptw_io_requestor_0_status_ie2;
  wire[1:0] ptw_io_requestor_0_status_prv1;
  wire ptw_io_requestor_0_status_ie1;
  wire[1:0] ptw_io_requestor_0_status_prv;
  wire ptw_io_requestor_0_status_ie;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_mem_req_valid;
  wire[39:0] ptw_io_mem_req_bits_addr;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_bits_phys;
  wire[63:0] ptw_io_mem_req_bits_data;
  wire icache_io_cpu_resp_valid;
  wire[39:0] icache_io_cpu_resp_bits_pc;
  wire[31:0] icache_io_cpu_resp_bits_data_0;
  wire icache_io_cpu_resp_bits_mask;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_bits_mask;
  wire icache_io_cpu_btb_resp_bits_bridx;
  wire[38:0] icache_io_cpu_btb_resp_bits_target;
  wire[2:0] icache_io_cpu_btb_resp_bits_entry;
  wire[3:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[39:0] icache_io_cpu_npc;
  wire icache_io_ptw_req_valid;
  wire[26:0] icache_io_ptw_req_bits_addr;
  wire[1:0] icache_io_ptw_req_bits_prv;
  wire icache_io_ptw_req_bits_store;
  wire icache_io_ptw_req_bits_fetch;
  wire icache_io_mem_acquire_valid;
  wire[25:0] icache_io_mem_acquire_bits_addr_block;
  wire[1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] icache_io_mem_acquire_bits_addr_beat;
  wire icache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] icache_io_mem_acquire_bits_a_type;
  wire[16:0] icache_io_mem_acquire_bits_union;
  wire[127:0] icache_io_mem_acquire_bits_data;
  wire icache_io_mem_grant_ready;
  wire dcache_io_cpu_req_ready;
  wire dcache_io_cpu_resp_valid;
  wire[39:0] dcache_io_cpu_resp_bits_addr;
  wire[8:0] dcache_io_cpu_resp_bits_tag;
  wire[4:0] dcache_io_cpu_resp_bits_cmd;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[63:0] dcache_io_cpu_resp_bits_data_word_bypass;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire dcache_io_cpu_replay_next_valid;
  wire[8:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_ordered;
  wire dcache_io_ptw_req_valid;
  wire[26:0] dcache_io_ptw_req_bits_addr;
  wire[1:0] dcache_io_ptw_req_bits_prv;
  wire dcache_io_ptw_req_bits_store;
  wire dcache_io_ptw_req_bits_fetch;
  wire dcache_io_mem_acquire_valid;
  wire[25:0] dcache_io_mem_acquire_bits_addr_block;
  wire[1:0] dcache_io_mem_acquire_bits_client_xact_id;
  wire[1:0] dcache_io_mem_acquire_bits_addr_beat;
  wire dcache_io_mem_acquire_bits_is_builtin_type;
  wire[2:0] dcache_io_mem_acquire_bits_a_type;
  wire[16:0] dcache_io_mem_acquire_bits_union;
  wire[127:0] dcache_io_mem_acquire_bits_data;
  wire dcache_io_mem_grant_ready;
  wire dcache_io_mem_probe_ready;
  wire dcache_io_mem_release_valid;
  wire[1:0] dcache_io_mem_release_bits_addr_beat;
  wire[25:0] dcache_io_mem_release_bits_addr_block;
  wire[1:0] dcache_io_mem_release_bits_client_xact_id;
  wire dcache_io_mem_release_bits_voluntary;
  wire[2:0] dcache_io_mem_release_bits_r_type;
  wire[127:0] dcache_io_mem_release_bits_data;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_dma_req_bits_length = {1{$random}};
//  assign io_dma_req_bits_dest = {1{$random}};
//  assign io_dma_req_bits_source = {1{$random}};
//  assign io_dma_req_bits_cmd = {1{$random}};
//  assign io_dma_req_bits_client_xact_id = {1{$random}};
// synthesis translate_on
`endif
  assign io_dma_resp_ready = 1'h0;
  assign io_dma_req_valid = 1'h0;
  assign io_host_debug_stats_csr = core_io_host_debug_stats_csr;
  assign io_host_csr_resp_bits = core_io_host_csr_resp_bits;
  assign io_host_csr_resp_valid = core_io_host_csr_resp_valid;
  assign io_host_csr_req_ready = core_io_host_csr_req_ready;
  assign io_uncached_0_grant_ready = icache_io_mem_grant_ready;
  assign io_uncached_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_uncached_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_uncached_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_uncached_0_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cached_0_release_bits_data = dcache_io_mem_release_bits_data;
  assign io_cached_0_release_bits_r_type = dcache_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_voluntary = dcache_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_client_xact_id = dcache_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_addr_block = dcache_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_addr_beat = dcache_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_valid = dcache_io_mem_release_valid;
  assign io_cached_0_probe_ready = dcache_io_mem_probe_ready;
  assign io_cached_0_grant_ready = dcache_io_mem_grant_ready;
  assign io_cached_0_acquire_bits_data = dcache_io_mem_acquire_bits_data;
  assign io_cached_0_acquire_bits_union = dcache_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_a_type = dcache_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_is_builtin_type = dcache_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_addr_beat = dcache_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_client_xact_id = dcache_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_block = dcache_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_valid = dcache_io_mem_acquire_valid;
  Rocket core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_csr_req_ready( core_io_host_csr_req_ready ),
       .io_host_csr_req_valid( io_host_csr_req_valid ),
       .io_host_csr_req_bits_rw( io_host_csr_req_bits_rw ),
       .io_host_csr_req_bits_addr( io_host_csr_req_bits_addr ),
       .io_host_csr_req_bits_data( io_host_csr_req_bits_data ),
       .io_host_csr_resp_ready( io_host_csr_resp_ready ),
       .io_host_csr_resp_valid( core_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( core_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( core_io_host_debug_stats_csr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_imem_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_imem_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_imem_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_imem_btb_update_bits_taken(  )
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_imem_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_imem_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_imem_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_imem_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_imem_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_imem_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_imem_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_imem_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_imem_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_imem_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_imem_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_imem_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_imem_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_imem_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_imem_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_imem_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_imem_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_imem_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_imem_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_imem_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_imem_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_imem_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_imem_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_imem_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_imem_npc( icache_io_cpu_npc ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_dmem_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_status_sd( core_io_ptw_status_sd ),
       .io_ptw_status_zero2( core_io_ptw_status_zero2 ),
       .io_ptw_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_ptw_status_zero1( core_io_ptw_status_zero1 ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_mprv( core_io_ptw_status_mprv ),
       .io_ptw_status_xs( core_io_ptw_status_xs ),
       .io_ptw_status_fs( core_io_ptw_status_fs ),
       .io_ptw_status_prv3( core_io_ptw_status_prv3 ),
       .io_ptw_status_ie3( core_io_ptw_status_ie3 ),
       .io_ptw_status_prv2( core_io_ptw_status_prv2 ),
       .io_ptw_status_ie2( core_io_ptw_status_ie2 ),
       .io_ptw_status_prv1( core_io_ptw_status_prv1 ),
       .io_ptw_status_ie1( core_io_ptw_status_ie1 ),
       .io_ptw_status_prv( core_io_ptw_status_prv ),
       .io_ptw_status_ie( core_io_ptw_status_ie )
       //.io_fpu_inst(  )
       //.io_fpu_fromint_data(  )
       //.io_fpu_fcsr_rm(  )
       //.io_fpu_fcsr_flags_valid(  )
       //.io_fpu_fcsr_flags_bits(  )
       //.io_fpu_store_data(  )
       //.io_fpu_toint_data(  )
       //.io_fpu_dmem_resp_val(  )
       //.io_fpu_dmem_resp_type(  )
       //.io_fpu_dmem_resp_tag(  )
       //.io_fpu_dmem_resp_data(  )
       //.io_fpu_valid(  )
       //.io_fpu_fcsr_rdy(  )
       //.io_fpu_nack_mem(  )
       //.io_fpu_illegal_rm(  )
       //.io_fpu_killx(  )
       //.io_fpu_killm(  )
       //.io_fpu_dec_cmd(  )
       //.io_fpu_dec_ldst(  )
       //.io_fpu_dec_wen(  )
       //.io_fpu_dec_ren1(  )
       //.io_fpu_dec_ren2(  )
       //.io_fpu_dec_ren3(  )
       //.io_fpu_dec_swap12(  )
       //.io_fpu_dec_swap23(  )
       //.io_fpu_dec_single(  )
       //.io_fpu_dec_fromint(  )
       //.io_fpu_dec_toint(  )
       //.io_fpu_dec_fastpipe(  )
       //.io_fpu_dec_fma(  )
       //.io_fpu_dec_div(  )
       //.io_fpu_dec_sqrt(  )
       //.io_fpu_dec_round(  )
       //.io_fpu_dec_wflags(  )
       //.io_fpu_sboard_set(  )
       //.io_fpu_sboard_clr(  )
       //.io_fpu_sboard_clra(  )
       //.io_fpu_cp_req_ready(  )
       //.io_fpu_cp_req_valid(  )
       //.io_fpu_cp_req_bits_cmd(  )
       //.io_fpu_cp_req_bits_ldst(  )
       //.io_fpu_cp_req_bits_wen(  )
       //.io_fpu_cp_req_bits_ren1(  )
       //.io_fpu_cp_req_bits_ren2(  )
       //.io_fpu_cp_req_bits_ren3(  )
       //.io_fpu_cp_req_bits_swap12(  )
       //.io_fpu_cp_req_bits_swap23(  )
       //.io_fpu_cp_req_bits_single(  )
       //.io_fpu_cp_req_bits_fromint(  )
       //.io_fpu_cp_req_bits_toint(  )
       //.io_fpu_cp_req_bits_fastpipe(  )
       //.io_fpu_cp_req_bits_fma(  )
       //.io_fpu_cp_req_bits_div(  )
       //.io_fpu_cp_req_bits_sqrt(  )
       //.io_fpu_cp_req_bits_round(  )
       //.io_fpu_cp_req_bits_wflags(  )
       //.io_fpu_cp_req_bits_rm(  )
       //.io_fpu_cp_req_bits_typ(  )
       //.io_fpu_cp_req_bits_in1(  )
       //.io_fpu_cp_req_bits_in2(  )
       //.io_fpu_cp_req_bits_in3(  )
       //.io_fpu_cp_resp_ready(  )
       //.io_fpu_cp_resp_valid(  )
       //.io_fpu_cp_resp_bits_data(  )
       //.io_fpu_cp_resp_bits_exc(  )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data_word_bypass(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_invalidate_lr(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_autl_acquire_ready(  )
       //.io_rocc_autl_acquire_valid(  )
       //.io_rocc_autl_acquire_bits_addr_block(  )
       //.io_rocc_autl_acquire_bits_client_xact_id(  )
       //.io_rocc_autl_acquire_bits_addr_beat(  )
       //.io_rocc_autl_acquire_bits_is_builtin_type(  )
       //.io_rocc_autl_acquire_bits_a_type(  )
       //.io_rocc_autl_acquire_bits_union(  )
       //.io_rocc_autl_acquire_bits_data(  )
       //.io_rocc_autl_grant_ready(  )
       //.io_rocc_autl_grant_valid(  )
       //.io_rocc_autl_grant_bits_addr_beat(  )
       //.io_rocc_autl_grant_bits_client_xact_id(  )
       //.io_rocc_autl_grant_bits_manager_xact_id(  )
       //.io_rocc_autl_grant_bits_is_builtin_type(  )
       //.io_rocc_autl_grant_bits_g_type(  )
       //.io_rocc_autl_grant_bits_data(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits_addr(  )
       //.io_rocc_iptw_req_bits_prv(  )
       //.io_rocc_iptw_req_bits_store(  )
       //.io_rocc_iptw_req_bits_fetch(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_pte_ppn(  )
       //.io_rocc_iptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_iptw_resp_bits_pte_d(  )
       //.io_rocc_iptw_resp_bits_pte_r(  )
       //.io_rocc_iptw_resp_bits_pte_typ(  )
       //.io_rocc_iptw_resp_bits_pte_v(  )
       //.io_rocc_iptw_status_sd(  )
       //.io_rocc_iptw_status_zero2(  )
       //.io_rocc_iptw_status_sd_rv32(  )
       //.io_rocc_iptw_status_zero1(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_mprv(  )
       //.io_rocc_iptw_status_xs(  )
       //.io_rocc_iptw_status_fs(  )
       //.io_rocc_iptw_status_prv3(  )
       //.io_rocc_iptw_status_ie3(  )
       //.io_rocc_iptw_status_prv2(  )
       //.io_rocc_iptw_status_ie2(  )
       //.io_rocc_iptw_status_prv1(  )
       //.io_rocc_iptw_status_ie1(  )
       //.io_rocc_iptw_status_prv(  )
       //.io_rocc_iptw_status_ie(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits_addr(  )
       //.io_rocc_dptw_req_bits_prv(  )
       //.io_rocc_dptw_req_bits_store(  )
       //.io_rocc_dptw_req_bits_fetch(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_pte_ppn(  )
       //.io_rocc_dptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_dptw_resp_bits_pte_d(  )
       //.io_rocc_dptw_resp_bits_pte_r(  )
       //.io_rocc_dptw_resp_bits_pte_typ(  )
       //.io_rocc_dptw_resp_bits_pte_v(  )
       //.io_rocc_dptw_status_sd(  )
       //.io_rocc_dptw_status_zero2(  )
       //.io_rocc_dptw_status_sd_rv32(  )
       //.io_rocc_dptw_status_zero1(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_mprv(  )
       //.io_rocc_dptw_status_xs(  )
       //.io_rocc_dptw_status_fs(  )
       //.io_rocc_dptw_status_prv3(  )
       //.io_rocc_dptw_status_ie3(  )
       //.io_rocc_dptw_status_prv2(  )
       //.io_rocc_dptw_status_ie2(  )
       //.io_rocc_dptw_status_prv1(  )
       //.io_rocc_dptw_status_ie1(  )
       //.io_rocc_dptw_status_prv(  )
       //.io_rocc_dptw_status_ie(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits_addr(  )
       //.io_rocc_pptw_req_bits_prv(  )
       //.io_rocc_pptw_req_bits_store(  )
       //.io_rocc_pptw_req_bits_fetch(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_pte_ppn(  )
       //.io_rocc_pptw_resp_bits_pte_reserved_for_software(  )
       //.io_rocc_pptw_resp_bits_pte_d(  )
       //.io_rocc_pptw_resp_bits_pte_r(  )
       //.io_rocc_pptw_resp_bits_pte_typ(  )
       //.io_rocc_pptw_resp_bits_pte_v(  )
       //.io_rocc_pptw_status_sd(  )
       //.io_rocc_pptw_status_zero2(  )
       //.io_rocc_pptw_status_sd_rv32(  )
       //.io_rocc_pptw_status_zero1(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_mprv(  )
       //.io_rocc_pptw_status_xs(  )
       //.io_rocc_pptw_status_fs(  )
       //.io_rocc_pptw_status_prv3(  )
       //.io_rocc_pptw_status_ie3(  )
       //.io_rocc_pptw_status_prv2(  )
       //.io_rocc_pptw_status_ie2(  )
       //.io_rocc_pptw_status_prv1(  )
       //.io_rocc_pptw_status_ie1(  )
       //.io_rocc_pptw_status_prv(  )
       //.io_rocc_pptw_status_ie(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_fpu_req_ready(  )
       //.io_rocc_fpu_req_valid(  )
       //.io_rocc_fpu_req_bits_cmd(  )
       //.io_rocc_fpu_req_bits_ldst(  )
       //.io_rocc_fpu_req_bits_wen(  )
       //.io_rocc_fpu_req_bits_ren1(  )
       //.io_rocc_fpu_req_bits_ren2(  )
       //.io_rocc_fpu_req_bits_ren3(  )
       //.io_rocc_fpu_req_bits_swap12(  )
       //.io_rocc_fpu_req_bits_swap23(  )
       //.io_rocc_fpu_req_bits_single(  )
       //.io_rocc_fpu_req_bits_fromint(  )
       //.io_rocc_fpu_req_bits_toint(  )
       //.io_rocc_fpu_req_bits_fastpipe(  )
       //.io_rocc_fpu_req_bits_fma(  )
       //.io_rocc_fpu_req_bits_div(  )
       //.io_rocc_fpu_req_bits_sqrt(  )
       //.io_rocc_fpu_req_bits_round(  )
       //.io_rocc_fpu_req_bits_wflags(  )
       //.io_rocc_fpu_req_bits_rm(  )
       //.io_rocc_fpu_req_bits_typ(  )
       //.io_rocc_fpu_req_bits_in1(  )
       //.io_rocc_fpu_req_bits_in2(  )
       //.io_rocc_fpu_req_bits_in3(  )
       //.io_rocc_fpu_resp_ready(  )
       //.io_rocc_fpu_resp_valid(  )
       //.io_rocc_fpu_resp_bits_data(  )
       //.io_rocc_fpu_resp_bits_exc(  )
       //.io_rocc_exception(  )
       //.io_rocc_dma_req_ready(  )
       //.io_rocc_dma_req_valid(  )
       //.io_rocc_dma_req_bits_client_xact_id(  )
       //.io_rocc_dma_req_bits_cmd(  )
       //.io_rocc_dma_req_bits_source(  )
       //.io_rocc_dma_req_bits_dest(  )
       //.io_rocc_dma_req_bits_length(  )
       //.io_rocc_dma_resp_ready(  )
       //.io_rocc_dma_resp_valid(  )
       //.io_rocc_dma_resp_bits_client_xact_id(  )
       //.io_rocc_dma_resp_bits_status(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign core.io_fpu_fcsr_flags_valid = {1{$random}};
    assign core.io_fpu_fcsr_flags_bits = {1{$random}};
    assign core.io_fpu_store_data = {2{$random}};
    assign core.io_fpu_toint_data = {2{$random}};
    assign core.io_fpu_nack_mem = {1{$random}};
    assign core.io_fpu_illegal_rm = {1{$random}};
    assign core.io_fpu_dec_wen = {1{$random}};
    assign core.io_fpu_dec_ren1 = {1{$random}};
    assign core.io_fpu_dec_ren2 = {1{$random}};
    assign core.io_fpu_dec_ren3 = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_invalidate_lr = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_autl_acquire_valid = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_addr_block = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_addr_beat = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_is_builtin_type = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_a_type = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_union = {1{$random}};
    assign core.io_rocc_autl_acquire_bits_data = {4{$random}};
    assign core.io_rocc_autl_grant_ready = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_iptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_iptw_req_bits_store = {1{$random}};
    assign core.io_rocc_iptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_dptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_dptw_req_bits_store = {1{$random}};
    assign core.io_rocc_dptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits_addr = {1{$random}};
    assign core.io_rocc_pptw_req_bits_prv = {1{$random}};
    assign core.io_rocc_pptw_req_bits_store = {1{$random}};
    assign core.io_rocc_pptw_req_bits_fetch = {1{$random}};
    assign core.io_rocc_fpu_req_valid = {1{$random}};
    assign core.io_rocc_fpu_req_bits_cmd = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ldst = {1{$random}};
    assign core.io_rocc_fpu_req_bits_wen = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren1 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren2 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_ren3 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_swap12 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_swap23 = {1{$random}};
    assign core.io_rocc_fpu_req_bits_single = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fromint = {1{$random}};
    assign core.io_rocc_fpu_req_bits_toint = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fastpipe = {1{$random}};
    assign core.io_rocc_fpu_req_bits_fma = {1{$random}};
    assign core.io_rocc_fpu_req_bits_div = {1{$random}};
    assign core.io_rocc_fpu_req_bits_sqrt = {1{$random}};
    assign core.io_rocc_fpu_req_bits_round = {1{$random}};
    assign core.io_rocc_fpu_req_bits_wflags = {1{$random}};
    assign core.io_rocc_fpu_req_bits_rm = {1{$random}};
    assign core.io_rocc_fpu_req_bits_typ = {1{$random}};
    assign core.io_rocc_fpu_req_bits_in1 = {3{$random}};
    assign core.io_rocc_fpu_req_bits_in2 = {3{$random}};
    assign core.io_rocc_fpu_req_bits_in3 = {3{$random}};
    assign core.io_rocc_fpu_resp_ready = {1{$random}};
    assign core.io_rocc_dma_req_valid = {1{$random}};
    assign core.io_rocc_dma_req_bits_client_xact_id = {1{$random}};
    assign core.io_rocc_dma_req_bits_cmd = {1{$random}};
    assign core.io_rocc_dma_req_bits_source = {1{$random}};
    assign core.io_rocc_dma_req_bits_dest = {1{$random}};
    assign core.io_rocc_dma_req_bits_length = {1{$random}};
    assign core.io_rocc_dma_resp_ready = {1{$random}};
// synthesis translate_on
`endif
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data_0( icache_io_cpu_resp_bits_data_0 ),
       .io_cpu_resp_bits_mask( icache_io_cpu_resp_bits_mask ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_mask( icache_io_cpu_btb_resp_bits_mask ),
       .io_cpu_btb_resp_bits_bridx( icache_io_cpu_btb_resp_bits_bridx ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_history( icache_io_cpu_btb_resp_bits_bht_history ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_mask( core_io_imem_btb_update_bits_prediction_bits_mask ),
       .io_cpu_btb_update_bits_prediction_bits_bridx( core_io_imem_btb_update_bits_prediction_bits_bridx ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_history( core_io_imem_btb_update_bits_prediction_bits_bht_history ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       //.io_cpu_btb_update_bits_taken(  )
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_br_pc( core_io_imem_btb_update_bits_br_pc ),
       .io_cpu_bht_update_valid( core_io_imem_bht_update_valid ),
       .io_cpu_bht_update_bits_prediction_valid( core_io_imem_bht_update_bits_prediction_valid ),
       .io_cpu_bht_update_bits_prediction_bits_taken( core_io_imem_bht_update_bits_prediction_bits_taken ),
       .io_cpu_bht_update_bits_prediction_bits_mask( core_io_imem_bht_update_bits_prediction_bits_mask ),
       .io_cpu_bht_update_bits_prediction_bits_bridx( core_io_imem_bht_update_bits_prediction_bits_bridx ),
       .io_cpu_bht_update_bits_prediction_bits_target( core_io_imem_bht_update_bits_prediction_bits_target ),
       .io_cpu_bht_update_bits_prediction_bits_entry( core_io_imem_bht_update_bits_prediction_bits_entry ),
       .io_cpu_bht_update_bits_prediction_bits_bht_history( core_io_imem_bht_update_bits_prediction_bits_bht_history ),
       .io_cpu_bht_update_bits_prediction_bits_bht_value( core_io_imem_bht_update_bits_prediction_bits_bht_value ),
       .io_cpu_bht_update_bits_pc( core_io_imem_bht_update_bits_pc ),
       .io_cpu_bht_update_bits_taken( core_io_imem_bht_update_bits_taken ),
       .io_cpu_bht_update_bits_mispredict( core_io_imem_bht_update_bits_mispredict ),
       .io_cpu_ras_update_valid( core_io_imem_ras_update_valid ),
       .io_cpu_ras_update_bits_isCall( core_io_imem_ras_update_bits_isCall ),
       .io_cpu_ras_update_bits_isReturn( core_io_imem_ras_update_bits_isReturn ),
       .io_cpu_ras_update_bits_returnAddr( core_io_imem_ras_update_bits_returnAddr ),
       .io_cpu_ras_update_bits_prediction_valid( core_io_imem_ras_update_bits_prediction_valid ),
       .io_cpu_ras_update_bits_prediction_bits_taken( core_io_imem_ras_update_bits_prediction_bits_taken ),
       .io_cpu_ras_update_bits_prediction_bits_mask( core_io_imem_ras_update_bits_prediction_bits_mask ),
       .io_cpu_ras_update_bits_prediction_bits_bridx( core_io_imem_ras_update_bits_prediction_bits_bridx ),
       .io_cpu_ras_update_bits_prediction_bits_target( core_io_imem_ras_update_bits_prediction_bits_target ),
       .io_cpu_ras_update_bits_prediction_bits_entry( core_io_imem_ras_update_bits_prediction_bits_entry ),
       .io_cpu_ras_update_bits_prediction_bits_bht_history( core_io_imem_ras_update_bits_prediction_bits_bht_history ),
       .io_cpu_ras_update_bits_prediction_bits_bht_value( core_io_imem_ras_update_bits_prediction_bits_bht_value ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_cpu_npc( icache_io_cpu_npc ),
       .io_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_ptw_req_valid( icache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_0_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_0_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_0_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_0_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_0_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_acquire_ready( io_uncached_0_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( icache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( icache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( icache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( icache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( icache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( icache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( icache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_uncached_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_uncached_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_uncached_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_uncached_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_uncached_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_uncached_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_uncached_0_grant_bits_data )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign icache.io_cpu_btb_update_bits_taken = {1{$random}};
// synthesis translate_on
`endif
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_ptw_req_valid( dcache_io_ptw_req_valid ),
       .io_ptw_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_ptw_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_ptw_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_ptw_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_ptw_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_ptw_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_ptw_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_ptw_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_ptw_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_ptw_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_ptw_status_sd( ptw_io_requestor_1_status_sd ),
       .io_ptw_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_ptw_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_ptw_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_ptw_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_ptw_status_xs( ptw_io_requestor_1_status_xs ),
       .io_ptw_status_fs( ptw_io_requestor_1_status_fs ),
       .io_ptw_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_ptw_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_ptw_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_ptw_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_ptw_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_ptw_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_ptw_status_prv( ptw_io_requestor_1_status_prv ),
       .io_ptw_status_ie( ptw_io_requestor_1_status_ie ),
       .io_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_mem_acquire_ready( io_cached_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_addr_block( dcache_io_mem_acquire_bits_addr_block ),
       .io_mem_acquire_bits_client_xact_id( dcache_io_mem_acquire_bits_client_xact_id ),
       .io_mem_acquire_bits_addr_beat( dcache_io_mem_acquire_bits_addr_beat ),
       .io_mem_acquire_bits_is_builtin_type( dcache_io_mem_acquire_bits_is_builtin_type ),
       .io_mem_acquire_bits_a_type( dcache_io_mem_acquire_bits_a_type ),
       .io_mem_acquire_bits_union( dcache_io_mem_acquire_bits_union ),
       .io_mem_acquire_bits_data( dcache_io_mem_acquire_bits_data ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_cached_0_grant_valid ),
       .io_mem_grant_bits_addr_beat( io_cached_0_grant_bits_addr_beat ),
       .io_mem_grant_bits_client_xact_id( io_cached_0_grant_bits_client_xact_id ),
       .io_mem_grant_bits_manager_xact_id( io_cached_0_grant_bits_manager_xact_id ),
       .io_mem_grant_bits_is_builtin_type( io_cached_0_grant_bits_is_builtin_type ),
       .io_mem_grant_bits_g_type( io_cached_0_grant_bits_g_type ),
       .io_mem_grant_bits_data( io_cached_0_grant_bits_data ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_cached_0_probe_valid ),
       .io_mem_probe_bits_addr_block( io_cached_0_probe_bits_addr_block ),
       .io_mem_probe_bits_p_type( io_cached_0_probe_bits_p_type ),
       .io_mem_release_ready( io_cached_0_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_addr_beat( dcache_io_mem_release_bits_addr_beat ),
       .io_mem_release_bits_addr_block( dcache_io_mem_release_bits_addr_block ),
       .io_mem_release_bits_client_xact_id( dcache_io_mem_release_bits_client_xact_id ),
       .io_mem_release_bits_voluntary( dcache_io_mem_release_bits_voluntary ),
       .io_mem_release_bits_r_type( dcache_io_mem_release_bits_r_type ),
       .io_mem_release_bits_data( dcache_io_mem_release_bits_data )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_ptw_req_valid ),
       .io_requestor_1_req_bits_addr( dcache_io_ptw_req_bits_addr ),
       .io_requestor_1_req_bits_prv( dcache_io_ptw_req_bits_prv ),
       .io_requestor_1_req_bits_store( dcache_io_ptw_req_bits_store ),
       .io_requestor_1_req_bits_fetch( dcache_io_ptw_req_bits_fetch ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_pte_ppn( ptw_io_requestor_1_resp_bits_pte_ppn ),
       .io_requestor_1_resp_bits_pte_reserved_for_software( ptw_io_requestor_1_resp_bits_pte_reserved_for_software ),
       .io_requestor_1_resp_bits_pte_d( ptw_io_requestor_1_resp_bits_pte_d ),
       .io_requestor_1_resp_bits_pte_r( ptw_io_requestor_1_resp_bits_pte_r ),
       .io_requestor_1_resp_bits_pte_typ( ptw_io_requestor_1_resp_bits_pte_typ ),
       .io_requestor_1_resp_bits_pte_v( ptw_io_requestor_1_resp_bits_pte_v ),
       .io_requestor_1_status_sd( ptw_io_requestor_1_status_sd ),
       .io_requestor_1_status_zero2( ptw_io_requestor_1_status_zero2 ),
       .io_requestor_1_status_sd_rv32( ptw_io_requestor_1_status_sd_rv32 ),
       .io_requestor_1_status_zero1( ptw_io_requestor_1_status_zero1 ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_mprv( ptw_io_requestor_1_status_mprv ),
       .io_requestor_1_status_xs( ptw_io_requestor_1_status_xs ),
       .io_requestor_1_status_fs( ptw_io_requestor_1_status_fs ),
       .io_requestor_1_status_prv3( ptw_io_requestor_1_status_prv3 ),
       .io_requestor_1_status_ie3( ptw_io_requestor_1_status_ie3 ),
       .io_requestor_1_status_prv2( ptw_io_requestor_1_status_prv2 ),
       .io_requestor_1_status_ie2( ptw_io_requestor_1_status_ie2 ),
       .io_requestor_1_status_prv1( ptw_io_requestor_1_status_prv1 ),
       .io_requestor_1_status_ie1( ptw_io_requestor_1_status_ie1 ),
       .io_requestor_1_status_prv( ptw_io_requestor_1_status_prv ),
       .io_requestor_1_status_ie( ptw_io_requestor_1_status_ie ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_ptw_req_valid ),
       .io_requestor_0_req_bits_addr( icache_io_ptw_req_bits_addr ),
       .io_requestor_0_req_bits_prv( icache_io_ptw_req_bits_prv ),
       .io_requestor_0_req_bits_store( icache_io_ptw_req_bits_store ),
       .io_requestor_0_req_bits_fetch( icache_io_ptw_req_bits_fetch ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_pte_ppn( ptw_io_requestor_0_resp_bits_pte_ppn ),
       .io_requestor_0_resp_bits_pte_reserved_for_software( ptw_io_requestor_0_resp_bits_pte_reserved_for_software ),
       .io_requestor_0_resp_bits_pte_d( ptw_io_requestor_0_resp_bits_pte_d ),
       .io_requestor_0_resp_bits_pte_r( ptw_io_requestor_0_resp_bits_pte_r ),
       .io_requestor_0_resp_bits_pte_typ( ptw_io_requestor_0_resp_bits_pte_typ ),
       .io_requestor_0_resp_bits_pte_v( ptw_io_requestor_0_resp_bits_pte_v ),
       .io_requestor_0_status_sd( ptw_io_requestor_0_status_sd ),
       .io_requestor_0_status_zero2( ptw_io_requestor_0_status_zero2 ),
       .io_requestor_0_status_sd_rv32( ptw_io_requestor_0_status_sd_rv32 ),
       .io_requestor_0_status_zero1( ptw_io_requestor_0_status_zero1 ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_mprv( ptw_io_requestor_0_status_mprv ),
       .io_requestor_0_status_xs( ptw_io_requestor_0_status_xs ),
       .io_requestor_0_status_fs( ptw_io_requestor_0_status_fs ),
       .io_requestor_0_status_prv3( ptw_io_requestor_0_status_prv3 ),
       .io_requestor_0_status_ie3( ptw_io_requestor_0_status_ie3 ),
       .io_requestor_0_status_prv2( ptw_io_requestor_0_status_prv2 ),
       .io_requestor_0_status_ie2( ptw_io_requestor_0_status_ie2 ),
       .io_requestor_0_status_prv1( ptw_io_requestor_0_status_prv1 ),
       .io_requestor_0_status_ie1( ptw_io_requestor_0_status_ie1 ),
       .io_requestor_0_status_prv( ptw_io_requestor_0_status_prv ),
       .io_requestor_0_status_ie( ptw_io_requestor_0_status_ie ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_status_sd( core_io_ptw_status_sd ),
       .io_dpath_status_zero2( core_io_ptw_status_zero2 ),
       .io_dpath_status_sd_rv32( core_io_ptw_status_sd_rv32 ),
       .io_dpath_status_zero1( core_io_ptw_status_zero1 ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_mprv( core_io_ptw_status_mprv ),
       .io_dpath_status_xs( core_io_ptw_status_xs ),
       .io_dpath_status_fs( core_io_ptw_status_fs ),
       .io_dpath_status_prv3( core_io_ptw_status_prv3 ),
       .io_dpath_status_ie3( core_io_ptw_status_ie3 ),
       .io_dpath_status_prv2( core_io_ptw_status_prv2 ),
       .io_dpath_status_ie2( core_io_ptw_status_ie2 ),
       .io_dpath_status_prv1( core_io_ptw_status_prv1 ),
       .io_dpath_status_ie1( core_io_ptw_status_ie1 ),
       .io_dpath_status_prv( core_io_ptw_status_prv ),
       .io_dpath_status_ie( core_io_ptw_status_ie )
  );
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data_word_bypass( dcArb_io_requestor_1_resp_bits_data_word_bypass ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       .io_requestor_1_invalidate_lr( core_io_dmem_invalidate_lr ),
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_data( ptw_io_mem_req_bits_data ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data_word_bypass( dcArb_io_requestor_0_resp_bits_data_word_bypass ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_invalidate_lr(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data_word_bypass( dcache_io_cpu_resp_bits_data_word_bypass ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_invalidate_lr(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
// synthesis translate_on
`endif
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [11:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[11:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T21;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T22;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T23;
  wire T8;
  wire T9;
  wire[63:0] T10;
  wire[76:0] T11;
  reg [76:0] ram [1:0];
  wire[76:0] T12;
  wire[76:0] T13;
  wire[76:0] T14;
  wire[75:0] T15;
  wire[11:0] T16;
  wire T17;
  wire T18;
  wire empty;
  wire T19;
  wire T20;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T21 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T22 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T23 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_data = T10;
  assign T10 = T11[6'h3f:1'h0];
  assign T11 = ram[R1];
  assign T13 = T14;
  assign T14 = {io_enq_bits_rw, T15};
  assign T15 = {io_enq_bits_addr, io_enq_bits_data};
  assign io_deq_bits_addr = T16;
  assign T16 = T11[7'h4b:7'h40];
  assign io_deq_bits_rw = T17;
  assign T17 = T11[7'h4c:7'h4c];
  assign io_deq_valid = T18;
  assign T18 = empty ^ 1'h1;
  assign empty = ptr_match & T19;
  assign T19 = maybe_full ^ 1'h1;
  assign io_enq_ready = T20;
  assign T20 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= T13;
  end
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T15;
  wire T2;
  wire T3;
  wire do_deq;
  reg  R4;
  wire T16;
  wire T5;
  wire T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T17;
  wire T8;
  wire T9;
  wire[63:0] T10;
  reg [63:0] ram [1:0];
  wire[63:0] T11;
  wire T12;
  wire empty;
  wire T13;
  wire T14;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R4 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T15 = reset ? 1'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T16 = reset ? 1'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T17 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits = T10;
  assign T10 = ram[R1];
  assign io_deq_valid = T12;
  assign T12 = empty ^ 1'h1;
  assign empty = ptr_match & T13;
  assign T13 = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 1'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits;
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_csr,
    input  io_mem_backup_ctrl_en,
    input  io_mem_backup_ctrl_in_valid,
    input  io_mem_backup_ctrl_out_ready,
    output io_mem_backup_ctrl_out_valid,
    input  io_mem_0_aw_ready,
    output io_mem_0_aw_valid,
    output[31:0] io_mem_0_aw_bits_addr,
    output[7:0] io_mem_0_aw_bits_len,
    output[2:0] io_mem_0_aw_bits_size,
    output[1:0] io_mem_0_aw_bits_burst,
    output io_mem_0_aw_bits_lock,
    output[3:0] io_mem_0_aw_bits_cache,
    output[2:0] io_mem_0_aw_bits_prot,
    output[3:0] io_mem_0_aw_bits_qos,
    output[3:0] io_mem_0_aw_bits_region,
    output[3:0] io_mem_0_aw_bits_id,
    output io_mem_0_aw_bits_user,
    input  io_mem_0_w_ready,
    output io_mem_0_w_valid,
    output[63:0] io_mem_0_w_bits_data,
    output io_mem_0_w_bits_last,
    output[7:0] io_mem_0_w_bits_strb,
    output io_mem_0_w_bits_user,
    output io_mem_0_b_ready,
    input  io_mem_0_b_valid,
    input [1:0] io_mem_0_b_bits_resp,
    input [3:0] io_mem_0_b_bits_id,
    input  io_mem_0_b_bits_user,
    input  io_mem_0_ar_ready,
    output io_mem_0_ar_valid,
    output[31:0] io_mem_0_ar_bits_addr,
    output[7:0] io_mem_0_ar_bits_len,
    output[2:0] io_mem_0_ar_bits_size,
    output[1:0] io_mem_0_ar_bits_burst,
    output io_mem_0_ar_bits_lock,
    output[3:0] io_mem_0_ar_bits_cache,
    output[2:0] io_mem_0_ar_bits_prot,
    output[3:0] io_mem_0_ar_bits_qos,
    output[3:0] io_mem_0_ar_bits_region,
    output[3:0] io_mem_0_ar_bits_id,
    output io_mem_0_ar_bits_user,
    output io_mem_0_r_ready,
    input  io_mem_0_r_valid,
    input [1:0] io_mem_0_r_bits_resp,
    input [63:0] io_mem_0_r_bits_data,
    input  io_mem_0_r_bits_last,
    input [3:0] io_mem_0_r_bits_id,
    input  io_mem_0_r_bits_user
);

  reg  R0;
  reg  R1;
  wire Queue_io_enq_ready;
  wire Queue_io_deq_valid;
  wire Queue_io_deq_bits_rw;
  wire[11:0] Queue_io_deq_bits_addr;
  wire[63:0] Queue_io_deq_bits_data;
  wire Queue_1_io_enq_ready;
  wire Queue_1_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_2_io_enq_ready;
  wire Queue_2_io_deq_valid;
  wire[31:0] Queue_2_io_deq_bits_addr;
  wire[7:0] Queue_2_io_deq_bits_len;
  wire[2:0] Queue_2_io_deq_bits_size;
  wire[1:0] Queue_2_io_deq_bits_burst;
  wire Queue_2_io_deq_bits_lock;
  wire[2:0] Queue_2_io_deq_bits_prot;
  wire[3:0] Queue_2_io_deq_bits_qos;
  wire[3:0] Queue_2_io_deq_bits_region;
  wire[3:0] Queue_2_io_deq_bits_id;
  wire Queue_2_io_deq_bits_user;
  wire Queue_3_io_enq_ready;
  wire Queue_3_io_deq_valid;
  wire[31:0] Queue_3_io_deq_bits_addr;
  wire[7:0] Queue_3_io_deq_bits_len;
  wire[2:0] Queue_3_io_deq_bits_size;
  wire[1:0] Queue_3_io_deq_bits_burst;
  wire Queue_3_io_deq_bits_lock;
  wire[2:0] Queue_3_io_deq_bits_prot;
  wire[3:0] Queue_3_io_deq_bits_qos;
  wire[3:0] Queue_3_io_deq_bits_region;
  wire[3:0] Queue_3_io_deq_bits_id;
  wire Queue_3_io_deq_bits_user;
  wire Queue_4_io_enq_ready;
  wire Queue_4_io_deq_valid;
  wire[63:0] Queue_4_io_deq_bits_data;
  wire Queue_4_io_deq_bits_last;
  wire[7:0] Queue_4_io_deq_bits_strb;
  wire Queue_4_io_deq_bits_user;
  wire Queue_5_io_enq_ready;
  wire Queue_5_io_deq_valid;
  wire[1:0] Queue_5_io_deq_bits_resp;
  wire[63:0] Queue_5_io_deq_bits_data;
  wire Queue_5_io_deq_bits_last;
  wire[3:0] Queue_5_io_deq_bits_id;
  wire Queue_5_io_deq_bits_user;
  wire Queue_6_io_enq_ready;
  wire Queue_6_io_deq_valid;
  wire[1:0] Queue_6_io_deq_bits_resp;
  wire[3:0] Queue_6_io_deq_bits_id;
  wire Queue_6_io_deq_bits_user;
  wire errslave_io_aw_ready;
  wire errslave_io_w_ready;
  wire errslave_io_b_valid;
  wire[1:0] errslave_io_b_bits_resp;
  wire[3:0] errslave_io_b_bits_id;
  wire errslave_io_ar_ready;
  wire errslave_io_r_valid;
  wire[1:0] errslave_io_r_bits_resp;
  wire[63:0] errslave_io_r_bits_data;
  wire errslave_io_r_bits_last;
  wire[3:0] errslave_io_r_bits_id;
  wire RocketTile_io_cached_0_acquire_valid;
  wire[25:0] RocketTile_io_cached_0_acquire_bits_addr_block;
  wire[1:0] RocketTile_io_cached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_cached_0_acquire_bits_addr_beat;
  wire RocketTile_io_cached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_cached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_cached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_cached_0_acquire_bits_data;
  wire RocketTile_io_cached_0_grant_ready;
  wire RocketTile_io_cached_0_probe_ready;
  wire RocketTile_io_cached_0_release_valid;
  wire[1:0] RocketTile_io_cached_0_release_bits_addr_beat;
  wire[25:0] RocketTile_io_cached_0_release_bits_addr_block;
  wire[1:0] RocketTile_io_cached_0_release_bits_client_xact_id;
  wire RocketTile_io_cached_0_release_bits_voluntary;
  wire[2:0] RocketTile_io_cached_0_release_bits_r_type;
  wire[127:0] RocketTile_io_cached_0_release_bits_data;
  wire RocketTile_io_uncached_0_acquire_valid;
  wire[25:0] RocketTile_io_uncached_0_acquire_bits_addr_block;
  wire[1:0] RocketTile_io_uncached_0_acquire_bits_client_xact_id;
  wire[1:0] RocketTile_io_uncached_0_acquire_bits_addr_beat;
  wire RocketTile_io_uncached_0_acquire_bits_is_builtin_type;
  wire[2:0] RocketTile_io_uncached_0_acquire_bits_a_type;
  wire[16:0] RocketTile_io_uncached_0_acquire_bits_union;
  wire[127:0] RocketTile_io_uncached_0_acquire_bits_data;
  wire RocketTile_io_uncached_0_grant_ready;
  wire RocketTile_io_host_csr_req_ready;
  wire RocketTile_io_host_csr_resp_valid;
  wire[63:0] RocketTile_io_host_csr_resp_bits;
  wire RocketTile_io_host_debug_stats_csr;
  wire uncore_io_host_in_ready;
  wire uncore_io_host_out_valid;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_debug_stats_csr;
  wire uncore_io_mem_0_aw_valid;
  wire[31:0] uncore_io_mem_0_aw_bits_addr;
  wire[7:0] uncore_io_mem_0_aw_bits_len;
  wire[2:0] uncore_io_mem_0_aw_bits_size;
  wire[1:0] uncore_io_mem_0_aw_bits_burst;
  wire uncore_io_mem_0_aw_bits_lock;
  wire[3:0] uncore_io_mem_0_aw_bits_cache;
  wire[2:0] uncore_io_mem_0_aw_bits_prot;
  wire[3:0] uncore_io_mem_0_aw_bits_qos;
  wire[3:0] uncore_io_mem_0_aw_bits_region;
  wire[3:0] uncore_io_mem_0_aw_bits_id;
  wire uncore_io_mem_0_aw_bits_user;
  wire uncore_io_mem_0_w_valid;
  wire[63:0] uncore_io_mem_0_w_bits_data;
  wire uncore_io_mem_0_w_bits_last;
  wire[7:0] uncore_io_mem_0_w_bits_strb;
  wire uncore_io_mem_0_w_bits_user;
  wire uncore_io_mem_0_b_ready;
  wire uncore_io_mem_0_ar_valid;
  wire[31:0] uncore_io_mem_0_ar_bits_addr;
  wire[7:0] uncore_io_mem_0_ar_bits_len;
  wire[2:0] uncore_io_mem_0_ar_bits_size;
  wire[1:0] uncore_io_mem_0_ar_bits_burst;
  wire uncore_io_mem_0_ar_bits_lock;
  wire[3:0] uncore_io_mem_0_ar_bits_cache;
  wire[2:0] uncore_io_mem_0_ar_bits_prot;
  wire[3:0] uncore_io_mem_0_ar_bits_qos;
  wire[3:0] uncore_io_mem_0_ar_bits_region;
  wire[3:0] uncore_io_mem_0_ar_bits_id;
  wire uncore_io_mem_0_ar_bits_user;
  wire uncore_io_mem_0_r_ready;
  wire uncore_io_tiles_cached_0_acquire_ready;
  wire uncore_io_tiles_cached_0_grant_valid;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire[1:0] uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire[2:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire uncore_io_tiles_cached_0_probe_valid;
  wire[25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire[1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire uncore_io_tiles_cached_0_release_ready;
  wire uncore_io_tiles_uncached_0_acquire_ready;
  wire uncore_io_tiles_uncached_0_grant_valid;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire[1:0] uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire[2:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire[3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire[127:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire uncore_io_htif_0_reset;
  wire uncore_io_htif_0_csr_req_valid;
  wire uncore_io_htif_0_csr_req_bits_rw;
  wire[11:0] uncore_io_htif_0_csr_req_bits_addr;
  wire[63:0] uncore_io_htif_0_csr_req_bits_data;
  wire uncore_io_htif_0_csr_resp_ready;
  wire uncore_io_mmio_aw_valid;
  wire[31:0] uncore_io_mmio_aw_bits_addr;
  wire[7:0] uncore_io_mmio_aw_bits_len;
  wire[2:0] uncore_io_mmio_aw_bits_size;
  wire[1:0] uncore_io_mmio_aw_bits_burst;
  wire uncore_io_mmio_aw_bits_lock;
  wire[3:0] uncore_io_mmio_aw_bits_cache;
  wire[2:0] uncore_io_mmio_aw_bits_prot;
  wire[3:0] uncore_io_mmio_aw_bits_qos;
  wire[3:0] uncore_io_mmio_aw_bits_region;
  wire[3:0] uncore_io_mmio_aw_bits_id;
  wire uncore_io_mmio_aw_bits_user;
  wire uncore_io_mmio_w_valid;
  wire[63:0] uncore_io_mmio_w_bits_data;
  wire uncore_io_mmio_w_bits_last;
  wire[7:0] uncore_io_mmio_w_bits_strb;
  wire uncore_io_mmio_w_bits_user;
  wire uncore_io_mmio_b_ready;
  wire uncore_io_mmio_ar_valid;
  wire[31:0] uncore_io_mmio_ar_bits_addr;
  wire[7:0] uncore_io_mmio_ar_bits_len;
  wire[2:0] uncore_io_mmio_ar_bits_size;
  wire[1:0] uncore_io_mmio_ar_bits_burst;
  wire uncore_io_mmio_ar_bits_lock;
  wire[3:0] uncore_io_mmio_ar_bits_cache;
  wire[2:0] uncore_io_mmio_ar_bits_prot;
  wire[3:0] uncore_io_mmio_ar_bits_qos;
  wire[3:0] uncore_io_mmio_ar_bits_region;
  wire[3:0] uncore_io_mmio_ar_bits_id;
  wire uncore_io_mmio_ar_bits_user;
  wire uncore_io_mmio_r_ready;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_mem_backup_ctrl_out_valid = {1{$random}};
//  assign io_host_clk_edge = {1{$random}};
//  assign io_host_clk = {1{$random}};
// synthesis translate_on
`endif
  assign io_mem_0_r_ready = Queue_5_io_enq_ready;
  assign io_mem_0_ar_bits_user = Queue_2_io_deq_bits_user;
  assign io_mem_0_ar_bits_id = Queue_2_io_deq_bits_id;
  assign io_mem_0_ar_bits_region = Queue_2_io_deq_bits_region;
  assign io_mem_0_ar_bits_qos = Queue_2_io_deq_bits_qos;
  assign io_mem_0_ar_bits_prot = Queue_2_io_deq_bits_prot;
  assign io_mem_0_ar_bits_cache = 4'h3;
  assign io_mem_0_ar_bits_lock = Queue_2_io_deq_bits_lock;
  assign io_mem_0_ar_bits_burst = Queue_2_io_deq_bits_burst;
  assign io_mem_0_ar_bits_size = Queue_2_io_deq_bits_size;
  assign io_mem_0_ar_bits_len = Queue_2_io_deq_bits_len;
  assign io_mem_0_ar_bits_addr = Queue_2_io_deq_bits_addr;
  assign io_mem_0_ar_valid = Queue_2_io_deq_valid;
  assign io_mem_0_b_ready = Queue_6_io_enq_ready;
  assign io_mem_0_w_bits_user = Queue_4_io_deq_bits_user;
  assign io_mem_0_w_bits_strb = Queue_4_io_deq_bits_strb;
  assign io_mem_0_w_bits_last = Queue_4_io_deq_bits_last;
  assign io_mem_0_w_bits_data = Queue_4_io_deq_bits_data;
  assign io_mem_0_w_valid = Queue_4_io_deq_valid;
  assign io_mem_0_aw_bits_user = Queue_3_io_deq_bits_user;
  assign io_mem_0_aw_bits_id = Queue_3_io_deq_bits_id;
  assign io_mem_0_aw_bits_region = Queue_3_io_deq_bits_region;
  assign io_mem_0_aw_bits_qos = Queue_3_io_deq_bits_qos;
  assign io_mem_0_aw_bits_prot = Queue_3_io_deq_bits_prot;
  assign io_mem_0_aw_bits_cache = 4'h3;
  assign io_mem_0_aw_bits_lock = Queue_3_io_deq_bits_lock;
  assign io_mem_0_aw_bits_burst = Queue_3_io_deq_bits_burst;
  assign io_mem_0_aw_bits_size = Queue_3_io_deq_bits_size;
  assign io_mem_0_aw_bits_len = Queue_3_io_deq_bits_len;
  assign io_mem_0_aw_bits_addr = Queue_3_io_deq_bits_addr;
  assign io_mem_0_aw_valid = Queue_3_io_deq_valid;
  assign io_host_debug_stats_csr = uncore_io_host_debug_stats_csr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_csr( uncore_io_host_debug_stats_csr ),
       .io_mem_0_aw_ready( Queue_3_io_enq_ready ),
       .io_mem_0_aw_valid( uncore_io_mem_0_aw_valid ),
       .io_mem_0_aw_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_mem_0_aw_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_mem_0_aw_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_mem_0_aw_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_mem_0_aw_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_mem_0_aw_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_mem_0_aw_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_mem_0_aw_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_mem_0_aw_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_mem_0_aw_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_mem_0_aw_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_mem_0_w_ready( Queue_4_io_enq_ready ),
       .io_mem_0_w_valid( uncore_io_mem_0_w_valid ),
       .io_mem_0_w_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_mem_0_w_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_mem_0_w_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_mem_0_w_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_mem_0_b_ready( uncore_io_mem_0_b_ready ),
       .io_mem_0_b_valid( Queue_6_io_deq_valid ),
       .io_mem_0_b_bits_resp( Queue_6_io_deq_bits_resp ),
       .io_mem_0_b_bits_id( Queue_6_io_deq_bits_id ),
       .io_mem_0_b_bits_user( Queue_6_io_deq_bits_user ),
       .io_mem_0_ar_ready( Queue_2_io_enq_ready ),
       .io_mem_0_ar_valid( uncore_io_mem_0_ar_valid ),
       .io_mem_0_ar_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_mem_0_ar_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_mem_0_ar_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_mem_0_ar_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_mem_0_ar_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_mem_0_ar_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_mem_0_ar_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_mem_0_ar_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_mem_0_ar_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_mem_0_ar_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_mem_0_ar_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_mem_0_r_ready( uncore_io_mem_0_r_ready ),
       .io_mem_0_r_valid( Queue_5_io_deq_valid ),
       .io_mem_0_r_bits_resp( Queue_5_io_deq_bits_resp ),
       .io_mem_0_r_bits_data( Queue_5_io_deq_bits_data ),
       .io_mem_0_r_bits_last( Queue_5_io_deq_bits_last ),
       .io_mem_0_r_bits_id( Queue_5_io_deq_bits_id ),
       .io_mem_0_r_bits_user( Queue_5_io_deq_bits_user ),
       .io_tiles_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_tiles_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_tiles_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_tiles_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_tiles_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_tiles_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_tiles_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_tiles_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_tiles_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_tiles_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_tiles_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_tiles_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_tiles_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_tiles_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_tiles_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_tiles_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_tiles_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_tiles_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_tiles_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_tiles_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_tiles_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_tiles_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_tiles_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_tiles_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_tiles_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_tiles_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_tiles_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_tiles_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_tiles_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_tiles_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_tiles_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_tiles_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_tiles_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_tiles_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_tiles_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_tiles_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_tiles_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_tiles_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_tiles_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_tiles_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_tiles_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_tiles_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_tiles_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_tiles_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_tiles_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_tiles_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_csr_req_ready( Queue_io_enq_ready ),
       .io_htif_0_csr_req_valid( uncore_io_htif_0_csr_req_valid ),
       .io_htif_0_csr_req_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_htif_0_csr_req_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_htif_0_csr_req_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_htif_0_csr_resp_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_htif_0_csr_resp_valid( Queue_1_io_deq_valid ),
       .io_htif_0_csr_resp_bits( Queue_1_io_deq_bits ),
       .io_htif_0_debug_stats_csr( RocketTile_io_host_debug_stats_csr ),
       //.io_mem_backup_ctrl_en(  )
       //.io_mem_backup_ctrl_in_valid(  )
       //.io_mem_backup_ctrl_out_ready(  )
       //.io_mem_backup_ctrl_out_valid(  )
       .io_mmio_aw_ready( errslave_io_aw_ready ),
       .io_mmio_aw_valid( uncore_io_mmio_aw_valid ),
       .io_mmio_aw_bits_addr( uncore_io_mmio_aw_bits_addr ),
       .io_mmio_aw_bits_len( uncore_io_mmio_aw_bits_len ),
       .io_mmio_aw_bits_size( uncore_io_mmio_aw_bits_size ),
       .io_mmio_aw_bits_burst( uncore_io_mmio_aw_bits_burst ),
       .io_mmio_aw_bits_lock( uncore_io_mmio_aw_bits_lock ),
       .io_mmio_aw_bits_cache( uncore_io_mmio_aw_bits_cache ),
       .io_mmio_aw_bits_prot( uncore_io_mmio_aw_bits_prot ),
       .io_mmio_aw_bits_qos( uncore_io_mmio_aw_bits_qos ),
       .io_mmio_aw_bits_region( uncore_io_mmio_aw_bits_region ),
       .io_mmio_aw_bits_id( uncore_io_mmio_aw_bits_id ),
       .io_mmio_aw_bits_user( uncore_io_mmio_aw_bits_user ),
       .io_mmio_w_ready( errslave_io_w_ready ),
       .io_mmio_w_valid( uncore_io_mmio_w_valid ),
       .io_mmio_w_bits_data( uncore_io_mmio_w_bits_data ),
       .io_mmio_w_bits_last( uncore_io_mmio_w_bits_last ),
       .io_mmio_w_bits_strb( uncore_io_mmio_w_bits_strb ),
       .io_mmio_w_bits_user( uncore_io_mmio_w_bits_user ),
       .io_mmio_b_ready( uncore_io_mmio_b_ready ),
       .io_mmio_b_valid( errslave_io_b_valid ),
       .io_mmio_b_bits_resp( errslave_io_b_bits_resp ),
       .io_mmio_b_bits_id( errslave_io_b_bits_id ),
       //.io_mmio_b_bits_user(  )
       .io_mmio_ar_ready( errslave_io_ar_ready ),
       .io_mmio_ar_valid( uncore_io_mmio_ar_valid ),
       .io_mmio_ar_bits_addr( uncore_io_mmio_ar_bits_addr ),
       .io_mmio_ar_bits_len( uncore_io_mmio_ar_bits_len ),
       .io_mmio_ar_bits_size( uncore_io_mmio_ar_bits_size ),
       .io_mmio_ar_bits_burst( uncore_io_mmio_ar_bits_burst ),
       .io_mmio_ar_bits_lock( uncore_io_mmio_ar_bits_lock ),
       .io_mmio_ar_bits_cache( uncore_io_mmio_ar_bits_cache ),
       .io_mmio_ar_bits_prot( uncore_io_mmio_ar_bits_prot ),
       .io_mmio_ar_bits_qos( uncore_io_mmio_ar_bits_qos ),
       .io_mmio_ar_bits_region( uncore_io_mmio_ar_bits_region ),
       .io_mmio_ar_bits_id( uncore_io_mmio_ar_bits_id ),
       .io_mmio_ar_bits_user( uncore_io_mmio_ar_bits_user ),
       .io_mmio_r_ready( uncore_io_mmio_r_ready ),
       .io_mmio_r_valid( errslave_io_r_valid ),
       .io_mmio_r_bits_resp( errslave_io_r_bits_resp ),
       .io_mmio_r_bits_data( errslave_io_r_bits_data ),
       .io_mmio_r_bits_last( errslave_io_r_bits_last ),
       .io_mmio_r_bits_id( errslave_io_r_bits_id )
       //.io_mmio_r_bits_user(  )
       //.io_dma_0_req_ready(  )
       //.io_dma_0_req_valid(  )
       //.io_dma_0_req_bits_client_xact_id(  )
       //.io_dma_0_req_bits_cmd(  )
       //.io_dma_0_req_bits_source(  )
       //.io_dma_0_req_bits_dest(  )
       //.io_dma_0_req_bits_length(  )
       //.io_dma_0_resp_ready(  )
       //.io_dma_0_resp_valid(  )
       //.io_dma_0_resp_bits_client_xact_id(  )
       //.io_dma_0_resp_bits_status(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign uncore.io_mmio_b_bits_user = {1{$random}};
    assign uncore.io_mmio_r_bits_user = {1{$random}};
// synthesis translate_on
`endif
  RocketTile RocketTile(.clk(clk), .reset(uncore_io_htif_0_reset),
       .io_cached_0_acquire_ready( uncore_io_tiles_cached_0_acquire_ready ),
       .io_cached_0_acquire_valid( RocketTile_io_cached_0_acquire_valid ),
       .io_cached_0_acquire_bits_addr_block( RocketTile_io_cached_0_acquire_bits_addr_block ),
       .io_cached_0_acquire_bits_client_xact_id( RocketTile_io_cached_0_acquire_bits_client_xact_id ),
       .io_cached_0_acquire_bits_addr_beat( RocketTile_io_cached_0_acquire_bits_addr_beat ),
       .io_cached_0_acquire_bits_is_builtin_type( RocketTile_io_cached_0_acquire_bits_is_builtin_type ),
       .io_cached_0_acquire_bits_a_type( RocketTile_io_cached_0_acquire_bits_a_type ),
       .io_cached_0_acquire_bits_union( RocketTile_io_cached_0_acquire_bits_union ),
       .io_cached_0_acquire_bits_data( RocketTile_io_cached_0_acquire_bits_data ),
       .io_cached_0_grant_ready( RocketTile_io_cached_0_grant_ready ),
       .io_cached_0_grant_valid( uncore_io_tiles_cached_0_grant_valid ),
       .io_cached_0_grant_bits_addr_beat( uncore_io_tiles_cached_0_grant_bits_addr_beat ),
       .io_cached_0_grant_bits_client_xact_id( uncore_io_tiles_cached_0_grant_bits_client_xact_id ),
       .io_cached_0_grant_bits_manager_xact_id( uncore_io_tiles_cached_0_grant_bits_manager_xact_id ),
       .io_cached_0_grant_bits_is_builtin_type( uncore_io_tiles_cached_0_grant_bits_is_builtin_type ),
       .io_cached_0_grant_bits_g_type( uncore_io_tiles_cached_0_grant_bits_g_type ),
       .io_cached_0_grant_bits_data( uncore_io_tiles_cached_0_grant_bits_data ),
       .io_cached_0_probe_ready( RocketTile_io_cached_0_probe_ready ),
       .io_cached_0_probe_valid( uncore_io_tiles_cached_0_probe_valid ),
       .io_cached_0_probe_bits_addr_block( uncore_io_tiles_cached_0_probe_bits_addr_block ),
       .io_cached_0_probe_bits_p_type( uncore_io_tiles_cached_0_probe_bits_p_type ),
       .io_cached_0_release_ready( uncore_io_tiles_cached_0_release_ready ),
       .io_cached_0_release_valid( RocketTile_io_cached_0_release_valid ),
       .io_cached_0_release_bits_addr_beat( RocketTile_io_cached_0_release_bits_addr_beat ),
       .io_cached_0_release_bits_addr_block( RocketTile_io_cached_0_release_bits_addr_block ),
       .io_cached_0_release_bits_client_xact_id( RocketTile_io_cached_0_release_bits_client_xact_id ),
       .io_cached_0_release_bits_voluntary( RocketTile_io_cached_0_release_bits_voluntary ),
       .io_cached_0_release_bits_r_type( RocketTile_io_cached_0_release_bits_r_type ),
       .io_cached_0_release_bits_data( RocketTile_io_cached_0_release_bits_data ),
       .io_uncached_0_acquire_ready( uncore_io_tiles_uncached_0_acquire_ready ),
       .io_uncached_0_acquire_valid( RocketTile_io_uncached_0_acquire_valid ),
       .io_uncached_0_acquire_bits_addr_block( RocketTile_io_uncached_0_acquire_bits_addr_block ),
       .io_uncached_0_acquire_bits_client_xact_id( RocketTile_io_uncached_0_acquire_bits_client_xact_id ),
       .io_uncached_0_acquire_bits_addr_beat( RocketTile_io_uncached_0_acquire_bits_addr_beat ),
       .io_uncached_0_acquire_bits_is_builtin_type( RocketTile_io_uncached_0_acquire_bits_is_builtin_type ),
       .io_uncached_0_acquire_bits_a_type( RocketTile_io_uncached_0_acquire_bits_a_type ),
       .io_uncached_0_acquire_bits_union( RocketTile_io_uncached_0_acquire_bits_union ),
       .io_uncached_0_acquire_bits_data( RocketTile_io_uncached_0_acquire_bits_data ),
       .io_uncached_0_grant_ready( RocketTile_io_uncached_0_grant_ready ),
       .io_uncached_0_grant_valid( uncore_io_tiles_uncached_0_grant_valid ),
       .io_uncached_0_grant_bits_addr_beat( uncore_io_tiles_uncached_0_grant_bits_addr_beat ),
       .io_uncached_0_grant_bits_client_xact_id( uncore_io_tiles_uncached_0_grant_bits_client_xact_id ),
       .io_uncached_0_grant_bits_manager_xact_id( uncore_io_tiles_uncached_0_grant_bits_manager_xact_id ),
       .io_uncached_0_grant_bits_is_builtin_type( uncore_io_tiles_uncached_0_grant_bits_is_builtin_type ),
       .io_uncached_0_grant_bits_g_type( uncore_io_tiles_uncached_0_grant_bits_g_type ),
       .io_uncached_0_grant_bits_data( uncore_io_tiles_uncached_0_grant_bits_data ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_csr_req_ready( RocketTile_io_host_csr_req_ready ),
       .io_host_csr_req_valid( Queue_io_deq_valid ),
       .io_host_csr_req_bits_rw( Queue_io_deq_bits_rw ),
       .io_host_csr_req_bits_addr( Queue_io_deq_bits_addr ),
       .io_host_csr_req_bits_data( Queue_io_deq_bits_data ),
       .io_host_csr_resp_ready( Queue_1_io_enq_ready ),
       .io_host_csr_resp_valid( RocketTile_io_host_csr_resp_valid ),
       .io_host_csr_resp_bits( RocketTile_io_host_csr_resp_bits ),
       .io_host_debug_stats_csr( RocketTile_io_host_debug_stats_csr )
       //.io_dma_req_ready(  )
       //.io_dma_req_valid(  )
       //.io_dma_req_bits_client_xact_id(  )
       //.io_dma_req_bits_cmd(  )
       //.io_dma_req_bits_source(  )
       //.io_dma_req_bits_dest(  )
       //.io_dma_req_bits_length(  )
       //.io_dma_resp_ready(  )
       //.io_dma_resp_valid(  )
       //.io_dma_resp_bits_client_xact_id(  )
       //.io_dma_resp_bits_status(  )
  );
  Queue_0 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_csr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_csr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_csr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_csr_req_bits_data ),
       .io_deq_ready( RocketTile_io_host_csr_req_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_rw( Queue_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_io_deq_bits_data )
       //.io_count(  )
  );
  Queue_1 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( RocketTile_io_host_csr_resp_valid ),
       .io_enq_bits( RocketTile_io_host_csr_resp_bits ),
       .io_deq_ready( uncore_io_htif_0_csr_resp_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
       //.io_count(  )
  );
  Queue_2 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_ar_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_ar_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_ar_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_ar_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_ar_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_ar_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_ar_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_ar_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_ar_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_ar_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_ar_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_ar_bits_user ),
       .io_deq_ready( io_mem_0_ar_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_addr( Queue_2_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_2_io_deq_bits_len ),
       .io_deq_bits_size( Queue_2_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_2_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_2_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_2_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_2_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_2_io_deq_bits_region ),
       .io_deq_bits_id( Queue_2_io_deq_bits_id ),
       .io_deq_bits_user( Queue_2_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_2 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_aw_valid ),
       .io_enq_bits_addr( uncore_io_mem_0_aw_bits_addr ),
       .io_enq_bits_len( uncore_io_mem_0_aw_bits_len ),
       .io_enq_bits_size( uncore_io_mem_0_aw_bits_size ),
       .io_enq_bits_burst( uncore_io_mem_0_aw_bits_burst ),
       .io_enq_bits_lock( uncore_io_mem_0_aw_bits_lock ),
       .io_enq_bits_cache( uncore_io_mem_0_aw_bits_cache ),
       .io_enq_bits_prot( uncore_io_mem_0_aw_bits_prot ),
       .io_enq_bits_qos( uncore_io_mem_0_aw_bits_qos ),
       .io_enq_bits_region( uncore_io_mem_0_aw_bits_region ),
       .io_enq_bits_id( uncore_io_mem_0_aw_bits_id ),
       .io_enq_bits_user( uncore_io_mem_0_aw_bits_user ),
       .io_deq_ready( io_mem_0_aw_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_addr( Queue_3_io_deq_bits_addr ),
       .io_deq_bits_len( Queue_3_io_deq_bits_len ),
       .io_deq_bits_size( Queue_3_io_deq_bits_size ),
       .io_deq_bits_burst( Queue_3_io_deq_bits_burst ),
       .io_deq_bits_lock( Queue_3_io_deq_bits_lock ),
       //.io_deq_bits_cache(  )
       .io_deq_bits_prot( Queue_3_io_deq_bits_prot ),
       .io_deq_bits_qos( Queue_3_io_deq_bits_qos ),
       .io_deq_bits_region( Queue_3_io_deq_bits_region ),
       .io_deq_bits_id( Queue_3_io_deq_bits_id ),
       .io_deq_bits_user( Queue_3_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_3 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( uncore_io_mem_0_w_valid ),
       .io_enq_bits_data( uncore_io_mem_0_w_bits_data ),
       .io_enq_bits_last( uncore_io_mem_0_w_bits_last ),
       .io_enq_bits_strb( uncore_io_mem_0_w_bits_strb ),
       .io_enq_bits_user( uncore_io_mem_0_w_bits_user ),
       .io_deq_ready( io_mem_0_w_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_data( Queue_4_io_deq_bits_data ),
       .io_deq_bits_last( Queue_4_io_deq_bits_last ),
       .io_deq_bits_strb( Queue_4_io_deq_bits_strb ),
       .io_deq_bits_user( Queue_4_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_4 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( io_mem_0_r_valid ),
       .io_enq_bits_resp( io_mem_0_r_bits_resp ),
       .io_enq_bits_data( io_mem_0_r_bits_data ),
       .io_enq_bits_last( io_mem_0_r_bits_last ),
       .io_enq_bits_id( io_mem_0_r_bits_id ),
       .io_enq_bits_user( io_mem_0_r_bits_user ),
       .io_deq_ready( uncore_io_mem_0_r_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_resp( Queue_5_io_deq_bits_resp ),
       .io_deq_bits_data( Queue_5_io_deq_bits_data ),
       .io_deq_bits_last( Queue_5_io_deq_bits_last ),
       .io_deq_bits_id( Queue_5_io_deq_bits_id ),
       .io_deq_bits_user( Queue_5_io_deq_bits_user )
       //.io_count(  )
  );
  Queue_5 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( io_mem_0_b_valid ),
       .io_enq_bits_resp( io_mem_0_b_bits_resp ),
       .io_enq_bits_id( io_mem_0_b_bits_id ),
       .io_enq_bits_user( io_mem_0_b_bits_user ),
       .io_deq_ready( uncore_io_mem_0_b_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_resp( Queue_6_io_deq_bits_resp ),
       .io_deq_bits_id( Queue_6_io_deq_bits_id ),
       .io_deq_bits_user( Queue_6_io_deq_bits_user )
       //.io_count(  )
  );
  NastiErrorSlave errslave(.clk(clk), .reset(reset),
       .io_aw_ready( errslave_io_aw_ready ),
       .io_aw_valid( uncore_io_mmio_aw_valid ),
       .io_aw_bits_addr( uncore_io_mmio_aw_bits_addr ),
       .io_aw_bits_len( uncore_io_mmio_aw_bits_len ),
       .io_aw_bits_size( uncore_io_mmio_aw_bits_size ),
       .io_aw_bits_burst( uncore_io_mmio_aw_bits_burst ),
       .io_aw_bits_lock( uncore_io_mmio_aw_bits_lock ),
       .io_aw_bits_cache( uncore_io_mmio_aw_bits_cache ),
       .io_aw_bits_prot( uncore_io_mmio_aw_bits_prot ),
       .io_aw_bits_qos( uncore_io_mmio_aw_bits_qos ),
       .io_aw_bits_region( uncore_io_mmio_aw_bits_region ),
       .io_aw_bits_id( uncore_io_mmio_aw_bits_id ),
       .io_aw_bits_user( uncore_io_mmio_aw_bits_user ),
       .io_w_ready( errslave_io_w_ready ),
       .io_w_valid( uncore_io_mmio_w_valid ),
       .io_w_bits_data( uncore_io_mmio_w_bits_data ),
       .io_w_bits_last( uncore_io_mmio_w_bits_last ),
       .io_w_bits_strb( uncore_io_mmio_w_bits_strb ),
       .io_w_bits_user( uncore_io_mmio_w_bits_user ),
       .io_b_ready( uncore_io_mmio_b_ready ),
       .io_b_valid( errslave_io_b_valid ),
       .io_b_bits_resp( errslave_io_b_bits_resp ),
       .io_b_bits_id( errslave_io_b_bits_id ),
       //.io_b_bits_user(  )
       .io_ar_ready( errslave_io_ar_ready ),
       .io_ar_valid( uncore_io_mmio_ar_valid ),
       .io_ar_bits_addr( uncore_io_mmio_ar_bits_addr ),
       .io_ar_bits_len( uncore_io_mmio_ar_bits_len ),
       .io_ar_bits_size( uncore_io_mmio_ar_bits_size ),
       .io_ar_bits_burst( uncore_io_mmio_ar_bits_burst ),
       .io_ar_bits_lock( uncore_io_mmio_ar_bits_lock ),
       .io_ar_bits_cache( uncore_io_mmio_ar_bits_cache ),
       .io_ar_bits_prot( uncore_io_mmio_ar_bits_prot ),
       .io_ar_bits_qos( uncore_io_mmio_ar_bits_qos ),
       .io_ar_bits_region( uncore_io_mmio_ar_bits_region ),
       .io_ar_bits_id( uncore_io_mmio_ar_bits_id ),
       .io_ar_bits_user( uncore_io_mmio_ar_bits_user ),
       .io_r_ready( uncore_io_mmio_r_ready ),
       .io_r_valid( errslave_io_r_valid ),
       .io_r_bits_resp( errslave_io_r_bits_resp ),
       .io_r_bits_data( errslave_io_r_bits_data ),
       .io_r_bits_last( errslave_io_r_bits_last ),
       .io_r_bits_id( errslave_io_r_bits_id )
       //.io_r_bits_user(  )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T4(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [21:0] W0I,
  input [21:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [21:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+22) begin
    for (j=1; j<22; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [21:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][21:0] <= W0I[21:0];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [19:0] RW0M,
  input [19:0] RW0I,
  output [19:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+20) begin
    for (j=1; j<20; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [19:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][19:0] <= RW0I[19:0];
end
assign RW0O = ram[reg_RW0A];

endmodule


module ICache_T97(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


