`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module ZynqAdapter(
  input   clk,
  input   reset,
  output  io_nasti_aw_ready,
  input   io_nasti_aw_valid,
  input  [31:0] io_nasti_aw_bits_addr,
  input  [7:0] io_nasti_aw_bits_len,
  input  [2:0] io_nasti_aw_bits_size,
  input  [1:0] io_nasti_aw_bits_burst,
  input   io_nasti_aw_bits_lock,
  input  [3:0] io_nasti_aw_bits_cache,
  input  [2:0] io_nasti_aw_bits_prot,
  input  [3:0] io_nasti_aw_bits_qos,
  input  [3:0] io_nasti_aw_bits_region,
  input  [11:0] io_nasti_aw_bits_id,
  input   io_nasti_aw_bits_user,
  output  io_nasti_w_ready,
  input   io_nasti_w_valid,
  input  [31:0] io_nasti_w_bits_data,
  input   io_nasti_w_bits_last,
  input  [11:0] io_nasti_w_bits_id,
  input  [3:0] io_nasti_w_bits_strb,
  input   io_nasti_w_bits_user,
  input   io_nasti_b_ready,
  output  io_nasti_b_valid,
  output [1:0] io_nasti_b_bits_resp,
  output [11:0] io_nasti_b_bits_id,
  output  io_nasti_b_bits_user,
  output  io_nasti_ar_ready,
  input   io_nasti_ar_valid,
  input  [31:0] io_nasti_ar_bits_addr,
  input  [7:0] io_nasti_ar_bits_len,
  input  [2:0] io_nasti_ar_bits_size,
  input  [1:0] io_nasti_ar_bits_burst,
  input   io_nasti_ar_bits_lock,
  input  [3:0] io_nasti_ar_bits_cache,
  input  [2:0] io_nasti_ar_bits_prot,
  input  [3:0] io_nasti_ar_bits_qos,
  input  [3:0] io_nasti_ar_bits_region,
  input  [11:0] io_nasti_ar_bits_id,
  input   io_nasti_ar_bits_user,
  input   io_nasti_r_ready,
  output  io_nasti_r_valid,
  output [1:0] io_nasti_r_bits_resp,
  output [31:0] io_nasti_r_bits_data,
  output  io_nasti_r_bits_last,
  output [11:0] io_nasti_r_bits_id,
  output  io_nasti_r_bits_user,
  output  io_reset,
  input   io_debug_req_ready,
  output  io_debug_req_valid,
  output [4:0] io_debug_req_bits_addr,
  output [33:0] io_debug_req_bits_data,
  output [1:0] io_debug_req_bits_op,
  output  io_debug_resp_ready,
  input   io_debug_resp_valid,
  input  [33:0] io_debug_resp_bits_data,
  input  [1:0] io_debug_resp_bits_resp
);
  wire  T_371_valid;
  wire [4:0] T_371_bits_addr;
  wire [33:0] T_371_bits_data;
  wire [1:0] T_371_bits_op;
  reg  reqReg_valid;
  reg [31:0] GEN_39;
  reg [4:0] reqReg_bits_addr;
  reg [31:0] GEN_40;
  reg [33:0] reqReg_bits_data;
  reg [63:0] GEN_41;
  reg [1:0] reqReg_bits_op;
  reg [31:0] GEN_42;
  wire  T_402_valid;
  wire [33:0] T_402_bits_data;
  wire [1:0] T_402_bits_resp;
  reg  respReg_valid;
  reg [31:0] GEN_43;
  reg [33:0] respReg_bits_data;
  reg [63:0] GEN_44;
  reg [1:0] respReg_bits_resp;
  reg [31:0] GEN_45;
  wire  T_420;
  reg  awReady;
  reg [31:0] GEN_46;
  wire  GEN_0;
  wire  T_423;
  wire  T_424;
  reg  wReady;
  reg [31:0] GEN_47;
  wire  GEN_1;
  reg  arReady;
  reg [31:0] GEN_48;
  reg  rValid;
  reg [31:0] GEN_49;
  reg  bValid;
  reg [31:0] GEN_50;
  reg [11:0] bId;
  reg [31:0] GEN_51;
  wire [11:0] GEN_2;
  wire  T_429;
  reg [11:0] rId;
  reg [31:0] GEN_52;
  wire [11:0] GEN_3;
  reg [31:0] wData;
  reg [31:0] GEN_53;
  wire [31:0] GEN_4;
  wire [5:0] T_432;
  reg [5:0] wAddr;
  reg [31:0] GEN_54;
  wire [5:0] GEN_5;
  wire [5:0] T_434;
  reg [5:0] rAddr;
  reg [31:0] GEN_55;
  wire [5:0] GEN_6;
  reg  resetReg;
  reg [31:0] GEN_56;
  wire  T_437;
  wire [1:0] T_438;
  wire [3:0] T_439;
  wire [31:0] T_440;
  wire [31:0] rData;
  wire  T_443;
  wire  T_444;
  wire  T_447;
  wire  T_448;
  wire  T_449;
  wire  GEN_7;
  wire  T_451;
  wire  T_453;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_457;
  wire  T_459;
  wire  T_460;
  wire  GEN_10;
  wire  T_465;
  wire  T_466;
  wire  T_467;
  wire [4:0] T_468;
  wire [1:0] T_469;
  wire [1:0] T_470;
  wire [31:0] T_471;
  wire [33:0] T_472;
  wire [4:0] GEN_11;
  wire [1:0] GEN_12;
  wire [33:0] GEN_13;
  wire  T_474;
  wire [1:0] T_475;
  wire [33:0] T_476;
  wire [33:0] GEN_14;
  wire [4:0] GEN_15;
  wire [1:0] GEN_16;
  wire [33:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [4:0] GEN_21;
  wire [1:0] GEN_22;
  wire [33:0] GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  T_482;
  wire  T_483;
  wire  GEN_28;
  wire  T_485;
  wire  GEN_29;
  wire  T_487;
  wire  GEN_30;
  wire [33:0] GEN_31;
  wire [1:0] GEN_32;
  wire  GEN_33;
  wire [1:0] T_498_resp;
  wire [31:0] T_498_data;
  wire  T_498_last;
  wire [11:0] T_498_id;
  wire  T_498_user;
  wire [1:0] T_510_resp;
  wire [11:0] T_510_id;
  wire  T_510_user;
  wire  T_515;
  wire  T_517;
  wire [3:0] T_518;
  wire  T_520;
  wire  T_521;
  wire  T_522;
  wire  T_524;
  wire  T_526;
  wire  T_528;
  wire  T_529;
  wire  T_537;
  wire  T_538;
  wire  T_539;
  wire  T_541;
  wire  T_543;
  wire  T_545;
  wire  T_546;
  wire  T_547;
  wire  T_548;
  wire  T_549;
  wire  T_551;
  wire [4:0] GEN_34;
  reg [31:0] GEN_57;
  wire [33:0] GEN_35;
  reg [63:0] GEN_58;
  wire [1:0] GEN_36;
  reg [31:0] GEN_59;
  wire [33:0] GEN_37;
  reg [63:0] GEN_60;
  wire [1:0] GEN_38;
  reg [31:0] GEN_61;
  assign io_nasti_aw_ready = awReady;
  assign io_nasti_w_ready = wReady;
  assign io_nasti_b_valid = bValid;
  assign io_nasti_b_bits_resp = T_510_resp;
  assign io_nasti_b_bits_id = T_510_id;
  assign io_nasti_b_bits_user = T_510_user;
  assign io_nasti_ar_ready = respReg_valid;
  assign io_nasti_r_valid = rValid;
  assign io_nasti_r_bits_resp = T_498_resp;
  assign io_nasti_r_bits_data = T_498_data;
  assign io_nasti_r_bits_last = T_498_last;
  assign io_nasti_r_bits_id = T_498_id;
  assign io_nasti_r_bits_user = T_498_user;
  assign io_reset = resetReg;
  assign io_debug_req_valid = reqReg_valid;
  assign io_debug_req_bits_addr = reqReg_bits_addr;
  assign io_debug_req_bits_data = reqReg_bits_data;
  assign io_debug_req_bits_op = reqReg_bits_op;
  assign io_debug_resp_ready = T_515;
  assign T_371_valid = 1'h0;
  assign T_371_bits_addr = GEN_34;
  assign T_371_bits_data = GEN_35;
  assign T_371_bits_op = GEN_36;
  assign T_402_valid = 1'h0;
  assign T_402_bits_data = GEN_37;
  assign T_402_bits_resp = GEN_38;
  assign T_420 = io_nasti_aw_ready & io_nasti_aw_valid;
  assign GEN_0 = T_420 ? 1'h0 : awReady;
  assign T_423 = io_nasti_w_ready & io_nasti_w_valid;
  assign T_424 = T_423 & io_nasti_w_bits_last;
  assign GEN_1 = T_424 ? 1'h0 : wReady;
  assign GEN_2 = T_420 ? io_nasti_aw_bits_id : bId;
  assign T_429 = io_nasti_ar_ready & io_nasti_ar_valid;
  assign GEN_3 = T_429 ? io_nasti_ar_bits_id : rId;
  assign GEN_4 = T_424 ? io_nasti_w_bits_data : wData;
  assign T_432 = io_nasti_aw_bits_addr[5:0];
  assign GEN_5 = T_420 ? T_432 : wAddr;
  assign T_434 = io_nasti_ar_bits_addr[5:0];
  assign GEN_6 = T_429 ? T_434 : rAddr;
  assign T_437 = rAddr[2];
  assign T_438 = respReg_bits_data[33:32];
  assign T_439 = {respReg_bits_resp,T_438};
  assign T_440 = respReg_bits_data[31:0];
  assign rData = T_437 ? {{28'd0}, T_439} : T_440;
  assign T_443 = ~ io_nasti_aw_ready;
  assign T_444 = T_420 | T_443;
  assign T_447 = ~ io_nasti_w_ready;
  assign T_448 = T_424 | T_447;
  assign T_449 = T_444 & T_448;
  assign GEN_7 = T_449 ? 1'h1 : bValid;
  assign T_451 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_453 = wAddr == 6'h8;
  assign GEN_8 = T_453 ? 1'h1 : reqReg_valid;
  assign GEN_9 = T_453 ? 1'h0 : respReg_valid;
  assign T_457 = wAddr == 6'h20;
  assign T_459 = T_453 == 1'h0;
  assign T_460 = T_459 & T_457;
  assign GEN_10 = T_460 ? 1'h1 : resetReg;
  assign T_465 = T_457 == 1'h0;
  assign T_466 = T_459 & T_465;
  assign T_467 = wAddr[2];
  assign T_468 = wData[8:4];
  assign T_469 = wData[3:2];
  assign T_470 = wData[1:0];
  assign T_471 = reqReg_bits_data[31:0];
  assign T_472 = {T_470,T_471};
  assign GEN_11 = T_467 ? T_468 : reqReg_bits_addr;
  assign GEN_12 = T_467 ? T_469 : reqReg_bits_op;
  assign GEN_13 = T_467 ? T_472 : reqReg_bits_data;
  assign T_474 = T_467 == 1'h0;
  assign T_475 = reqReg_bits_data[33:32];
  assign T_476 = {T_475,wData};
  assign GEN_14 = T_474 ? T_476 : GEN_13;
  assign GEN_15 = T_466 ? GEN_11 : reqReg_bits_addr;
  assign GEN_16 = T_466 ? GEN_12 : reqReg_bits_op;
  assign GEN_17 = T_466 ? GEN_14 : reqReg_bits_data;
  assign GEN_18 = T_451 ? GEN_8 : reqReg_valid;
  assign GEN_19 = T_451 ? GEN_9 : respReg_valid;
  assign GEN_20 = T_451 ? GEN_10 : resetReg;
  assign GEN_21 = T_451 ? GEN_15 : reqReg_bits_addr;
  assign GEN_22 = T_451 ? GEN_16 : reqReg_bits_op;
  assign GEN_23 = T_451 ? GEN_17 : reqReg_bits_data;
  assign GEN_24 = T_451 ? 1'h1 : GEN_0;
  assign GEN_25 = T_451 ? 1'h1 : GEN_1;
  assign GEN_26 = T_451 ? 1'h0 : GEN_7;
  assign GEN_27 = T_429 ? 1'h1 : rValid;
  assign T_482 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_483 = T_482 & io_nasti_r_bits_last;
  assign GEN_28 = T_483 ? 1'h0 : GEN_27;
  assign T_485 = io_debug_req_ready & io_debug_req_valid;
  assign GEN_29 = T_485 ? 1'h0 : GEN_18;
  assign T_487 = io_debug_resp_ready & io_debug_resp_valid;
  assign GEN_30 = T_487 ? 1'h1 : GEN_19;
  assign GEN_31 = T_487 ? io_debug_resp_bits_data : respReg_bits_data;
  assign GEN_32 = T_487 ? io_debug_resp_bits_resp : respReg_bits_resp;
  assign GEN_33 = resetReg ? 1'h0 : GEN_20;
  assign T_498_resp = 2'h0;
  assign T_498_data = rData;
  assign T_498_last = 1'h1;
  assign T_498_id = rId;
  assign T_498_user = 1'h0;
  assign T_510_resp = 2'h0;
  assign T_510_id = bId;
  assign T_510_user = 1'h0;
  assign T_515 = ~ respReg_valid;
  assign T_517 = io_nasti_w_valid == 1'h0;
  assign T_518 = ~ io_nasti_w_bits_strb;
  assign T_520 = T_518 == 4'h0;
  assign T_521 = T_517 | T_520;
  assign T_522 = T_521 | reset;
  assign T_524 = T_522 == 1'h0;
  assign T_526 = io_nasti_ar_valid == 1'h0;
  assign T_528 = io_nasti_ar_bits_len == 8'h0;
  assign T_529 = T_526 | T_528;
  assign T_537 = io_nasti_ar_bits_burst == 2'h0;
  assign T_538 = T_529 | T_537;
  assign T_539 = T_538 | reset;
  assign T_541 = T_539 == 1'h0;
  assign T_543 = io_nasti_aw_valid == 1'h0;
  assign T_545 = io_nasti_aw_bits_len == 8'h0;
  assign T_546 = T_543 | T_545;
  assign T_547 = io_nasti_aw_bits_burst == 2'h0;
  assign T_548 = T_546 | T_547;
  assign T_549 = T_548 | reset;
  assign T_551 = T_549 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_57[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_58[33:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_59[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_60[33:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_61[1:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  reqReg_valid = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  reqReg_bits_addr = GEN_40[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {2{$random}};
  reqReg_bits_data = GEN_41[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  reqReg_bits_op = GEN_42[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  respReg_valid = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {2{$random}};
  respReg_bits_data = GEN_44[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  respReg_bits_resp = GEN_45[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  awReady = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  wReady = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  arReady = GEN_48[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  rValid = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  bValid = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  bId = GEN_51[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  rId = GEN_52[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  wData = GEN_53[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  wAddr = GEN_54[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  rAddr = GEN_55[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  resetReg = GEN_56[0:0];
  `endif
  GEN_57 = {1{$random}};
  GEN_58 = {2{$random}};
  GEN_59 = {1{$random}};
  GEN_60 = {2{$random}};
  GEN_61 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reqReg_valid <= T_371_valid;
    end else begin
      if(T_485) begin
        reqReg_valid <= 1'h0;
      end else begin
        if(T_451) begin
          if(T_453) begin
            reqReg_valid <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_addr <= T_371_bits_addr;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_467) begin
            reqReg_bits_addr <= T_468;
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_data <= T_371_bits_data;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_474) begin
            reqReg_bits_data <= T_476;
          end else begin
            if(T_467) begin
              reqReg_bits_data <= T_472;
            end
          end
        end
      end
    end
    if(reset) begin
      reqReg_bits_op <= T_371_bits_op;
    end else begin
      if(T_451) begin
        if(T_466) begin
          if(T_467) begin
            reqReg_bits_op <= T_469;
          end
        end
      end
    end
    if(reset) begin
      respReg_valid <= T_402_valid;
    end else begin
      if(T_487) begin
        respReg_valid <= 1'h1;
      end else begin
        if(T_451) begin
          if(T_453) begin
            respReg_valid <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      respReg_bits_data <= T_402_bits_data;
    end else begin
      if(T_487) begin
        respReg_bits_data <= io_debug_resp_bits_data;
      end
    end
    if(reset) begin
      respReg_bits_resp <= T_402_bits_resp;
    end else begin
      if(T_487) begin
        respReg_bits_resp <= io_debug_resp_bits_resp;
      end
    end
    if(reset) begin
      awReady <= 1'h1;
    end else begin
      if(T_451) begin
        awReady <= 1'h1;
      end else begin
        if(T_420) begin
          awReady <= 1'h0;
        end
      end
    end
    if(reset) begin
      wReady <= 1'h1;
    end else begin
      if(T_451) begin
        wReady <= 1'h1;
      end else begin
        if(T_424) begin
          wReady <= 1'h0;
        end
      end
    end
    if(reset) begin
      arReady <= 1'h0;
    end
    if(reset) begin
      rValid <= 1'h0;
    end else begin
      if(T_483) begin
        rValid <= 1'h0;
      end else begin
        if(T_429) begin
          rValid <= 1'h1;
        end
      end
    end
    if(reset) begin
      bValid <= 1'h0;
    end else begin
      if(T_451) begin
        bValid <= 1'h0;
      end else begin
        if(T_449) begin
          bValid <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_420) begin
        bId <= io_nasti_aw_bits_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_429) begin
        rId <= io_nasti_ar_bits_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_424) begin
        wData <= io_nasti_w_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_420) begin
        wAddr <= T_432;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_429) begin
        rAddr <= T_434;
      end
    end
    if(reset) begin
      resetReg <= 1'h0;
    end else begin
      if(resetReg) begin
        resetReg <= 1'h0;
      end else begin
        if(T_451) begin
          if(T_460) begin
            resetReg <= 1'h1;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_524) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter cannot take partial writes\n    at Adapter.scala:129 assert(!w.valid || w.bits.strb.andR,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_524) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_541) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter can only take fixed bursts\n    at Adapter.scala:131 assert(!ar.valid ||\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_541) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_551) begin
          $fwrite(32'h80000002,"Assertion failed: Nasti to DebugBusIO converter can only take fixed bursts\n    at Adapter.scala:135 assert(!aw.valid ||\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_551) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module RVCExpander(
  input   clk,
  input   reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0] io_out_rd,
  output [4:0] io_out_rs1,
  output [4:0] io_out_rs2,
  output [4:0] io_out_rs3,
  output  io_rvc
);
  wire [1:0] T_8;
  wire  T_10;
  wire [7:0] T_11;
  wire  T_13;
  wire [6:0] T_16;
  wire [3:0] T_17;
  wire [1:0] T_18;
  wire  T_19;
  wire  T_20;
  wire [2:0] T_22;
  wire [5:0] T_23;
  wire [6:0] T_24;
  wire [9:0] T_25;
  wire [2:0] T_29;
  wire [4:0] T_30;
  wire [11:0] T_31;
  wire [14:0] T_32;
  wire [17:0] T_33;
  wire [29:0] T_34;
  wire [4:0] T_42;
  wire [31:0] T_49_bits;
  wire [4:0] T_49_rd;
  wire [4:0] T_49_rs1;
  wire [4:0] T_49_rs2;
  wire [4:0] T_49_rs3;
  wire [1:0] T_55;
  wire [2:0] T_56;
  wire [4:0] T_58;
  wire [7:0] T_59;
  wire [2:0] T_61;
  wire [4:0] T_62;
  wire [11:0] T_68;
  wire [12:0] T_69;
  wire [15:0] T_70;
  wire [27:0] T_71;
  wire [31:0] T_88_bits;
  wire [4:0] T_88_rd;
  wire [4:0] T_88_rs1;
  wire [4:0] T_88_rs2;
  wire [4:0] T_88_rs3;
  wire [3:0] T_99;
  wire [6:0] T_100;
  wire [11:0] T_109;
  wire [11:0] T_110;
  wire [14:0] T_111;
  wire [26:0] T_112;
  wire [31:0] T_129_bits;
  wire [4:0] T_129_rd;
  wire [4:0] T_129_rs1;
  wire [4:0] T_129_rs2;
  wire [4:0] T_129_rs3;
  wire [27:0] T_151;
  wire [31:0] T_168_bits;
  wire [4:0] T_168_rd;
  wire [4:0] T_168_rs1;
  wire [4:0] T_168_rs2;
  wire [4:0] T_168_rs3;
  wire [1:0] T_181;
  wire [4:0] T_196;
  wire [7:0] T_198;
  wire [14:0] T_199;
  wire [6:0] T_200;
  wire [11:0] T_201;
  wire [26:0] T_202;
  wire [31:0] T_219_bits;
  wire [4:0] T_219_rd;
  wire [4:0] T_219_rs1;
  wire [4:0] T_219_rs2;
  wire [4:0] T_219_rs3;
  wire [2:0] T_230;
  wire [4:0] T_243;
  wire [7:0] T_245;
  wire [14:0] T_246;
  wire [7:0] T_247;
  wire [12:0] T_248;
  wire [27:0] T_249;
  wire [31:0] T_266_bits;
  wire [4:0] T_266_rd;
  wire [4:0] T_266_rs1;
  wire [4:0] T_266_rs2;
  wire [4:0] T_266_rs3;
  wire [14:0] T_297;
  wire [26:0] T_300;
  wire [31:0] T_317_bits;
  wire [4:0] T_317_rd;
  wire [4:0] T_317_rs1;
  wire [4:0] T_317_rs2;
  wire [4:0] T_317_rs3;
  wire [14:0] T_344;
  wire [27:0] T_347;
  wire [31:0] T_364_bits;
  wire [4:0] T_364_rd;
  wire [4:0] T_364_rs1;
  wire [4:0] T_364_rs2;
  wire [4:0] T_364_rs3;
  wire  T_370;
  wire [6:0] T_374;
  wire [4:0] T_375;
  wire [11:0] T_376;
  wire [4:0] T_377;
  wire [11:0] T_381;
  wire [16:0] T_382;
  wire [19:0] T_383;
  wire [31:0] T_384;
  wire [31:0] T_397_bits;
  wire [4:0] T_397_rd;
  wire [4:0] T_397_rs1;
  wire [4:0] T_397_rs2;
  wire [4:0] T_397_rs3;
  wire  T_405;
  wire [6:0] T_408;
  wire [11:0] T_419;
  wire [31:0] T_422;
  wire [31:0] T_435_bits;
  wire [4:0] T_435_rd;
  wire [4:0] T_435_rs1;
  wire [4:0] T_435_rs2;
  wire [4:0] T_435_rs3;
  wire [16:0] T_453;
  wire [19:0] T_454;
  wire [31:0] T_455;
  wire [31:0] T_468_bits;
  wire [4:0] T_468_rd;
  wire [4:0] T_468_rs1;
  wire [4:0] T_468_rs2;
  wire [4:0] T_468_rs3;
  wire  T_482;
  wire [6:0] T_485;
  wire [14:0] T_490;
  wire [19:0] T_493;
  wire [31:0] T_494;
  wire [19:0] T_495;
  wire [24:0] T_497;
  wire [31:0] T_498;
  wire [31:0] T_511_bits;
  wire [4:0] T_511_rd;
  wire [4:0] T_511_rs1;
  wire [4:0] T_511_rs2;
  wire [4:0] T_511_rs3;
  wire  T_519;
  wire  T_522;
  wire  T_523;
  wire [6:0] T_535;
  wire [2:0] T_540;
  wire [1:0] T_541;
  wire  T_543;
  wire [1:0] T_546;
  wire [5:0] T_547;
  wire [4:0] T_548;
  wire [5:0] T_549;
  wire [11:0] T_550;
  wire [11:0] T_554;
  wire [16:0] T_555;
  wire [19:0] T_556;
  wire [31:0] T_557;
  wire [31:0] T_570_bits;
  wire [4:0] T_570_rd;
  wire [4:0] T_570_rs1;
  wire [4:0] T_570_rs2;
  wire [4:0] T_570_rs3;
  wire [31:0] T_576_bits;
  wire [4:0] T_576_rd;
  wire [4:0] T_576_rs1;
  wire [4:0] T_576_rs2;
  wire [4:0] T_576_rs3;
  wire [5:0] T_584;
  wire [11:0] T_593;
  wire [10:0] T_594;
  wire [13:0] T_595;
  wire [25:0] T_596;
  wire [30:0] GEN_0;
  wire [30:0] T_613;
  wire [16:0] T_630;
  wire [19:0] T_631;
  wire [31:0] T_632;
  wire [2:0] T_643;
  wire [2:0] T_645;
  wire  T_647;
  wire [2:0] T_649;
  wire  T_651;
  wire  T_655;
  wire [1:0] T_656;
  wire [1:0] T_662;
  wire [2:0] T_671;
  wire [2:0] T_676;
  wire [2:0] T_677;
  wire [2:0] T_678;
  wire  T_681;
  wire [30:0] T_684;
  wire [6:0] T_688;
  wire [11:0] T_698;
  wire [9:0] T_699;
  wire [12:0] T_700;
  wire [24:0] T_701;
  wire [30:0] GEN_1;
  wire [30:0] T_702;
  wire [1:0] T_703;
  wire [1:0] T_705;
  wire  T_707;
  wire  T_711;
  wire [31:0] T_712;
  wire [30:0] T_717;
  wire [31:0] T_718;
  wire [31:0] T_735_bits;
  wire [4:0] T_735_rd;
  wire [4:0] T_735_rs1;
  wire [4:0] T_735_rs2;
  wire [4:0] T_735_rs3;
  wire [9:0] T_745;
  wire  T_746;
  wire [1:0] T_747;
  wire  T_749;
  wire  T_751;
  wire [2:0] T_752;
  wire [3:0] T_754;
  wire [1:0] T_755;
  wire [5:0] T_756;
  wire [1:0] T_757;
  wire [10:0] T_758;
  wire [12:0] T_759;
  wire [14:0] T_760;
  wire [20:0] T_761;
  wire  T_762;
  wire [9:0] T_784;
  wire  T_806;
  wire [7:0] T_828;
  wire [12:0] T_831;
  wire [19:0] T_832;
  wire [10:0] T_833;
  wire [11:0] T_834;
  wire [31:0] T_835;
  wire [31:0] T_850_bits;
  wire [4:0] T_850_rd;
  wire [4:0] T_850_rs1;
  wire [4:0] T_850_rs2;
  wire [4:0] T_850_rs3;
  wire [4:0] T_860;
  wire [3:0] T_866;
  wire [4:0] T_867;
  wire [6:0] T_868;
  wire [7:0] T_869;
  wire [12:0] T_870;
  wire  T_871;
  wire [5:0] T_887;
  wire [3:0] T_908;
  wire  T_924;
  wire [7:0] T_926;
  wire [6:0] T_927;
  wire [14:0] T_928;
  wire [9:0] T_929;
  wire [6:0] T_930;
  wire [16:0] T_931;
  wire [31:0] T_932;
  wire [31:0] T_947_bits;
  wire [4:0] T_947_rd;
  wire [4:0] T_947_rs1;
  wire [4:0] T_947_rs2;
  wire [4:0] T_947_rs3;
  wire [6:0] T_1024;
  wire [14:0] T_1025;
  wire [31:0] T_1029;
  wire [31:0] T_1042_bits;
  wire [4:0] T_1042_rd;
  wire [4:0] T_1042_rs1;
  wire [4:0] T_1042_rs2;
  wire [4:0] T_1042_rs3;
  wire [10:0] T_1056;
  wire [13:0] T_1057;
  wire [25:0] T_1058;
  wire [31:0] T_1069_bits;
  wire [4:0] T_1069_rd;
  wire [4:0] T_1069_rs1;
  wire [4:0] T_1069_rs2;
  wire [4:0] T_1069_rs3;
  wire [4:0] T_1079;
  wire [3:0] T_1080;
  wire [8:0] T_1081;
  wire [11:0] T_1086;
  wire [13:0] T_1087;
  wire [16:0] T_1088;
  wire [28:0] T_1089;
  wire [31:0] T_1100_bits;
  wire [4:0] T_1100_rd;
  wire [4:0] T_1100_rs1;
  wire [4:0] T_1100_rs2;
  wire [4:0] T_1100_rs3;
  wire [1:0] T_1106;
  wire [2:0] T_1108;
  wire [4:0] T_1110;
  wire [2:0] T_1111;
  wire [7:0] T_1112;
  wire [11:0] T_1117;
  wire [12:0] T_1118;
  wire [15:0] T_1119;
  wire [27:0] T_1120;
  wire [31:0] T_1131_bits;
  wire [4:0] T_1131_rd;
  wire [4:0] T_1131_rs1;
  wire [4:0] T_1131_rs2;
  wire [4:0] T_1131_rs3;
  wire [28:0] T_1151;
  wire [31:0] T_1162_bits;
  wire [4:0] T_1162_rd;
  wire [4:0] T_1162_rs1;
  wire [4:0] T_1162_rs2;
  wire [4:0] T_1162_rs3;
  wire [11:0] T_1173;
  wire [9:0] T_1174;
  wire [12:0] T_1175;
  wire [24:0] T_1176;
  wire [31:0] T_1187_bits;
  wire [4:0] T_1187_rd;
  wire [4:0] T_1187_rs1;
  wire [4:0] T_1187_rs2;
  wire [4:0] T_1187_rs3;
  wire [9:0] T_1199;
  wire [12:0] T_1200;
  wire [24:0] T_1201;
  wire [31:0] T_1212_bits;
  wire [4:0] T_1212_rd;
  wire [4:0] T_1212_rs1;
  wire [4:0] T_1212_rs2;
  wire [4:0] T_1212_rs3;
  wire [24:0] T_1226;
  wire [17:0] T_1227;
  wire [24:0] T_1229;
  wire [24:0] T_1233;
  wire [31:0] T_1244_bits;
  wire [4:0] T_1244_rd;
  wire [4:0] T_1244_rs1;
  wire [4:0] T_1244_rs2;
  wire [4:0] T_1244_rs3;
  wire  T_1252;
  wire [31:0] T_1253_bits;
  wire [4:0] T_1253_rd;
  wire [4:0] T_1253_rs1;
  wire [4:0] T_1253_rs2;
  wire [4:0] T_1253_rs3;
  wire [24:0] T_1267;
  wire [24:0] T_1270;
  wire [24:0] T_1272;
  wire [24:0] T_1276;
  wire [31:0] T_1287_bits;
  wire [4:0] T_1287_rd;
  wire [4:0] T_1287_rs1;
  wire [4:0] T_1287_rs2;
  wire [4:0] T_1287_rs3;
  wire [31:0] T_1296_bits;
  wire [4:0] T_1296_rd;
  wire [4:0] T_1296_rs1;
  wire [4:0] T_1296_rs2;
  wire [4:0] T_1296_rs3;
  wire [31:0] T_1303_bits;
  wire [4:0] T_1303_rd;
  wire [4:0] T_1303_rs1;
  wire [4:0] T_1303_rs2;
  wire [4:0] T_1303_rs3;
  wire [5:0] T_1312;
  wire [8:0] T_1313;
  wire [3:0] T_1314;
  wire [4:0] T_1323;
  wire [7:0] T_1325;
  wire [14:0] T_1326;
  wire [8:0] T_1327;
  wire [13:0] T_1328;
  wire [28:0] T_1329;
  wire [31:0] T_1340_bits;
  wire [4:0] T_1340_rd;
  wire [4:0] T_1340_rs1;
  wire [4:0] T_1340_rs2;
  wire [4:0] T_1340_rs3;
  wire [1:0] T_1346;
  wire [3:0] T_1347;
  wire [5:0] T_1349;
  wire [7:0] T_1350;
  wire [2:0] T_1351;
  wire [4:0] T_1360;
  wire [7:0] T_1362;
  wire [14:0] T_1363;
  wire [7:0] T_1364;
  wire [12:0] T_1365;
  wire [27:0] T_1366;
  wire [31:0] T_1377_bits;
  wire [4:0] T_1377_rd;
  wire [4:0] T_1377_rs1;
  wire [4:0] T_1377_rs2;
  wire [4:0] T_1377_rs3;
  wire [14:0] T_1400;
  wire [28:0] T_1403;
  wire [31:0] T_1414_bits;
  wire [4:0] T_1414_rd;
  wire [4:0] T_1414_rs1;
  wire [4:0] T_1414_rs2;
  wire [4:0] T_1414_rs3;
  wire [4:0] T_1421;
  wire [4:0] T_1422;
  wire [31:0] T_1430_bits;
  wire [4:0] T_1430_rd;
  wire [4:0] T_1430_rs1;
  wire [4:0] T_1430_rs2;
  wire [4:0] T_1430_rs3;
  wire [31:0] T_1446_bits;
  wire [4:0] T_1446_rd;
  wire [4:0] T_1446_rs1;
  wire [4:0] T_1446_rs2;
  wire [4:0] T_1446_rs3;
  wire [31:0] T_1462_bits;
  wire [4:0] T_1462_rd;
  wire [4:0] T_1462_rs1;
  wire [4:0] T_1462_rs2;
  wire [4:0] T_1462_rs3;
  wire [31:0] T_1478_bits;
  wire [4:0] T_1478_rd;
  wire [4:0] T_1478_rs1;
  wire [4:0] T_1478_rs2;
  wire [4:0] T_1478_rs3;
  wire [31:0] T_1494_bits;
  wire [4:0] T_1494_rd;
  wire [4:0] T_1494_rs1;
  wire [4:0] T_1494_rs2;
  wire [4:0] T_1494_rs3;
  wire [31:0] T_1510_bits;
  wire [4:0] T_1510_rd;
  wire [4:0] T_1510_rs1;
  wire [4:0] T_1510_rs2;
  wire [4:0] T_1510_rs3;
  wire [31:0] T_1526_bits;
  wire [4:0] T_1526_rd;
  wire [4:0] T_1526_rs1;
  wire [4:0] T_1526_rs2;
  wire [4:0] T_1526_rs3;
  wire [31:0] T_1542_bits;
  wire [4:0] T_1542_rd;
  wire [4:0] T_1542_rs1;
  wire [4:0] T_1542_rs2;
  wire [4:0] T_1542_rs3;
  wire [2:0] T_1549;
  wire [4:0] T_1550;
  wire [4:0] T_1552;
  wire  T_1554;
  wire [4:0] T_1556;
  wire  T_1558;
  wire [4:0] T_1560;
  wire  T_1562;
  wire [4:0] T_1564;
  wire  T_1566;
  wire  T_1570;
  wire [31:0] T_1571_bits;
  wire [4:0] T_1571_rd;
  wire [4:0] T_1571_rs1;
  wire [4:0] T_1571_rs2;
  wire [4:0] T_1571_rs3;
  wire [31:0] T_1581_bits;
  wire [4:0] T_1581_rd;
  wire [4:0] T_1581_rs1;
  wire [4:0] T_1581_rs2;
  wire [4:0] T_1581_rs3;
  wire [31:0] T_1587_bits;
  wire [4:0] T_1587_rd;
  wire [4:0] T_1587_rs1;
  wire [4:0] T_1587_rs2;
  wire [4:0] T_1587_rs3;
  wire [31:0] T_1601_bits;
  wire [4:0] T_1601_rd;
  wire [4:0] T_1601_rs1;
  wire [4:0] T_1601_rs2;
  wire [4:0] T_1601_rs3;
  wire [31:0] T_1611_bits;
  wire [4:0] T_1611_rd;
  wire [4:0] T_1611_rs1;
  wire [4:0] T_1611_rs2;
  wire [4:0] T_1611_rs3;
  wire [31:0] T_1617_bits;
  wire [4:0] T_1617_rd;
  wire [4:0] T_1617_rs1;
  wire [4:0] T_1617_rs2;
  wire [4:0] T_1617_rs3;
  wire [31:0] T_1623_bits;
  wire [4:0] T_1623_rd;
  wire [4:0] T_1623_rs1;
  wire [4:0] T_1623_rs2;
  wire [4:0] T_1623_rs3;
  wire [31:0] T_1641_bits;
  wire [4:0] T_1641_rd;
  wire [4:0] T_1641_rs1;
  wire [4:0] T_1641_rs2;
  wire [4:0] T_1641_rs3;
  wire [31:0] T_1651_bits;
  wire [4:0] T_1651_rd;
  wire [4:0] T_1651_rs1;
  wire [4:0] T_1651_rs2;
  wire [4:0] T_1651_rs3;
  wire [31:0] T_1657_bits;
  wire [4:0] T_1657_rd;
  wire [4:0] T_1657_rs1;
  wire [4:0] T_1657_rs2;
  wire [4:0] T_1657_rs3;
  wire [31:0] T_1671_bits;
  wire [4:0] T_1671_rd;
  wire [4:0] T_1671_rs1;
  wire [4:0] T_1671_rs2;
  wire [4:0] T_1671_rs3;
  wire [31:0] T_1681_bits;
  wire [4:0] T_1681_rd;
  wire [4:0] T_1681_rs1;
  wire [4:0] T_1681_rs2;
  wire [4:0] T_1681_rs3;
  wire [31:0] T_1687_bits;
  wire [4:0] T_1687_rd;
  wire [4:0] T_1687_rs1;
  wire [4:0] T_1687_rs2;
  wire [4:0] T_1687_rs3;
  wire [31:0] T_1693_bits;
  wire [4:0] T_1693_rd;
  wire [4:0] T_1693_rs1;
  wire [4:0] T_1693_rs2;
  wire [4:0] T_1693_rs3;
  wire [31:0] T_1699_bits;
  wire [4:0] T_1699_rd;
  wire [4:0] T_1699_rs1;
  wire [4:0] T_1699_rs2;
  wire [4:0] T_1699_rs3;
  wire [31:0] T_1721_bits;
  wire [4:0] T_1721_rd;
  wire [4:0] T_1721_rs1;
  wire [4:0] T_1721_rs2;
  wire [4:0] T_1721_rs3;
  wire [31:0] T_1731_bits;
  wire [4:0] T_1731_rd;
  wire [4:0] T_1731_rs1;
  wire [4:0] T_1731_rs2;
  wire [4:0] T_1731_rs3;
  wire [31:0] T_1737_bits;
  wire [4:0] T_1737_rd;
  wire [4:0] T_1737_rs1;
  wire [4:0] T_1737_rs2;
  wire [4:0] T_1737_rs3;
  wire [31:0] T_1751_bits;
  wire [4:0] T_1751_rd;
  wire [4:0] T_1751_rs1;
  wire [4:0] T_1751_rs2;
  wire [4:0] T_1751_rs3;
  wire [31:0] T_1761_bits;
  wire [4:0] T_1761_rd;
  wire [4:0] T_1761_rs1;
  wire [4:0] T_1761_rs2;
  wire [4:0] T_1761_rs3;
  wire [31:0] T_1767_bits;
  wire [4:0] T_1767_rd;
  wire [4:0] T_1767_rs1;
  wire [4:0] T_1767_rs2;
  wire [4:0] T_1767_rs3;
  wire [31:0] T_1773_bits;
  wire [4:0] T_1773_rd;
  wire [4:0] T_1773_rs1;
  wire [4:0] T_1773_rs2;
  wire [4:0] T_1773_rs3;
  wire [31:0] T_1791_bits;
  wire [4:0] T_1791_rd;
  wire [4:0] T_1791_rs1;
  wire [4:0] T_1791_rs2;
  wire [4:0] T_1791_rs3;
  wire [31:0] T_1801_bits;
  wire [4:0] T_1801_rd;
  wire [4:0] T_1801_rs1;
  wire [4:0] T_1801_rs2;
  wire [4:0] T_1801_rs3;
  wire [31:0] T_1807_bits;
  wire [4:0] T_1807_rd;
  wire [4:0] T_1807_rs1;
  wire [4:0] T_1807_rs2;
  wire [4:0] T_1807_rs3;
  wire [31:0] T_1821_bits;
  wire [4:0] T_1821_rd;
  wire [4:0] T_1821_rs1;
  wire [4:0] T_1821_rs2;
  wire [4:0] T_1821_rs3;
  wire [31:0] T_1831_bits;
  wire [4:0] T_1831_rd;
  wire [4:0] T_1831_rs1;
  wire [4:0] T_1831_rs2;
  wire [4:0] T_1831_rs3;
  wire [31:0] T_1837_bits;
  wire [4:0] T_1837_rd;
  wire [4:0] T_1837_rs1;
  wire [4:0] T_1837_rs2;
  wire [4:0] T_1837_rs3;
  wire [31:0] T_1843_bits;
  wire [4:0] T_1843_rd;
  wire [4:0] T_1843_rs1;
  wire [4:0] T_1843_rs2;
  wire [4:0] T_1843_rs3;
  wire [31:0] T_1849_bits;
  wire [4:0] T_1849_rd;
  wire [4:0] T_1849_rs1;
  wire [4:0] T_1849_rs2;
  wire [4:0] T_1849_rs3;
  wire [31:0] T_1855_bits;
  wire [4:0] T_1855_rd;
  wire [4:0] T_1855_rs1;
  wire [4:0] T_1855_rs2;
  wire [4:0] T_1855_rs3;
  assign io_out_bits = T_1855_bits;
  assign io_out_rd = T_1855_rd;
  assign io_out_rs1 = T_1855_rs1;
  assign io_out_rs2 = T_1855_rs2;
  assign io_out_rs3 = T_1855_rs3;
  assign io_rvc = T_10;
  assign T_8 = io_in[1:0];
  assign T_10 = T_8 != 2'h3;
  assign T_11 = io_in[12:5];
  assign T_13 = T_11 != 8'h0;
  assign T_16 = T_13 ? 7'h13 : 7'h1f;
  assign T_17 = io_in[10:7];
  assign T_18 = io_in[12:11];
  assign T_19 = io_in[5];
  assign T_20 = io_in[6];
  assign T_22 = {T_20,2'h0};
  assign T_23 = {T_17,T_18};
  assign T_24 = {T_23,T_19};
  assign T_25 = {T_24,T_22};
  assign T_29 = io_in[4:2];
  assign T_30 = {2'h1,T_29};
  assign T_31 = {T_30,T_16};
  assign T_32 = {T_25,5'h2};
  assign T_33 = {T_32,3'h0};
  assign T_34 = {T_33,T_31};
  assign T_42 = io_in[31:27];
  assign T_49_bits = {{2'd0}, T_34};
  assign T_49_rd = T_30;
  assign T_49_rs1 = 5'h2;
  assign T_49_rs2 = T_30;
  assign T_49_rs3 = T_42;
  assign T_55 = io_in[6:5];
  assign T_56 = io_in[12:10];
  assign T_58 = {T_55,T_56};
  assign T_59 = {T_58,3'h0};
  assign T_61 = io_in[9:7];
  assign T_62 = {2'h1,T_61};
  assign T_68 = {T_30,7'h7};
  assign T_69 = {T_59,T_62};
  assign T_70 = {T_69,3'h3};
  assign T_71 = {T_70,T_68};
  assign T_88_bits = {{4'd0}, T_71};
  assign T_88_rd = T_30;
  assign T_88_rs1 = T_62;
  assign T_88_rs2 = T_30;
  assign T_88_rs3 = T_42;
  assign T_99 = {T_19,T_56};
  assign T_100 = {T_99,T_22};
  assign T_109 = {T_30,7'h3};
  assign T_110 = {T_100,T_62};
  assign T_111 = {T_110,3'h2};
  assign T_112 = {T_111,T_109};
  assign T_129_bits = {{5'd0}, T_112};
  assign T_129_rd = T_30;
  assign T_129_rs1 = T_62;
  assign T_129_rs2 = T_30;
  assign T_129_rs3 = T_42;
  assign T_151 = {T_70,T_109};
  assign T_168_bits = {{4'd0}, T_151};
  assign T_168_rd = T_30;
  assign T_168_rs1 = T_62;
  assign T_168_rs2 = T_30;
  assign T_168_rs3 = T_42;
  assign T_181 = T_100[6:5];
  assign T_196 = T_100[4:0];
  assign T_198 = {3'h2,T_196};
  assign T_199 = {T_198,7'h2f};
  assign T_200 = {T_181,T_30};
  assign T_201 = {T_200,T_62};
  assign T_202 = {T_201,T_199};
  assign T_219_bits = {{5'd0}, T_202};
  assign T_219_rd = T_30;
  assign T_219_rs1 = T_62;
  assign T_219_rs2 = T_30;
  assign T_219_rs3 = T_42;
  assign T_230 = T_59[7:5];
  assign T_243 = T_59[4:0];
  assign T_245 = {3'h3,T_243};
  assign T_246 = {T_245,7'h27};
  assign T_247 = {T_230,T_30};
  assign T_248 = {T_247,T_62};
  assign T_249 = {T_248,T_246};
  assign T_266_bits = {{4'd0}, T_249};
  assign T_266_rd = T_30;
  assign T_266_rs1 = T_62;
  assign T_266_rs2 = T_30;
  assign T_266_rs3 = T_42;
  assign T_297 = {T_198,7'h23};
  assign T_300 = {T_201,T_297};
  assign T_317_bits = {{5'd0}, T_300};
  assign T_317_rd = T_30;
  assign T_317_rs1 = T_62;
  assign T_317_rs2 = T_30;
  assign T_317_rs3 = T_42;
  assign T_344 = {T_245,7'h23};
  assign T_347 = {T_248,T_344};
  assign T_364_bits = {{4'd0}, T_347};
  assign T_364_rd = T_30;
  assign T_364_rs1 = T_62;
  assign T_364_rs2 = T_30;
  assign T_364_rs3 = T_42;
  assign T_370 = io_in[12];
  assign T_374 = T_370 ? 7'h7f : 7'h0;
  assign T_375 = io_in[6:2];
  assign T_376 = {T_374,T_375};
  assign T_377 = io_in[11:7];
  assign T_381 = {T_377,7'h13};
  assign T_382 = {T_376,T_377};
  assign T_383 = {T_382,3'h0};
  assign T_384 = {T_383,T_381};
  assign T_397_bits = T_384;
  assign T_397_rd = T_377;
  assign T_397_rs1 = T_377;
  assign T_397_rs2 = T_30;
  assign T_397_rs3 = T_42;
  assign T_405 = T_377 != 5'h0;
  assign T_408 = T_405 ? 7'h1b : 7'h1f;
  assign T_419 = {T_377,T_408};
  assign T_422 = {T_383,T_419};
  assign T_435_bits = T_422;
  assign T_435_rd = T_377;
  assign T_435_rs1 = T_377;
  assign T_435_rs2 = T_30;
  assign T_435_rs3 = T_42;
  assign T_453 = {T_376,5'h0};
  assign T_454 = {T_453,3'h0};
  assign T_455 = {T_454,T_381};
  assign T_468_bits = T_455;
  assign T_468_rd = T_377;
  assign T_468_rs1 = 5'h0;
  assign T_468_rs2 = T_30;
  assign T_468_rs3 = T_42;
  assign T_482 = T_376 != 12'h0;
  assign T_485 = T_482 ? 7'h37 : 7'h3f;
  assign T_490 = T_370 ? 15'h7fff : 15'h0;
  assign T_493 = {T_490,T_375};
  assign T_494 = {T_493,12'h0};
  assign T_495 = T_494[31:12];
  assign T_497 = {T_495,T_377};
  assign T_498 = {T_497,T_485};
  assign T_511_bits = T_498;
  assign T_511_rd = T_377;
  assign T_511_rs1 = T_377;
  assign T_511_rs2 = T_30;
  assign T_511_rs3 = T_42;
  assign T_519 = T_377 == 5'h0;
  assign T_522 = T_377 == 5'h2;
  assign T_523 = T_519 | T_522;
  assign T_535 = T_482 ? 7'h13 : 7'h1f;
  assign T_540 = T_370 ? 3'h7 : 3'h0;
  assign T_541 = io_in[4:3];
  assign T_543 = io_in[2];
  assign T_546 = {T_543,T_20};
  assign T_547 = {T_546,4'h0};
  assign T_548 = {T_540,T_541};
  assign T_549 = {T_548,T_19};
  assign T_550 = {T_549,T_547};
  assign T_554 = {T_377,T_535};
  assign T_555 = {T_550,T_377};
  assign T_556 = {T_555,3'h0};
  assign T_557 = {T_556,T_554};
  assign T_570_bits = T_557;
  assign T_570_rd = T_377;
  assign T_570_rs1 = T_377;
  assign T_570_rs2 = T_30;
  assign T_570_rs3 = T_42;
  assign T_576_bits = T_523 ? T_570_bits : T_511_bits;
  assign T_576_rd = T_523 ? T_570_rd : T_511_rd;
  assign T_576_rs1 = T_523 ? T_570_rs1 : T_511_rs1;
  assign T_576_rs2 = T_523 ? T_570_rs2 : T_511_rs2;
  assign T_576_rs3 = T_523 ? T_570_rs3 : T_511_rs3;
  assign T_584 = {T_370,T_375};
  assign T_593 = {T_62,7'h13};
  assign T_594 = {T_584,T_62};
  assign T_595 = {T_594,3'h5};
  assign T_596 = {T_595,T_593};
  assign GEN_0 = {{5'd0}, T_596};
  assign T_613 = GEN_0 | 31'h40000000;
  assign T_630 = {T_376,T_62};
  assign T_631 = {T_630,3'h7};
  assign T_632 = {T_631,T_593};
  assign T_643 = {T_370,T_55};
  assign T_645 = T_643 & 3'h3;
  assign T_647 = T_643 >= 3'h4;
  assign T_649 = T_645 & 3'h1;
  assign T_651 = T_645 >= 3'h2;
  assign T_655 = T_649 >= 3'h1;
  assign T_656 = T_655 ? 2'h3 : 2'h2;
  assign T_662 = T_651 ? T_656 : 2'h0;
  assign T_671 = T_655 ? 3'h7 : 3'h6;
  assign T_676 = T_655 ? 3'h4 : 3'h0;
  assign T_677 = T_651 ? T_671 : T_676;
  assign T_678 = T_647 ? {{1'd0}, T_662} : T_677;
  assign T_681 = T_55 == 2'h0;
  assign T_684 = T_681 ? 31'h40000000 : 31'h0;
  assign T_688 = T_370 ? 7'h3b : 7'h33;
  assign T_698 = {T_62,T_688};
  assign T_699 = {T_30,T_62};
  assign T_700 = {T_699,T_678};
  assign T_701 = {T_700,T_698};
  assign GEN_1 = {{6'd0}, T_701};
  assign T_702 = GEN_1 | T_684;
  assign T_703 = io_in[11:10];
  assign T_705 = T_703 & 2'h1;
  assign T_707 = T_703 >= 2'h2;
  assign T_711 = T_705 >= 2'h1;
  assign T_712 = T_711 ? {{1'd0}, T_702} : T_632;
  assign T_717 = T_711 ? T_613 : {{5'd0}, T_596};
  assign T_718 = T_707 ? T_712 : {{1'd0}, T_717};
  assign T_735_bits = T_718;
  assign T_735_rd = T_62;
  assign T_735_rs1 = T_62;
  assign T_735_rs2 = T_30;
  assign T_735_rs3 = T_42;
  assign T_745 = T_370 ? 10'h3ff : 10'h0;
  assign T_746 = io_in[8];
  assign T_747 = io_in[10:9];
  assign T_749 = io_in[7];
  assign T_751 = io_in[11];
  assign T_752 = io_in[5:3];
  assign T_754 = {T_752,1'h0};
  assign T_755 = {T_543,T_751};
  assign T_756 = {T_755,T_754};
  assign T_757 = {T_20,T_749};
  assign T_758 = {T_745,T_746};
  assign T_759 = {T_758,T_747};
  assign T_760 = {T_759,T_757};
  assign T_761 = {T_760,T_756};
  assign T_762 = T_761[20];
  assign T_784 = T_761[10:1];
  assign T_806 = T_761[11];
  assign T_828 = T_761[19:12];
  assign T_831 = {T_828,5'h0};
  assign T_832 = {T_831,7'h6f};
  assign T_833 = {T_762,T_784};
  assign T_834 = {T_833,T_806};
  assign T_835 = {T_834,T_832};
  assign T_850_bits = T_835;
  assign T_850_rd = 5'h0;
  assign T_850_rs1 = T_62;
  assign T_850_rs2 = T_30;
  assign T_850_rs3 = T_42;
  assign T_860 = T_370 ? 5'h1f : 5'h0;
  assign T_866 = {T_703,T_541};
  assign T_867 = {T_866,1'h0};
  assign T_868 = {T_860,T_55};
  assign T_869 = {T_868,T_543};
  assign T_870 = {T_869,T_867};
  assign T_871 = T_870[12];
  assign T_887 = T_870[10:5];
  assign T_908 = T_870[4:1];
  assign T_924 = T_870[11];
  assign T_926 = {T_924,7'h63};
  assign T_927 = {3'h0,T_908};
  assign T_928 = {T_927,T_926};
  assign T_929 = {5'h0,T_62};
  assign T_930 = {T_871,T_887};
  assign T_931 = {T_930,T_929};
  assign T_932 = {T_931,T_928};
  assign T_947_bits = T_932;
  assign T_947_rd = T_62;
  assign T_947_rs1 = T_62;
  assign T_947_rs2 = 5'h0;
  assign T_947_rs3 = T_42;
  assign T_1024 = {3'h1,T_908};
  assign T_1025 = {T_1024,T_926};
  assign T_1029 = {T_931,T_1025};
  assign T_1042_bits = T_1029;
  assign T_1042_rd = 5'h0;
  assign T_1042_rs1 = T_62;
  assign T_1042_rs2 = 5'h0;
  assign T_1042_rs3 = T_42;
  assign T_1056 = {T_584,T_377};
  assign T_1057 = {T_1056,3'h1};
  assign T_1058 = {T_1057,T_381};
  assign T_1069_bits = {{6'd0}, T_1058};
  assign T_1069_rd = T_377;
  assign T_1069_rs1 = T_377;
  assign T_1069_rs2 = T_375;
  assign T_1069_rs3 = T_42;
  assign T_1079 = {T_55,3'h0};
  assign T_1080 = {T_29,T_370};
  assign T_1081 = {T_1080,T_1079};
  assign T_1086 = {T_377,7'h7};
  assign T_1087 = {T_1081,5'h2};
  assign T_1088 = {T_1087,3'h3};
  assign T_1089 = {T_1088,T_1086};
  assign T_1100_bits = {{3'd0}, T_1089};
  assign T_1100_rd = T_377;
  assign T_1100_rs1 = 5'h2;
  assign T_1100_rs2 = T_375;
  assign T_1100_rs3 = T_42;
  assign T_1106 = io_in[3:2];
  assign T_1108 = io_in[6:4];
  assign T_1110 = {T_1108,2'h0};
  assign T_1111 = {T_1106,T_370};
  assign T_1112 = {T_1111,T_1110};
  assign T_1117 = {T_377,7'h3};
  assign T_1118 = {T_1112,5'h2};
  assign T_1119 = {T_1118,3'h2};
  assign T_1120 = {T_1119,T_1117};
  assign T_1131_bits = {{4'd0}, T_1120};
  assign T_1131_rd = T_377;
  assign T_1131_rs1 = 5'h2;
  assign T_1131_rs2 = T_375;
  assign T_1131_rs3 = T_42;
  assign T_1151 = {T_1088,T_1117};
  assign T_1162_bits = {{3'd0}, T_1151};
  assign T_1162_rd = T_377;
  assign T_1162_rs1 = 5'h2;
  assign T_1162_rs2 = T_375;
  assign T_1162_rs3 = T_42;
  assign T_1173 = {T_377,7'h33};
  assign T_1174 = {T_375,5'h0};
  assign T_1175 = {T_1174,3'h0};
  assign T_1176 = {T_1175,T_1173};
  assign T_1187_bits = {{7'd0}, T_1176};
  assign T_1187_rd = T_377;
  assign T_1187_rs1 = 5'h0;
  assign T_1187_rs2 = T_375;
  assign T_1187_rs3 = T_42;
  assign T_1199 = {T_375,T_377};
  assign T_1200 = {T_1199,3'h0};
  assign T_1201 = {T_1200,T_1173};
  assign T_1212_bits = {{7'd0}, T_1201};
  assign T_1212_rd = T_377;
  assign T_1212_rs1 = T_377;
  assign T_1212_rs2 = T_375;
  assign T_1212_rs3 = T_42;
  assign T_1226 = {T_1200,12'h67};
  assign T_1227 = T_1226[24:7];
  assign T_1229 = {T_1227,7'h1f};
  assign T_1233 = T_405 ? T_1226 : T_1229;
  assign T_1244_bits = {{7'd0}, T_1233};
  assign T_1244_rd = 5'h0;
  assign T_1244_rs1 = T_377;
  assign T_1244_rs2 = T_375;
  assign T_1244_rs3 = T_42;
  assign T_1252 = T_375 != 5'h0;
  assign T_1253_bits = T_1252 ? T_1187_bits : T_1244_bits;
  assign T_1253_rd = T_1252 ? T_1187_rd : T_1244_rd;
  assign T_1253_rs1 = T_1252 ? T_1187_rs1 : T_1244_rs1;
  assign T_1253_rs2 = T_1252 ? T_1187_rs2 : T_1244_rs2;
  assign T_1253_rs3 = T_1252 ? T_1187_rs3 : T_1244_rs3;
  assign T_1267 = {T_1200,12'he7};
  assign T_1270 = {T_1227,7'h73};
  assign T_1272 = T_1270 | 25'h100000;
  assign T_1276 = T_405 ? T_1267 : T_1272;
  assign T_1287_bits = {{7'd0}, T_1276};
  assign T_1287_rd = 5'h1;
  assign T_1287_rs1 = T_377;
  assign T_1287_rs2 = T_375;
  assign T_1287_rs3 = T_42;
  assign T_1296_bits = T_1252 ? T_1212_bits : T_1287_bits;
  assign T_1296_rd = T_1252 ? T_1212_rd : T_1287_rd;
  assign T_1296_rs1 = T_1252 ? T_1212_rs1 : T_1287_rs1;
  assign T_1296_rs2 = T_1252 ? T_1212_rs2 : T_1287_rs2;
  assign T_1296_rs3 = T_1252 ? T_1212_rs3 : T_1287_rs3;
  assign T_1303_bits = T_370 ? T_1296_bits : T_1253_bits;
  assign T_1303_rd = T_370 ? T_1296_rd : T_1253_rd;
  assign T_1303_rs1 = T_370 ? T_1296_rs1 : T_1253_rs1;
  assign T_1303_rs2 = T_370 ? T_1296_rs2 : T_1253_rs2;
  assign T_1303_rs3 = T_370 ? T_1296_rs3 : T_1253_rs3;
  assign T_1312 = {T_61,T_56};
  assign T_1313 = {T_1312,3'h0};
  assign T_1314 = T_1313[8:5];
  assign T_1323 = T_1313[4:0];
  assign T_1325 = {3'h3,T_1323};
  assign T_1326 = {T_1325,7'h27};
  assign T_1327 = {T_1314,T_375};
  assign T_1328 = {T_1327,5'h2};
  assign T_1329 = {T_1328,T_1326};
  assign T_1340_bits = {{3'd0}, T_1329};
  assign T_1340_rd = T_377;
  assign T_1340_rs1 = 5'h2;
  assign T_1340_rs2 = T_375;
  assign T_1340_rs3 = T_42;
  assign T_1346 = io_in[8:7];
  assign T_1347 = io_in[12:9];
  assign T_1349 = {T_1346,T_1347};
  assign T_1350 = {T_1349,2'h0};
  assign T_1351 = T_1350[7:5];
  assign T_1360 = T_1350[4:0];
  assign T_1362 = {3'h2,T_1360};
  assign T_1363 = {T_1362,7'h23};
  assign T_1364 = {T_1351,T_375};
  assign T_1365 = {T_1364,5'h2};
  assign T_1366 = {T_1365,T_1363};
  assign T_1377_bits = {{4'd0}, T_1366};
  assign T_1377_rd = T_377;
  assign T_1377_rs1 = 5'h2;
  assign T_1377_rs2 = T_375;
  assign T_1377_rs3 = T_42;
  assign T_1400 = {T_1325,7'h23};
  assign T_1403 = {T_1328,T_1400};
  assign T_1414_bits = {{3'd0}, T_1403};
  assign T_1414_rd = T_377;
  assign T_1414_rs1 = 5'h2;
  assign T_1414_rs2 = T_375;
  assign T_1414_rs3 = T_42;
  assign T_1421 = io_in[19:15];
  assign T_1422 = io_in[24:20];
  assign T_1430_bits = io_in;
  assign T_1430_rd = T_377;
  assign T_1430_rs1 = T_1421;
  assign T_1430_rs2 = T_1422;
  assign T_1430_rs3 = T_42;
  assign T_1446_bits = io_in;
  assign T_1446_rd = T_377;
  assign T_1446_rs1 = T_1421;
  assign T_1446_rs2 = T_1422;
  assign T_1446_rs3 = T_42;
  assign T_1462_bits = io_in;
  assign T_1462_rd = T_377;
  assign T_1462_rs1 = T_1421;
  assign T_1462_rs2 = T_1422;
  assign T_1462_rs3 = T_42;
  assign T_1478_bits = io_in;
  assign T_1478_rd = T_377;
  assign T_1478_rs1 = T_1421;
  assign T_1478_rs2 = T_1422;
  assign T_1478_rs3 = T_42;
  assign T_1494_bits = io_in;
  assign T_1494_rd = T_377;
  assign T_1494_rs1 = T_1421;
  assign T_1494_rs2 = T_1422;
  assign T_1494_rs3 = T_42;
  assign T_1510_bits = io_in;
  assign T_1510_rd = T_377;
  assign T_1510_rs1 = T_1421;
  assign T_1510_rs2 = T_1422;
  assign T_1510_rs3 = T_42;
  assign T_1526_bits = io_in;
  assign T_1526_rd = T_377;
  assign T_1526_rs1 = T_1421;
  assign T_1526_rs2 = T_1422;
  assign T_1526_rs3 = T_42;
  assign T_1542_bits = io_in;
  assign T_1542_rd = T_377;
  assign T_1542_rs1 = T_1421;
  assign T_1542_rs2 = T_1422;
  assign T_1542_rs3 = T_42;
  assign T_1549 = io_in[15:13];
  assign T_1550 = {T_8,T_1549};
  assign T_1552 = T_1550 & 5'hf;
  assign T_1554 = T_1550 >= 5'h10;
  assign T_1556 = T_1552 & 5'h7;
  assign T_1558 = T_1552 >= 5'h8;
  assign T_1560 = T_1556 & 5'h3;
  assign T_1562 = T_1556 >= 5'h4;
  assign T_1564 = T_1560 & 5'h1;
  assign T_1566 = T_1560 >= 5'h2;
  assign T_1570 = T_1564 >= 5'h1;
  assign T_1571_bits = T_1570 ? T_1542_bits : T_1526_bits;
  assign T_1571_rd = T_1570 ? T_1542_rd : T_1526_rd;
  assign T_1571_rs1 = T_1570 ? T_1542_rs1 : T_1526_rs1;
  assign T_1571_rs2 = T_1570 ? T_1542_rs2 : T_1526_rs2;
  assign T_1571_rs3 = T_1570 ? T_1542_rs3 : T_1526_rs3;
  assign T_1581_bits = T_1570 ? T_1510_bits : T_1494_bits;
  assign T_1581_rd = T_1570 ? T_1510_rd : T_1494_rd;
  assign T_1581_rs1 = T_1570 ? T_1510_rs1 : T_1494_rs1;
  assign T_1581_rs2 = T_1570 ? T_1510_rs2 : T_1494_rs2;
  assign T_1581_rs3 = T_1570 ? T_1510_rs3 : T_1494_rs3;
  assign T_1587_bits = T_1566 ? T_1571_bits : T_1581_bits;
  assign T_1587_rd = T_1566 ? T_1571_rd : T_1581_rd;
  assign T_1587_rs1 = T_1566 ? T_1571_rs1 : T_1581_rs1;
  assign T_1587_rs2 = T_1566 ? T_1571_rs2 : T_1581_rs2;
  assign T_1587_rs3 = T_1566 ? T_1571_rs3 : T_1581_rs3;
  assign T_1601_bits = T_1570 ? T_1478_bits : T_1462_bits;
  assign T_1601_rd = T_1570 ? T_1478_rd : T_1462_rd;
  assign T_1601_rs1 = T_1570 ? T_1478_rs1 : T_1462_rs1;
  assign T_1601_rs2 = T_1570 ? T_1478_rs2 : T_1462_rs2;
  assign T_1601_rs3 = T_1570 ? T_1478_rs3 : T_1462_rs3;
  assign T_1611_bits = T_1570 ? T_1446_bits : T_1430_bits;
  assign T_1611_rd = T_1570 ? T_1446_rd : T_1430_rd;
  assign T_1611_rs1 = T_1570 ? T_1446_rs1 : T_1430_rs1;
  assign T_1611_rs2 = T_1570 ? T_1446_rs2 : T_1430_rs2;
  assign T_1611_rs3 = T_1570 ? T_1446_rs3 : T_1430_rs3;
  assign T_1617_bits = T_1566 ? T_1601_bits : T_1611_bits;
  assign T_1617_rd = T_1566 ? T_1601_rd : T_1611_rd;
  assign T_1617_rs1 = T_1566 ? T_1601_rs1 : T_1611_rs1;
  assign T_1617_rs2 = T_1566 ? T_1601_rs2 : T_1611_rs2;
  assign T_1617_rs3 = T_1566 ? T_1601_rs3 : T_1611_rs3;
  assign T_1623_bits = T_1562 ? T_1587_bits : T_1617_bits;
  assign T_1623_rd = T_1562 ? T_1587_rd : T_1617_rd;
  assign T_1623_rs1 = T_1562 ? T_1587_rs1 : T_1617_rs1;
  assign T_1623_rs2 = T_1562 ? T_1587_rs2 : T_1617_rs2;
  assign T_1623_rs3 = T_1562 ? T_1587_rs3 : T_1617_rs3;
  assign T_1641_bits = T_1570 ? T_1414_bits : T_1377_bits;
  assign T_1641_rd = T_1570 ? T_1414_rd : T_1377_rd;
  assign T_1641_rs1 = T_1570 ? T_1414_rs1 : T_1377_rs1;
  assign T_1641_rs2 = T_1570 ? T_1414_rs2 : T_1377_rs2;
  assign T_1641_rs3 = T_1570 ? T_1414_rs3 : T_1377_rs3;
  assign T_1651_bits = T_1570 ? T_1340_bits : T_1303_bits;
  assign T_1651_rd = T_1570 ? T_1340_rd : T_1303_rd;
  assign T_1651_rs1 = T_1570 ? T_1340_rs1 : T_1303_rs1;
  assign T_1651_rs2 = T_1570 ? T_1340_rs2 : T_1303_rs2;
  assign T_1651_rs3 = T_1570 ? T_1340_rs3 : T_1303_rs3;
  assign T_1657_bits = T_1566 ? T_1641_bits : T_1651_bits;
  assign T_1657_rd = T_1566 ? T_1641_rd : T_1651_rd;
  assign T_1657_rs1 = T_1566 ? T_1641_rs1 : T_1651_rs1;
  assign T_1657_rs2 = T_1566 ? T_1641_rs2 : T_1651_rs2;
  assign T_1657_rs3 = T_1566 ? T_1641_rs3 : T_1651_rs3;
  assign T_1671_bits = T_1570 ? T_1162_bits : T_1131_bits;
  assign T_1671_rd = T_1570 ? T_1162_rd : T_1131_rd;
  assign T_1671_rs1 = T_1570 ? T_1162_rs1 : T_1131_rs1;
  assign T_1671_rs2 = T_1570 ? T_1162_rs2 : T_1131_rs2;
  assign T_1671_rs3 = T_1570 ? T_1162_rs3 : T_1131_rs3;
  assign T_1681_bits = T_1570 ? T_1100_bits : T_1069_bits;
  assign T_1681_rd = T_1570 ? T_1100_rd : T_1069_rd;
  assign T_1681_rs1 = T_1570 ? T_1100_rs1 : T_1069_rs1;
  assign T_1681_rs2 = T_1570 ? T_1100_rs2 : T_1069_rs2;
  assign T_1681_rs3 = T_1570 ? T_1100_rs3 : T_1069_rs3;
  assign T_1687_bits = T_1566 ? T_1671_bits : T_1681_bits;
  assign T_1687_rd = T_1566 ? T_1671_rd : T_1681_rd;
  assign T_1687_rs1 = T_1566 ? T_1671_rs1 : T_1681_rs1;
  assign T_1687_rs2 = T_1566 ? T_1671_rs2 : T_1681_rs2;
  assign T_1687_rs3 = T_1566 ? T_1671_rs3 : T_1681_rs3;
  assign T_1693_bits = T_1562 ? T_1657_bits : T_1687_bits;
  assign T_1693_rd = T_1562 ? T_1657_rd : T_1687_rd;
  assign T_1693_rs1 = T_1562 ? T_1657_rs1 : T_1687_rs1;
  assign T_1693_rs2 = T_1562 ? T_1657_rs2 : T_1687_rs2;
  assign T_1693_rs3 = T_1562 ? T_1657_rs3 : T_1687_rs3;
  assign T_1699_bits = T_1558 ? T_1623_bits : T_1693_bits;
  assign T_1699_rd = T_1558 ? T_1623_rd : T_1693_rd;
  assign T_1699_rs1 = T_1558 ? T_1623_rs1 : T_1693_rs1;
  assign T_1699_rs2 = T_1558 ? T_1623_rs2 : T_1693_rs2;
  assign T_1699_rs3 = T_1558 ? T_1623_rs3 : T_1693_rs3;
  assign T_1721_bits = T_1570 ? T_1042_bits : T_947_bits;
  assign T_1721_rd = T_1570 ? T_1042_rd : T_947_rd;
  assign T_1721_rs1 = T_1570 ? T_1042_rs1 : T_947_rs1;
  assign T_1721_rs2 = T_1570 ? T_1042_rs2 : T_947_rs2;
  assign T_1721_rs3 = T_1570 ? T_1042_rs3 : T_947_rs3;
  assign T_1731_bits = T_1570 ? T_850_bits : T_735_bits;
  assign T_1731_rd = T_1570 ? T_850_rd : T_735_rd;
  assign T_1731_rs1 = T_1570 ? T_850_rs1 : T_735_rs1;
  assign T_1731_rs2 = T_1570 ? T_850_rs2 : T_735_rs2;
  assign T_1731_rs3 = T_1570 ? T_850_rs3 : T_735_rs3;
  assign T_1737_bits = T_1566 ? T_1721_bits : T_1731_bits;
  assign T_1737_rd = T_1566 ? T_1721_rd : T_1731_rd;
  assign T_1737_rs1 = T_1566 ? T_1721_rs1 : T_1731_rs1;
  assign T_1737_rs2 = T_1566 ? T_1721_rs2 : T_1731_rs2;
  assign T_1737_rs3 = T_1566 ? T_1721_rs3 : T_1731_rs3;
  assign T_1751_bits = T_1570 ? T_576_bits : T_468_bits;
  assign T_1751_rd = T_1570 ? T_576_rd : T_468_rd;
  assign T_1751_rs1 = T_1570 ? T_576_rs1 : T_468_rs1;
  assign T_1751_rs2 = T_1570 ? T_576_rs2 : T_468_rs2;
  assign T_1751_rs3 = T_1570 ? T_576_rs3 : T_468_rs3;
  assign T_1761_bits = T_1570 ? T_435_bits : T_397_bits;
  assign T_1761_rd = T_1570 ? T_435_rd : T_397_rd;
  assign T_1761_rs1 = T_1570 ? T_435_rs1 : T_397_rs1;
  assign T_1761_rs2 = T_1570 ? T_435_rs2 : T_397_rs2;
  assign T_1761_rs3 = T_1570 ? T_435_rs3 : T_397_rs3;
  assign T_1767_bits = T_1566 ? T_1751_bits : T_1761_bits;
  assign T_1767_rd = T_1566 ? T_1751_rd : T_1761_rd;
  assign T_1767_rs1 = T_1566 ? T_1751_rs1 : T_1761_rs1;
  assign T_1767_rs2 = T_1566 ? T_1751_rs2 : T_1761_rs2;
  assign T_1767_rs3 = T_1566 ? T_1751_rs3 : T_1761_rs3;
  assign T_1773_bits = T_1562 ? T_1737_bits : T_1767_bits;
  assign T_1773_rd = T_1562 ? T_1737_rd : T_1767_rd;
  assign T_1773_rs1 = T_1562 ? T_1737_rs1 : T_1767_rs1;
  assign T_1773_rs2 = T_1562 ? T_1737_rs2 : T_1767_rs2;
  assign T_1773_rs3 = T_1562 ? T_1737_rs3 : T_1767_rs3;
  assign T_1791_bits = T_1570 ? T_364_bits : T_317_bits;
  assign T_1791_rd = T_1570 ? T_364_rd : T_317_rd;
  assign T_1791_rs1 = T_1570 ? T_364_rs1 : T_317_rs1;
  assign T_1791_rs2 = T_1570 ? T_364_rs2 : T_317_rs2;
  assign T_1791_rs3 = T_1570 ? T_364_rs3 : T_317_rs3;
  assign T_1801_bits = T_1570 ? T_266_bits : T_219_bits;
  assign T_1801_rd = T_1570 ? T_266_rd : T_219_rd;
  assign T_1801_rs1 = T_1570 ? T_266_rs1 : T_219_rs1;
  assign T_1801_rs2 = T_1570 ? T_266_rs2 : T_219_rs2;
  assign T_1801_rs3 = T_1570 ? T_266_rs3 : T_219_rs3;
  assign T_1807_bits = T_1566 ? T_1791_bits : T_1801_bits;
  assign T_1807_rd = T_1566 ? T_1791_rd : T_1801_rd;
  assign T_1807_rs1 = T_1566 ? T_1791_rs1 : T_1801_rs1;
  assign T_1807_rs2 = T_1566 ? T_1791_rs2 : T_1801_rs2;
  assign T_1807_rs3 = T_1566 ? T_1791_rs3 : T_1801_rs3;
  assign T_1821_bits = T_1570 ? T_168_bits : T_129_bits;
  assign T_1821_rd = T_1570 ? T_168_rd : T_129_rd;
  assign T_1821_rs1 = T_1570 ? T_168_rs1 : T_129_rs1;
  assign T_1821_rs2 = T_1570 ? T_168_rs2 : T_129_rs2;
  assign T_1821_rs3 = T_1570 ? T_168_rs3 : T_129_rs3;
  assign T_1831_bits = T_1570 ? T_88_bits : T_49_bits;
  assign T_1831_rd = T_1570 ? T_88_rd : T_49_rd;
  assign T_1831_rs1 = T_1570 ? T_88_rs1 : T_49_rs1;
  assign T_1831_rs2 = T_1570 ? T_88_rs2 : T_49_rs2;
  assign T_1831_rs3 = T_1570 ? T_88_rs3 : T_49_rs3;
  assign T_1837_bits = T_1566 ? T_1821_bits : T_1831_bits;
  assign T_1837_rd = T_1566 ? T_1821_rd : T_1831_rd;
  assign T_1837_rs1 = T_1566 ? T_1821_rs1 : T_1831_rs1;
  assign T_1837_rs2 = T_1566 ? T_1821_rs2 : T_1831_rs2;
  assign T_1837_rs3 = T_1566 ? T_1821_rs3 : T_1831_rs3;
  assign T_1843_bits = T_1562 ? T_1807_bits : T_1837_bits;
  assign T_1843_rd = T_1562 ? T_1807_rd : T_1837_rd;
  assign T_1843_rs1 = T_1562 ? T_1807_rs1 : T_1837_rs1;
  assign T_1843_rs2 = T_1562 ? T_1807_rs2 : T_1837_rs2;
  assign T_1843_rs3 = T_1562 ? T_1807_rs3 : T_1837_rs3;
  assign T_1849_bits = T_1558 ? T_1773_bits : T_1843_bits;
  assign T_1849_rd = T_1558 ? T_1773_rd : T_1843_rd;
  assign T_1849_rs1 = T_1558 ? T_1773_rs1 : T_1843_rs1;
  assign T_1849_rs2 = T_1558 ? T_1773_rs2 : T_1843_rs2;
  assign T_1849_rs3 = T_1558 ? T_1773_rs3 : T_1843_rs3;
  assign T_1855_bits = T_1554 ? T_1699_bits : T_1849_bits;
  assign T_1855_rd = T_1554 ? T_1699_rd : T_1849_rd;
  assign T_1855_rs1 = T_1554 ? T_1699_rs1 : T_1849_rs1;
  assign T_1855_rs2 = T_1554 ? T_1699_rs2 : T_1849_rs2;
  assign T_1855_rs3 = T_1554 ? T_1699_rs3 : T_1849_rs3;
endmodule
module IBuf(
  input   clk,
  input   reset,
  output  io_imem_ready,
  input   io_imem_valid,
  input   io_imem_bits_btb_valid,
  input   io_imem_bits_btb_bits_taken,
  input  [1:0] io_imem_bits_btb_bits_mask,
  input   io_imem_bits_btb_bits_bridx,
  input  [38:0] io_imem_bits_btb_bits_target,
  input  [5:0] io_imem_bits_btb_bits_entry,
  input  [6:0] io_imem_bits_btb_bits_bht_history,
  input  [1:0] io_imem_bits_btb_bits_bht_value,
  input  [39:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input  [1:0] io_imem_bits_mask,
  input   io_imem_bits_xcpt_if,
  input   io_imem_bits_replay,
  input   io_kill,
  output [39:0] io_pc,
  output  io_btb_resp_taken,
  output [1:0] io_btb_resp_mask,
  output  io_btb_resp_bridx,
  output [38:0] io_btb_resp_target,
  output [5:0] io_btb_resp_entry,
  output [6:0] io_btb_resp_bht_history,
  output [1:0] io_btb_resp_bht_value,
  input   io_inst_0_ready,
  output  io_inst_0_valid,
  output  io_inst_0_bits_pf0,
  output  io_inst_0_bits_pf1,
  output  io_inst_0_bits_replay,
  output  io_inst_0_bits_btb_hit,
  output  io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0] io_inst_0_bits_inst_rd,
  output [4:0] io_inst_0_bits_inst_rs1,
  output [4:0] io_inst_0_bits_inst_rs2,
  output [4:0] io_inst_0_bits_inst_rs3
);
  reg  nBufValid;
  reg [31:0] GEN_33;
  reg  buf_btb_valid;
  reg [31:0] GEN_34;
  reg  buf_btb_bits_taken;
  reg [31:0] GEN_35;
  reg [1:0] buf_btb_bits_mask;
  reg [31:0] GEN_36;
  reg  buf_btb_bits_bridx;
  reg [31:0] GEN_37;
  reg [38:0] buf_btb_bits_target;
  reg [63:0] GEN_38;
  reg [5:0] buf_btb_bits_entry;
  reg [31:0] GEN_43;
  reg [6:0] buf_btb_bits_bht_history;
  reg [31:0] GEN_44;
  reg [1:0] buf_btb_bits_bht_value;
  reg [31:0] GEN_48;
  reg [39:0] buf_pc;
  reg [63:0] GEN_51;
  reg [31:0] buf_data;
  reg [31:0] GEN_52;
  reg [1:0] buf_mask;
  reg [31:0] GEN_53;
  reg  buf_xcpt_if;
  reg [31:0] GEN_54;
  reg  buf_replay;
  reg [31:0] GEN_55;
  reg  ibufBTBHit;
  reg [31:0] GEN_56;
  reg  ibufBTBResp_taken;
  reg [31:0] GEN_57;
  reg [1:0] ibufBTBResp_mask;
  reg [31:0] GEN_58;
  reg  ibufBTBResp_bridx;
  reg [31:0] GEN_59;
  reg [38:0] ibufBTBResp_target;
  reg [63:0] GEN_60;
  reg [5:0] ibufBTBResp_entry;
  reg [31:0] GEN_61;
  reg [6:0] ibufBTBResp_bht_history;
  reg [31:0] GEN_62;
  reg [1:0] ibufBTBResp_bht_value;
  reg [31:0] GEN_63;
  wire  pcWordBits;
  wire [1:0] nReady;
  wire  T_375;
  wire [1:0] T_377;
  wire [1:0] T_379;
  wire [1:0] GEN_31;
  wire [2:0] T_380;
  wire [1:0] nIC;
  wire [1:0] GEN_32;
  wire [2:0] T_381;
  wire [1:0] nICReady;
  wire [1:0] T_383;
  wire [2:0] T_384;
  wire [1:0] nValid;
  wire  T_385;
  wire  T_386;
  wire [2:0] T_388;
  wire [1:0] T_389;
  wire  T_390;
  wire  T_391;
  wire  T_392;
  wire [2:0] T_395;
  wire [1:0] T_396;
  wire [1:0] T_397;
  wire  T_399;
  wire  T_400;
  wire  T_401;
  wire  T_406;
  wire [2:0] T_407;
  wire [1:0] T_408;
  wire [15:0] T_411;
  wire [31:0] T_412;
  wire [63:0] T_413;
  wire [5:0] GEN_39;
  wire [5:0] T_414;
  wire [63:0] T_415;
  wire [15:0] T_416;
  wire [39:0] T_418;
  wire [2:0] GEN_40;
  wire [2:0] T_419;
  wire [39:0] GEN_41;
  wire [40:0] T_420;
  wire [39:0] T_421;
  wire [39:0] T_422;
  wire [39:0] T_423;
  wire [1:0] GEN_42;
  wire [2:0] T_424;
  wire [1:0] T_425;
  wire  GEN_0;
  wire [1:0] GEN_1;
  wire [1:0] GEN_2;
  wire [38:0] GEN_3;
  wire [5:0] GEN_4;
  wire [6:0] GEN_5;
  wire [1:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire [5:0] GEN_13;
  wire [6:0] GEN_14;
  wire [1:0] GEN_15;
  wire [39:0] GEN_16;
  wire [31:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [38:0] GEN_25;
  wire [5:0] GEN_26;
  wire [6:0] GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [2:0] T_428;
  wire [1:0] T_429;
  wire [2:0] T_430;
  wire [1:0] T_431;
  wire [15:0] T_432;
  wire [31:0] T_433;
  wire [63:0] T_434;
  wire [15:0] T_435;
  wire [31:0] T_436;
  wire [63:0] T_437;
  wire [127:0] T_438;
  wire [5:0] GEN_45;
  wire [5:0] T_439;
  wire [190:0] GEN_46;
  wire [190:0] T_440;
  wire [31:0] icData;
  wire [4:0] GEN_47;
  wire [4:0] T_443;
  wire [62:0] T_444;
  wire [31:0] icMask;
  wire [31:0] T_445;
  wire [31:0] T_446;
  wire [31:0] T_447;
  wire [31:0] inst;
  wire [3:0] T_449;
  wire [4:0] T_451;
  wire [3:0] T_452;
  wire [1:0] valid;
  wire [1:0] T_454;
  wire [2:0] T_456;
  wire [1:0] bufMask;
  wire [1:0] T_458;
  wire [1:0] T_459;
  wire [1:0] T_461;
  wire [1:0] T_462;
  wire [1:0] xcpt_if;
  wire [1:0] T_464;
  wire [1:0] T_467;
  wire [1:0] T_468;
  wire [1:0] ic_replay;
  wire [1:0] T_470;
  wire [1:0] ibufBTBHitMask;
  wire [1:0] T_472;
  wire [2:0] T_473;
  wire [1:0] T_474;
  wire [3:0] T_476;
  wire [3:0] icBTBHitMask;
  wire [1:0] T_478;
  wire [3:0] GEN_49;
  wire [3:0] T_480;
  wire [3:0] GEN_50;
  wire [3:0] btbHitMask;
  wire  T_483;
  wire  T_484_taken;
  wire [1:0] T_484_mask;
  wire  T_484_bridx;
  wire [38:0] T_484_target;
  wire [5:0] T_484_entry;
  wire [6:0] T_484_bht_history;
  wire [1:0] T_484_bht_value;
  wire  T_494;
  wire [39:0] T_495;
  wire  RVCExpander_1_clk;
  wire  RVCExpander_1_reset;
  wire [31:0] RVCExpander_1_io_in;
  wire [31:0] RVCExpander_1_io_out_bits;
  wire [4:0] RVCExpander_1_io_out_rd;
  wire [4:0] RVCExpander_1_io_out_rs1;
  wire [4:0] RVCExpander_1_io_out_rs2;
  wire [4:0] RVCExpander_1_io_out_rs3;
  wire  RVCExpander_1_io_rvc;
  wire [1:0] T_497;
  wire  T_498;
  wire  T_500;
  wire [3:0] T_501;
  wire  T_502;
  wire [1:0] T_504;
  wire  T_505;
  wire [1:0] T_506;
  wire  T_507;
  wire  T_508;
  wire  T_509;
  wire  T_510;
  wire [1:0] T_511;
  wire  T_512;
  wire [1:0] T_516;
  wire  T_517;
  wire  T_518;
  wire [1:0] T_522;
  wire  T_523;
  wire  T_524;
  wire  T_525;
  wire  T_526;
  wire [1:0] T_527;
  wire  T_528;
  wire  T_536;
  wire [3:0] T_544;
  wire  T_545;
  wire  T_546;
  wire  T_547;
  wire  T_548;
  wire [2:0] T_553;
  wire [1:0] T_554;
  wire [1:0] T_555;
  wire [1:0] GEN_30;
  RVCExpander RVCExpander_1 (
    .clk(RVCExpander_1_clk),
    .reset(RVCExpander_1_reset),
    .io_in(RVCExpander_1_io_in),
    .io_out_bits(RVCExpander_1_io_out_bits),
    .io_out_rd(RVCExpander_1_io_out_rd),
    .io_out_rs1(RVCExpander_1_io_out_rs1),
    .io_out_rs2(RVCExpander_1_io_out_rs2),
    .io_out_rs3(RVCExpander_1_io_out_rs3),
    .io_rvc(RVCExpander_1_io_rvc)
  );
  assign io_imem_ready = T_392;
  assign io_pc = T_495;
  assign io_btb_resp_taken = T_484_taken;
  assign io_btb_resp_mask = T_484_mask;
  assign io_btb_resp_bridx = T_484_bridx;
  assign io_btb_resp_target = T_484_target;
  assign io_btb_resp_entry = T_484_entry;
  assign io_btb_resp_bht_history = T_484_bht_history;
  assign io_btb_resp_bht_value = T_484_bht_value;
  assign io_inst_0_valid = T_526;
  assign io_inst_0_bits_pf0 = T_528;
  assign io_inst_0_bits_pf1 = T_536;
  assign io_inst_0_bits_replay = T_510;
  assign io_inst_0_bits_btb_hit = T_547;
  assign io_inst_0_bits_rvc = RVCExpander_1_io_rvc;
  assign io_inst_0_bits_inst_bits = RVCExpander_1_io_out_bits;
  assign io_inst_0_bits_inst_rd = RVCExpander_1_io_out_rd;
  assign io_inst_0_bits_inst_rs1 = RVCExpander_1_io_out_rs1;
  assign io_inst_0_bits_inst_rs2 = RVCExpander_1_io_out_rs2;
  assign io_inst_0_bits_inst_rs3 = RVCExpander_1_io_out_rs3;
  assign pcWordBits = io_imem_bits_pc[1];
  assign nReady = GEN_30;
  assign T_375 = io_imem_bits_btb_valid & io_imem_bits_btb_bits_taken;
  assign T_377 = io_imem_bits_btb_bits_bridx + 1'h1;
  assign T_379 = T_375 ? T_377 : 2'h2;
  assign GEN_31 = {{1'd0}, pcWordBits};
  assign T_380 = T_379 - GEN_31;
  assign nIC = T_380[1:0];
  assign GEN_32 = {{1'd0}, nBufValid};
  assign T_381 = nReady - GEN_32;
  assign nICReady = T_381[1:0];
  assign T_383 = io_imem_valid ? nIC : 2'h0;
  assign T_384 = T_383 + GEN_32;
  assign nValid = T_384[1:0];
  assign T_385 = nReady >= GEN_32;
  assign T_386 = nICReady >= nIC;
  assign T_388 = nIC - nICReady;
  assign T_389 = T_388[1:0];
  assign T_390 = 2'h1 >= T_389;
  assign T_391 = T_386 | T_390;
  assign T_392 = T_385 & T_391;
  assign T_395 = GEN_32 - nReady;
  assign T_396 = T_395[1:0];
  assign T_397 = T_385 ? 2'h0 : T_396;
  assign T_399 = io_imem_valid & T_385;
  assign T_400 = nICReady < nIC;
  assign T_401 = T_399 & T_400;
  assign T_406 = T_401 & T_390;
  assign T_407 = GEN_31 + nICReady;
  assign T_408 = T_407[1:0];
  assign T_411 = io_imem_bits_data[31:16];
  assign T_412 = {T_411,T_411};
  assign T_413 = {T_412,io_imem_bits_data};
  assign GEN_39 = {{4'd0}, T_408};
  assign T_414 = GEN_39 << 4;
  assign T_415 = T_413 >> T_414;
  assign T_416 = T_415[15:0];
  assign T_418 = io_imem_bits_pc & 40'hfffffffffc;
  assign GEN_40 = {{1'd0}, nICReady};
  assign T_419 = GEN_40 << 1;
  assign GEN_41 = {{37'd0}, T_419};
  assign T_420 = io_imem_bits_pc + GEN_41;
  assign T_421 = T_420[39:0];
  assign T_422 = T_421 & 40'h3;
  assign T_423 = T_418 | T_422;
  assign GEN_42 = {{1'd0}, io_imem_bits_btb_bits_bridx};
  assign T_424 = GEN_42 + nICReady;
  assign T_425 = T_424[1:0];
  assign GEN_0 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_taken : ibufBTBResp_taken;
  assign GEN_1 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_mask : ibufBTBResp_mask;
  assign GEN_2 = io_imem_bits_btb_valid ? T_425 : {{1'd0}, ibufBTBResp_bridx};
  assign GEN_3 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_target : ibufBTBResp_target;
  assign GEN_4 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_entry : ibufBTBResp_entry;
  assign GEN_5 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_bht_history : ibufBTBResp_bht_history;
  assign GEN_6 = io_imem_bits_btb_valid ? io_imem_bits_btb_bits_bht_value : ibufBTBResp_bht_value;
  assign GEN_7 = T_406 ? T_389 : T_397;
  assign GEN_8 = T_406 ? io_imem_bits_btb_valid : buf_btb_valid;
  assign GEN_9 = T_406 ? io_imem_bits_btb_bits_taken : buf_btb_bits_taken;
  assign GEN_10 = T_406 ? io_imem_bits_btb_bits_mask : buf_btb_bits_mask;
  assign GEN_11 = T_406 ? io_imem_bits_btb_bits_bridx : buf_btb_bits_bridx;
  assign GEN_12 = T_406 ? io_imem_bits_btb_bits_target : buf_btb_bits_target;
  assign GEN_13 = T_406 ? io_imem_bits_btb_bits_entry : buf_btb_bits_entry;
  assign GEN_14 = T_406 ? io_imem_bits_btb_bits_bht_history : buf_btb_bits_bht_history;
  assign GEN_15 = T_406 ? io_imem_bits_btb_bits_bht_value : buf_btb_bits_bht_value;
  assign GEN_16 = T_406 ? T_423 : buf_pc;
  assign GEN_17 = T_406 ? {{16'd0}, T_416} : buf_data;
  assign GEN_18 = T_406 ? io_imem_bits_mask : buf_mask;
  assign GEN_19 = T_406 ? io_imem_bits_xcpt_if : buf_xcpt_if;
  assign GEN_20 = T_406 ? io_imem_bits_replay : buf_replay;
  assign GEN_21 = T_406 ? io_imem_bits_btb_valid : ibufBTBHit;
  assign GEN_22 = T_406 ? GEN_0 : ibufBTBResp_taken;
  assign GEN_23 = T_406 ? GEN_1 : ibufBTBResp_mask;
  assign GEN_24 = T_406 ? GEN_2 : {{1'd0}, ibufBTBResp_bridx};
  assign GEN_25 = T_406 ? GEN_3 : ibufBTBResp_target;
  assign GEN_26 = T_406 ? GEN_4 : ibufBTBResp_entry;
  assign GEN_27 = T_406 ? GEN_5 : ibufBTBResp_bht_history;
  assign GEN_28 = T_406 ? GEN_6 : ibufBTBResp_bht_value;
  assign GEN_29 = io_kill ? 2'h0 : GEN_7;
  assign T_428 = 2'h2 + GEN_32;
  assign T_429 = T_428[1:0];
  assign T_430 = T_429 - GEN_31;
  assign T_431 = T_430[1:0];
  assign T_432 = io_imem_bits_data[15:0];
  assign T_433 = {T_432,T_432};
  assign T_434 = {io_imem_bits_data,T_433};
  assign T_435 = T_434[63:48];
  assign T_436 = {T_435,T_435};
  assign T_437 = {T_436,T_436};
  assign T_438 = {T_437,T_434};
  assign GEN_45 = {{4'd0}, T_431};
  assign T_439 = GEN_45 << 4;
  assign GEN_46 = {{63'd0}, T_438};
  assign T_440 = GEN_46 << T_439;
  assign icData = T_440[95:64];
  assign GEN_47 = {{4'd0}, nBufValid};
  assign T_443 = GEN_47 << 4;
  assign T_444 = 63'hffffffff << T_443;
  assign icMask = T_444[31:0];
  assign T_445 = icData & icMask;
  assign T_446 = ~ icMask;
  assign T_447 = buf_data & T_446;
  assign inst = T_445 | T_447;
  assign T_449 = 4'h1 << nValid;
  assign T_451 = T_449 - 4'h1;
  assign T_452 = T_451[3:0];
  assign valid = T_452[1:0];
  assign T_454 = 2'h1 << nBufValid;
  assign T_456 = T_454 - 2'h1;
  assign bufMask = T_456[1:0];
  assign T_458 = buf_xcpt_if ? bufMask : 2'h0;
  assign T_459 = ~ bufMask;
  assign T_461 = io_imem_bits_xcpt_if ? T_459 : 2'h0;
  assign T_462 = T_458 | T_461;
  assign xcpt_if = valid & T_462;
  assign T_464 = buf_replay ? bufMask : 2'h0;
  assign T_467 = io_imem_bits_replay ? T_459 : 2'h0;
  assign T_468 = T_464 | T_467;
  assign ic_replay = valid & T_468;
  assign T_470 = 2'h1 << ibufBTBResp_bridx;
  assign ibufBTBHitMask = ibufBTBHit ? T_470 : 2'h0;
  assign T_472 = io_imem_bits_btb_bits_bridx + nBufValid;
  assign T_473 = T_472 - GEN_31;
  assign T_474 = T_473[1:0];
  assign T_476 = 4'h1 << T_474;
  assign icBTBHitMask = io_imem_bits_btb_valid ? T_476 : 4'h0;
  assign T_478 = ibufBTBHitMask & bufMask;
  assign GEN_49 = {{2'd0}, T_459};
  assign T_480 = icBTBHitMask & GEN_49;
  assign GEN_50 = {{2'd0}, T_478};
  assign btbHitMask = GEN_50 | T_480;
  assign T_483 = T_478 != 2'h0;
  assign T_484_taken = T_483 ? ibufBTBResp_taken : io_imem_bits_btb_bits_taken;
  assign T_484_mask = T_483 ? ibufBTBResp_mask : io_imem_bits_btb_bits_mask;
  assign T_484_bridx = T_483 ? ibufBTBResp_bridx : io_imem_bits_btb_bits_bridx;
  assign T_484_target = T_483 ? ibufBTBResp_target : io_imem_bits_btb_bits_target;
  assign T_484_entry = T_483 ? ibufBTBResp_entry : io_imem_bits_btb_bits_entry;
  assign T_484_bht_history = T_483 ? ibufBTBResp_bht_history : io_imem_bits_btb_bits_bht_history;
  assign T_484_bht_value = T_483 ? ibufBTBResp_bht_value : io_imem_bits_btb_bits_bht_value;
  assign T_494 = nBufValid > 1'h0;
  assign T_495 = T_494 ? buf_pc : io_imem_bits_pc;
  assign RVCExpander_1_clk = clk;
  assign RVCExpander_1_reset = reset;
  assign RVCExpander_1_io_in = inst;
  assign T_497 = ic_replay >> 1'h0;
  assign T_498 = T_497[0];
  assign T_500 = RVCExpander_1_io_rvc == 1'h0;
  assign T_501 = btbHitMask >> 1'h0;
  assign T_502 = T_501[0];
  assign T_504 = 1'h0 + 1'h1;
  assign T_505 = T_504[0:0];
  assign T_506 = ic_replay >> T_505;
  assign T_507 = T_506[0];
  assign T_508 = T_502 | T_507;
  assign T_509 = T_500 & T_508;
  assign T_510 = T_498 | T_509;
  assign T_511 = valid >> 1'h0;
  assign T_512 = T_511[0];
  assign T_516 = valid >> T_505;
  assign T_517 = T_516[0];
  assign T_518 = RVCExpander_1_io_rvc | T_517;
  assign T_522 = xcpt_if >> T_505;
  assign T_523 = T_522[0];
  assign T_524 = T_518 | T_523;
  assign T_525 = T_524 | T_510;
  assign T_526 = T_512 & T_525;
  assign T_527 = xcpt_if >> 1'h0;
  assign T_528 = T_527[0];
  assign T_536 = T_500 & T_523;
  assign T_544 = btbHitMask >> T_505;
  assign T_545 = T_544[0];
  assign T_546 = T_500 & T_545;
  assign T_547 = T_502 | T_546;
  assign T_548 = io_inst_0_ready & io_inst_0_valid;
  assign T_553 = 2'h0 + 2'h2;
  assign T_554 = T_553[1:0];
  assign T_555 = RVCExpander_1_io_rvc ? {{1'd0}, T_505} : T_554;
  assign GEN_30 = T_548 ? T_555 : 2'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  nBufValid = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  buf_btb_valid = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  buf_btb_bits_taken = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  buf_btb_bits_mask = GEN_36[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  buf_btb_bits_bridx = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {2{$random}};
  buf_btb_bits_target = GEN_38[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  buf_btb_bits_entry = GEN_43[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  buf_btb_bits_bht_history = GEN_44[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  buf_btb_bits_bht_value = GEN_48[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {2{$random}};
  buf_pc = GEN_51[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  buf_data = GEN_52[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  buf_mask = GEN_53[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  buf_xcpt_if = GEN_54[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  buf_replay = GEN_55[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  ibufBTBHit = GEN_56[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  ibufBTBResp_taken = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  ibufBTBResp_mask = GEN_58[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  ibufBTBResp_bridx = GEN_59[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {2{$random}};
  ibufBTBResp_target = GEN_60[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_61 = {1{$random}};
  ibufBTBResp_entry = GEN_61[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_62 = {1{$random}};
  ibufBTBResp_bht_history = GEN_62[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_63 = {1{$random}};
  ibufBTBResp_bht_value = GEN_63[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= GEN_29[0];
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_valid <= io_imem_bits_btb_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_taken <= io_imem_bits_btb_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_mask <= io_imem_bits_btb_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bridx <= io_imem_bits_btb_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_target <= io_imem_bits_btb_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_entry <= io_imem_bits_btb_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bht_history <= io_imem_bits_btb_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_btb_bits_bht_value <= io_imem_bits_btb_bits_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_pc <= T_423;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_data <= {{16'd0}, T_416};
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_mask <= io_imem_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_xcpt_if <= io_imem_bits_xcpt_if;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        buf_replay <= io_imem_bits_replay;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        ibufBTBHit <= io_imem_bits_btb_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_taken <= io_imem_bits_btb_bits_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_mask <= io_imem_bits_btb_bits_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ibufBTBResp_bridx <= GEN_24[0];
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_target <= io_imem_bits_btb_bits_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_entry <= io_imem_bits_btb_bits_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_bht_history <= io_imem_bits_btb_bits_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_406) begin
        if(io_imem_bits_btb_valid) begin
          ibufBTBResp_bht_value <= io_imem_bits_btb_bits_bht_value;
        end
      end
    end
  end
endmodule
module CSRFile(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  input  [11:0] io_rw_addr,
  input  [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  output  io_csr_stall,
  output  io_csr_xcpt,
  output  io_eret,
  output  io_singleStep,
  output  io_status_debug,
  output [1:0] io_status_prv,
  output  io_status_sd,
  output [30:0] io_status_zero3,
  output  io_status_sd_rv32,
  output [1:0] io_status_zero2,
  output [4:0] io_status_vm,
  output [3:0] io_status_zero1,
  output  io_status_mxr,
  output  io_status_pum,
  output  io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_hpp,
  output  io_status_spp,
  output  io_status_mpie,
  output  io_status_hpie,
  output  io_status_spie,
  output  io_status_upie,
  output  io_status_mie,
  output  io_status_hie,
  output  io_status_sie,
  output  io_status_uie,
  output [6:0] io_ptbr_asid,
  output [37:0] io_ptbr_ppn,
  output [39:0] io_evec,
  input   io_exception,
  input   io_retire,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_badaddr,
  output  io_fatc,
  output [63:0] io_time,
  output [2:0] io_fcsr_rm,
  input   io_fcsr_flags_valid,
  input  [4:0] io_fcsr_flags_bits,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [6:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [6:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [10:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output  io_interrupt,
  output [63:0] io_interrupt_cause,
  output [3:0] io_bp_0_control_ttype,
  output  io_bp_0_control_dmode,
  output [5:0] io_bp_0_control_maskmax,
  output [39:0] io_bp_0_control_reserved,
  output  io_bp_0_control_action,
  output  io_bp_0_control_chain,
  output [1:0] io_bp_0_control_zero,
  output [1:0] io_bp_0_control_tmatch,
  output  io_bp_0_control_m,
  output  io_bp_0_control_h,
  output  io_bp_0_control_s,
  output  io_bp_0_control_u,
  output  io_bp_0_control_x,
  output  io_bp_0_control_w,
  output  io_bp_0_control_r,
  output [38:0] io_bp_0_address
);
  wire  T_4982_debug;
  wire [1:0] T_4982_prv;
  wire  T_4982_sd;
  wire [30:0] T_4982_zero3;
  wire  T_4982_sd_rv32;
  wire [1:0] T_4982_zero2;
  wire [4:0] T_4982_vm;
  wire [3:0] T_4982_zero1;
  wire  T_4982_mxr;
  wire  T_4982_pum;
  wire  T_4982_mprv;
  wire [1:0] T_4982_xs;
  wire [1:0] T_4982_fs;
  wire [1:0] T_4982_mpp;
  wire [1:0] T_4982_hpp;
  wire  T_4982_spp;
  wire  T_4982_mpie;
  wire  T_4982_hpie;
  wire  T_4982_spie;
  wire  T_4982_upie;
  wire  T_4982_mie;
  wire  T_4982_hie;
  wire  T_4982_sie;
  wire  T_4982_uie;
  wire [66:0] T_5008;
  wire  T_5009;
  wire  T_5010;
  wire  T_5011;
  wire  T_5012;
  wire  T_5013;
  wire  T_5014;
  wire  T_5015;
  wire  T_5016;
  wire  T_5017;
  wire [1:0] T_5018;
  wire [1:0] T_5019;
  wire [1:0] T_5020;
  wire [1:0] T_5021;
  wire  T_5022;
  wire  T_5023;
  wire  T_5024;
  wire [3:0] T_5025;
  wire [4:0] T_5026;
  wire [1:0] T_5027;
  wire  T_5028;
  wire [30:0] T_5029;
  wire  T_5030;
  wire [1:0] T_5031;
  wire  T_5032;
  wire  reset_mstatus_debug;
  wire [1:0] reset_mstatus_prv;
  wire  reset_mstatus_sd;
  wire [30:0] reset_mstatus_zero3;
  wire  reset_mstatus_sd_rv32;
  wire [1:0] reset_mstatus_zero2;
  wire [4:0] reset_mstatus_vm;
  wire [3:0] reset_mstatus_zero1;
  wire  reset_mstatus_mxr;
  wire  reset_mstatus_pum;
  wire  reset_mstatus_mprv;
  wire [1:0] reset_mstatus_xs;
  wire [1:0] reset_mstatus_fs;
  wire [1:0] reset_mstatus_mpp;
  wire [1:0] reset_mstatus_hpp;
  wire  reset_mstatus_spp;
  wire  reset_mstatus_mpie;
  wire  reset_mstatus_hpie;
  wire  reset_mstatus_spie;
  wire  reset_mstatus_upie;
  wire  reset_mstatus_mie;
  wire  reset_mstatus_hie;
  wire  reset_mstatus_sie;
  wire  reset_mstatus_uie;
  reg  reg_mstatus_debug;
  reg [31:0] GEN_124;
  reg [1:0] reg_mstatus_prv;
  reg [31:0] GEN_125;
  reg  reg_mstatus_sd;
  reg [31:0] GEN_126;
  reg [30:0] reg_mstatus_zero3;
  reg [31:0] GEN_127;
  reg  reg_mstatus_sd_rv32;
  reg [31:0] GEN_128;
  reg [1:0] reg_mstatus_zero2;
  reg [31:0] GEN_129;
  reg [4:0] reg_mstatus_vm;
  reg [31:0] GEN_130;
  reg [3:0] reg_mstatus_zero1;
  reg [31:0] GEN_131;
  reg  reg_mstatus_mxr;
  reg [31:0] GEN_132;
  reg  reg_mstatus_pum;
  reg [31:0] GEN_133;
  reg  reg_mstatus_mprv;
  reg [31:0] GEN_134;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] GEN_135;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] GEN_136;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] GEN_137;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] GEN_138;
  reg  reg_mstatus_spp;
  reg [31:0] GEN_139;
  reg  reg_mstatus_mpie;
  reg [31:0] GEN_140;
  reg  reg_mstatus_hpie;
  reg [31:0] GEN_141;
  reg  reg_mstatus_spie;
  reg [31:0] GEN_142;
  reg  reg_mstatus_upie;
  reg [31:0] GEN_143;
  reg  reg_mstatus_mie;
  reg [31:0] GEN_144;
  reg  reg_mstatus_hie;
  reg [31:0] GEN_145;
  reg  reg_mstatus_sie;
  reg [31:0] GEN_146;
  reg  reg_mstatus_uie;
  reg [31:0] GEN_147;
  wire [1:0] new_prv;
  wire  T_5084;
  wire [1:0] T_5086;
  wire [1:0] T_5124_xdebugver;
  wire  T_5124_ndreset;
  wire  T_5124_fullreset;
  wire [11:0] T_5124_zero3;
  wire  T_5124_ebreakm;
  wire  T_5124_ebreakh;
  wire  T_5124_ebreaks;
  wire  T_5124_ebreaku;
  wire  T_5124_zero2;
  wire  T_5124_stopcycle;
  wire  T_5124_stoptime;
  wire [2:0] T_5124_cause;
  wire  T_5124_debugint;
  wire  T_5124_zero1;
  wire  T_5124_halt;
  wire  T_5124_step;
  wire [1:0] T_5124_prv;
  wire [31:0] T_5143;
  wire [1:0] T_5144;
  wire  T_5145;
  wire  T_5146;
  wire  T_5147;
  wire  T_5148;
  wire [2:0] T_5149;
  wire  T_5150;
  wire  T_5151;
  wire  T_5152;
  wire  T_5153;
  wire  T_5154;
  wire  T_5155;
  wire  T_5156;
  wire [11:0] T_5157;
  wire  T_5158;
  wire  T_5159;
  wire [1:0] T_5160;
  wire [1:0] reset_dcsr_xdebugver;
  wire  reset_dcsr_ndreset;
  wire  reset_dcsr_fullreset;
  wire [11:0] reset_dcsr_zero3;
  wire  reset_dcsr_ebreakm;
  wire  reset_dcsr_ebreakh;
  wire  reset_dcsr_ebreaks;
  wire  reset_dcsr_ebreaku;
  wire  reset_dcsr_zero2;
  wire  reset_dcsr_stopcycle;
  wire  reset_dcsr_stoptime;
  wire [2:0] reset_dcsr_cause;
  wire  reset_dcsr_debugint;
  wire  reset_dcsr_zero1;
  wire  reset_dcsr_halt;
  wire  reset_dcsr_step;
  wire [1:0] reset_dcsr_prv;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] GEN_148;
  reg  reg_dcsr_ndreset;
  reg [31:0] GEN_149;
  reg  reg_dcsr_fullreset;
  reg [31:0] GEN_150;
  reg [11:0] reg_dcsr_zero3;
  reg [31:0] GEN_151;
  reg  reg_dcsr_ebreakm;
  reg [31:0] GEN_152;
  reg  reg_dcsr_ebreakh;
  reg [31:0] GEN_153;
  reg  reg_dcsr_ebreaks;
  reg [31:0] GEN_154;
  reg  reg_dcsr_ebreaku;
  reg [31:0] GEN_155;
  reg  reg_dcsr_zero2;
  reg [31:0] GEN_156;
  reg  reg_dcsr_stopcycle;
  reg [31:0] GEN_157;
  reg  reg_dcsr_stoptime;
  reg [31:0] GEN_158;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] GEN_159;
  reg  reg_dcsr_debugint;
  reg [31:0] GEN_160;
  reg  reg_dcsr_zero1;
  reg [31:0] GEN_161;
  reg  reg_dcsr_halt;
  reg [31:0] GEN_162;
  reg  reg_dcsr_step;
  reg [31:0] GEN_163;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] GEN_164;
  wire  T_5226_rocc;
  wire  T_5226_meip;
  wire  T_5226_heip;
  wire  T_5226_seip;
  wire  T_5226_ueip;
  wire  T_5226_mtip;
  wire  T_5226_htip;
  wire  T_5226_stip;
  wire  T_5226_utip;
  wire  T_5226_msip;
  wire  T_5226_hsip;
  wire  T_5226_ssip;
  wire  T_5226_usip;
  wire [12:0] T_5241;
  wire  T_5242;
  wire  T_5243;
  wire  T_5244;
  wire  T_5245;
  wire  T_5246;
  wire  T_5247;
  wire  T_5248;
  wire  T_5249;
  wire  T_5250;
  wire  T_5251;
  wire  T_5252;
  wire  T_5253;
  wire  T_5254;
  wire  T_5255_rocc;
  wire  T_5255_meip;
  wire  T_5255_heip;
  wire  T_5255_seip;
  wire  T_5255_ueip;
  wire  T_5255_mtip;
  wire  T_5255_htip;
  wire  T_5255_stip;
  wire  T_5255_utip;
  wire  T_5255_msip;
  wire  T_5255_hsip;
  wire  T_5255_ssip;
  wire  T_5255_usip;
  wire  T_5276_rocc;
  wire  T_5276_meip;
  wire  T_5276_heip;
  wire  T_5276_seip;
  wire  T_5276_ueip;
  wire  T_5276_mtip;
  wire  T_5276_htip;
  wire  T_5276_stip;
  wire  T_5276_utip;
  wire  T_5276_msip;
  wire  T_5276_hsip;
  wire  T_5276_ssip;
  wire  T_5276_usip;
  wire [1:0] T_5293;
  wire [2:0] T_5294;
  wire [1:0] T_5295;
  wire [2:0] T_5296;
  wire [5:0] T_5297;
  wire [1:0] T_5298;
  wire [2:0] T_5299;
  wire [1:0] T_5300;
  wire [1:0] T_5301;
  wire [3:0] T_5302;
  wire [6:0] T_5303;
  wire [12:0] supported_interrupts;
  wire [1:0] T_5304;
  wire [2:0] T_5305;
  wire [1:0] T_5306;
  wire [2:0] T_5307;
  wire [5:0] T_5308;
  wire [1:0] T_5309;
  wire [2:0] T_5310;
  wire [1:0] T_5311;
  wire [1:0] T_5312;
  wire [3:0] T_5313;
  wire [6:0] T_5314;
  wire [12:0] delegable_interrupts;
  wire  exception;
  reg  reg_debug;
  reg [31:0] GEN_165;
  reg [39:0] reg_dpc;
  reg [63:0] GEN_166;
  reg [63:0] reg_dscratch;
  reg [63:0] GEN_167;
  reg  reg_singleStepped;
  reg [31:0] GEN_168;
  wire  T_5320;
  wire  GEN_36;
  wire  T_5323;
  wire  GEN_37;
  wire  T_5334;
  wire  T_5336;
  wire  T_5337;
  wire  T_5338;
  wire  T_5340;
  reg  reg_tselect;
  reg [31:0] GEN_169;
  reg [3:0] reg_bp_0_control_ttype;
  reg [31:0] GEN_170;
  reg  reg_bp_0_control_dmode;
  reg [31:0] GEN_171;
  reg [5:0] reg_bp_0_control_maskmax;
  reg [31:0] GEN_172;
  reg [39:0] reg_bp_0_control_reserved;
  reg [63:0] GEN_173;
  reg  reg_bp_0_control_action;
  reg [31:0] GEN_174;
  reg  reg_bp_0_control_chain;
  reg [31:0] GEN_175;
  reg [1:0] reg_bp_0_control_zero;
  reg [31:0] GEN_176;
  reg [1:0] reg_bp_0_control_tmatch;
  reg [31:0] GEN_177;
  reg  reg_bp_0_control_m;
  reg [31:0] GEN_178;
  reg  reg_bp_0_control_h;
  reg [31:0] GEN_179;
  reg  reg_bp_0_control_s;
  reg [31:0] GEN_180;
  reg  reg_bp_0_control_u;
  reg [31:0] GEN_181;
  reg  reg_bp_0_control_x;
  reg [31:0] GEN_182;
  reg  reg_bp_0_control_w;
  reg [31:0] GEN_183;
  reg  reg_bp_0_control_r;
  reg [31:0] GEN_184;
  reg [38:0] reg_bp_0_address;
  reg [63:0] GEN_185;
  reg [3:0] reg_bp_1_control_ttype;
  reg [31:0] GEN_186;
  reg  reg_bp_1_control_dmode;
  reg [31:0] GEN_187;
  reg [5:0] reg_bp_1_control_maskmax;
  reg [31:0] GEN_188;
  reg [39:0] reg_bp_1_control_reserved;
  reg [63:0] GEN_189;
  reg  reg_bp_1_control_action;
  reg [31:0] GEN_190;
  reg  reg_bp_1_control_chain;
  reg [31:0] GEN_191;
  reg [1:0] reg_bp_1_control_zero;
  reg [31:0] GEN_192;
  reg [1:0] reg_bp_1_control_tmatch;
  reg [31:0] GEN_193;
  reg  reg_bp_1_control_m;
  reg [31:0] GEN_194;
  reg  reg_bp_1_control_h;
  reg [31:0] GEN_195;
  reg  reg_bp_1_control_s;
  reg [31:0] GEN_196;
  reg  reg_bp_1_control_u;
  reg [31:0] GEN_197;
  reg  reg_bp_1_control_x;
  reg [31:0] GEN_198;
  reg  reg_bp_1_control_w;
  reg [31:0] GEN_199;
  reg  reg_bp_1_control_r;
  reg [31:0] GEN_200;
  reg [38:0] reg_bp_1_address;
  reg [63:0] GEN_201;
  reg [63:0] reg_mie;
  reg [63:0] GEN_202;
  reg [63:0] reg_mideleg;
  reg [63:0] GEN_203;
  reg [63:0] reg_medeleg;
  reg [63:0] GEN_204;
  reg  reg_mip_rocc;
  reg [31:0] GEN_205;
  reg  reg_mip_meip;
  reg [31:0] GEN_206;
  reg  reg_mip_heip;
  reg [31:0] GEN_207;
  reg  reg_mip_seip;
  reg [31:0] GEN_208;
  reg  reg_mip_ueip;
  reg [31:0] GEN_209;
  reg  reg_mip_mtip;
  reg [31:0] GEN_210;
  reg  reg_mip_htip;
  reg [31:0] GEN_211;
  reg  reg_mip_stip;
  reg [31:0] GEN_212;
  reg  reg_mip_utip;
  reg [31:0] GEN_213;
  reg  reg_mip_msip;
  reg [31:0] GEN_214;
  reg  reg_mip_hsip;
  reg [31:0] GEN_215;
  reg  reg_mip_ssip;
  reg [31:0] GEN_216;
  reg  reg_mip_usip;
  reg [31:0] GEN_217;
  reg [39:0] reg_mepc;
  reg [63:0] GEN_218;
  reg [63:0] reg_mcause;
  reg [63:0] GEN_219;
  reg [39:0] reg_mbadaddr;
  reg [63:0] GEN_220;
  reg [63:0] reg_mscratch;
  reg [63:0] GEN_221;
  reg [31:0] reg_mtvec;
  reg [31:0] GEN_222;
  reg [31:0] reg_mucounteren;
  reg [31:0] GEN_223;
  reg [31:0] reg_mscounteren;
  reg [31:0] GEN_224;
  reg [39:0] reg_sepc;
  reg [63:0] GEN_225;
  reg [63:0] reg_scause;
  reg [63:0] GEN_226;
  reg [39:0] reg_sbadaddr;
  reg [63:0] GEN_227;
  reg [63:0] reg_sscratch;
  reg [63:0] GEN_228;
  reg [38:0] reg_stvec;
  reg [63:0] GEN_229;
  reg [6:0] reg_sptbr_asid;
  reg [31:0] GEN_230;
  reg [37:0] reg_sptbr_ppn;
  reg [63:0] GEN_231;
  reg  reg_wfi;
  reg [31:0] GEN_232;
  reg [4:0] reg_fflags;
  reg [31:0] GEN_233;
  reg [2:0] reg_frm;
  reg [31:0] GEN_234;
  reg [5:0] T_5570;
  reg [31:0] GEN_235;
  wire [5:0] GEN_0;
  wire [6:0] T_5571;
  reg [57:0] T_5573;
  reg [63:0] GEN_236;
  wire  T_5574;
  wire [58:0] T_5576;
  wire [57:0] T_5577;
  wire [57:0] GEN_38;
  wire [63:0] T_5578;
  reg [5:0] T_5581;
  reg [31:0] GEN_237;
  wire [6:0] T_5582;
  reg [57:0] T_5584;
  reg [63:0] GEN_238;
  wire  T_5585;
  wire [58:0] T_5587;
  wire [57:0] T_5588;
  wire [57:0] GEN_39;
  wire [63:0] T_5589;
  wire  mip_rocc;
  wire  mip_meip;
  wire  mip_heip;
  wire  mip_seip;
  wire  mip_ueip;
  wire  mip_mtip;
  wire  mip_htip;
  wire  mip_stip;
  wire  mip_utip;
  wire  mip_msip;
  wire  mip_hsip;
  wire  mip_ssip;
  wire  mip_usip;
  wire [1:0] T_5603;
  wire [2:0] T_5604;
  wire [1:0] T_5605;
  wire [2:0] T_5606;
  wire [5:0] T_5607;
  wire [1:0] T_5608;
  wire [2:0] T_5609;
  wire [1:0] T_5610;
  wire [1:0] T_5611;
  wire [3:0] T_5612;
  wire [6:0] T_5613;
  wire [12:0] T_5614;
  wire [12:0] read_mip;
  wire [63:0] GEN_1;
  wire [63:0] pending_interrupts;
  wire  T_5616;
  wire  T_5618;
  wire  T_5620;
  wire  T_5621;
  wire  T_5622;
  wire  T_5623;
  wire [63:0] T_5624;
  wire [63:0] T_5625;
  wire [63:0] m_interrupts;
  wire  T_5630;
  wire  T_5632;
  wire  T_5633;
  wire  T_5634;
  wire  T_5635;
  wire [63:0] T_5636;
  wire [63:0] s_interrupts;
  wire [63:0] all_interrupts;
  wire  T_5639;
  wire  T_5640;
  wire  T_5641;
  wire  T_5642;
  wire  T_5643;
  wire  T_5644;
  wire  T_5645;
  wire  T_5646;
  wire  T_5647;
  wire  T_5648;
  wire  T_5649;
  wire  T_5650;
  wire  T_5651;
  wire  T_5652;
  wire  T_5653;
  wire  T_5654;
  wire  T_5655;
  wire  T_5656;
  wire  T_5657;
  wire  T_5658;
  wire  T_5659;
  wire  T_5660;
  wire  T_5661;
  wire  T_5662;
  wire  T_5663;
  wire  T_5664;
  wire  T_5665;
  wire  T_5666;
  wire  T_5667;
  wire  T_5668;
  wire  T_5669;
  wire  T_5670;
  wire  T_5671;
  wire  T_5672;
  wire  T_5673;
  wire  T_5674;
  wire  T_5675;
  wire  T_5676;
  wire  T_5677;
  wire  T_5678;
  wire  T_5679;
  wire  T_5680;
  wire  T_5681;
  wire  T_5682;
  wire  T_5683;
  wire  T_5684;
  wire  T_5685;
  wire  T_5686;
  wire  T_5687;
  wire  T_5688;
  wire  T_5689;
  wire  T_5690;
  wire  T_5691;
  wire  T_5692;
  wire  T_5693;
  wire  T_5694;
  wire  T_5695;
  wire  T_5696;
  wire  T_5697;
  wire  T_5698;
  wire  T_5699;
  wire  T_5700;
  wire  T_5701;
  wire [5:0] T_5767;
  wire [5:0] T_5768;
  wire [5:0] T_5769;
  wire [5:0] T_5770;
  wire [5:0] T_5771;
  wire [5:0] T_5772;
  wire [5:0] T_5773;
  wire [5:0] T_5774;
  wire [5:0] T_5775;
  wire [5:0] T_5776;
  wire [5:0] T_5777;
  wire [5:0] T_5778;
  wire [5:0] T_5779;
  wire [5:0] T_5780;
  wire [5:0] T_5781;
  wire [5:0] T_5782;
  wire [5:0] T_5783;
  wire [5:0] T_5784;
  wire [5:0] T_5785;
  wire [5:0] T_5786;
  wire [5:0] T_5787;
  wire [5:0] T_5788;
  wire [5:0] T_5789;
  wire [5:0] T_5790;
  wire [5:0] T_5791;
  wire [5:0] T_5792;
  wire [5:0] T_5793;
  wire [5:0] T_5794;
  wire [5:0] T_5795;
  wire [5:0] T_5796;
  wire [5:0] T_5797;
  wire [5:0] T_5798;
  wire [5:0] T_5799;
  wire [5:0] T_5800;
  wire [5:0] T_5801;
  wire [5:0] T_5802;
  wire [5:0] T_5803;
  wire [5:0] T_5804;
  wire [5:0] T_5805;
  wire [5:0] T_5806;
  wire [5:0] T_5807;
  wire [5:0] T_5808;
  wire [5:0] T_5809;
  wire [5:0] T_5810;
  wire [5:0] T_5811;
  wire [5:0] T_5812;
  wire [5:0] T_5813;
  wire [5:0] T_5814;
  wire [5:0] T_5815;
  wire [5:0] T_5816;
  wire [5:0] T_5817;
  wire [5:0] T_5818;
  wire [5:0] T_5819;
  wire [5:0] T_5820;
  wire [5:0] T_5821;
  wire [5:0] T_5822;
  wire [5:0] T_5823;
  wire [5:0] T_5824;
  wire [5:0] T_5825;
  wire [5:0] T_5826;
  wire [5:0] T_5827;
  wire [5:0] T_5828;
  wire [5:0] T_5829;
  wire [63:0] GEN_2;
  wire [64:0] T_5830;
  wire [63:0] interruptCause;
  wire  T_5832;
  wire  T_5835;
  wire  T_5836;
  wire  T_5841;
  wire  GEN_40;
  wire [63:0] GEN_41;
  wire  system_insn;
  wire  T_5844;
  wire  T_5846;
  wire  cpu_ren;
  wire  T_5847;
  wire  cpu_wen;
  wire [1:0] T_5848;
  wire [2:0] T_5849;
  wire [1:0] T_5850;
  wire [2:0] T_5851;
  wire [5:0] T_5852;
  wire [1:0] T_5853;
  wire [2:0] T_5854;
  wire [3:0] T_5855;
  wire [5:0] T_5856;
  wire [8:0] T_5857;
  wire [14:0] T_5858;
  wire [1:0] T_5859;
  wire [3:0] T_5860;
  wire [8:0] T_5861;
  wire [9:0] T_5862;
  wire [13:0] T_5863;
  wire [31:0] T_5864;
  wire [33:0] T_5865;
  wire [2:0] T_5866;
  wire [3:0] T_5867;
  wire [37:0] T_5868;
  wire [51:0] T_5869;
  wire [66:0] T_5870;
  wire [63:0] read_mstatus;
  wire [3:0] GEN_0_control_ttype;
  wire  GEN_0_control_dmode;
  wire [5:0] GEN_0_control_maskmax;
  wire [39:0] GEN_0_control_reserved;
  wire  GEN_0_control_action;
  wire  GEN_0_control_chain;
  wire [1:0] GEN_0_control_zero;
  wire [1:0] GEN_0_control_tmatch;
  wire  GEN_0_control_m;
  wire  GEN_0_control_h;
  wire  GEN_0_control_s;
  wire  GEN_0_control_u;
  wire  GEN_0_control_x;
  wire  GEN_0_control_w;
  wire  GEN_0_control_r;
  wire [38:0] GEN_0_address;
  wire [3:0] GEN_42;
  wire  GEN_43;
  wire [5:0] GEN_44;
  wire [39:0] GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire [1:0] GEN_48;
  wire [1:0] GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire [38:0] GEN_57;
  wire [3:0] GEN_1_control_ttype;
  wire  GEN_1_control_dmode;
  wire [5:0] GEN_1_control_maskmax;
  wire [39:0] GEN_1_control_reserved;
  wire  GEN_1_control_action;
  wire  GEN_1_control_chain;
  wire [1:0] GEN_1_control_zero;
  wire [1:0] GEN_1_control_tmatch;
  wire  GEN_1_control_m;
  wire  GEN_1_control_h;
  wire  GEN_1_control_s;
  wire  GEN_1_control_u;
  wire  GEN_1_control_x;
  wire  GEN_1_control_w;
  wire  GEN_1_control_r;
  wire [38:0] GEN_1_address;
  wire [1:0] T_5888;
  wire [3:0] GEN_2_control_ttype;
  wire  GEN_2_control_dmode;
  wire [5:0] GEN_2_control_maskmax;
  wire [39:0] GEN_2_control_reserved;
  wire  GEN_2_control_action;
  wire  GEN_2_control_chain;
  wire [1:0] GEN_2_control_zero;
  wire [1:0] GEN_2_control_tmatch;
  wire  GEN_2_control_m;
  wire  GEN_2_control_h;
  wire  GEN_2_control_s;
  wire  GEN_2_control_u;
  wire  GEN_2_control_x;
  wire  GEN_2_control_w;
  wire  GEN_2_control_r;
  wire [38:0] GEN_2_address;
  wire [2:0] T_5889;
  wire [3:0] GEN_3_control_ttype;
  wire  GEN_3_control_dmode;
  wire [5:0] GEN_3_control_maskmax;
  wire [39:0] GEN_3_control_reserved;
  wire  GEN_3_control_action;
  wire  GEN_3_control_chain;
  wire [1:0] GEN_3_control_zero;
  wire [1:0] GEN_3_control_tmatch;
  wire  GEN_3_control_m;
  wire  GEN_3_control_h;
  wire  GEN_3_control_s;
  wire  GEN_3_control_u;
  wire  GEN_3_control_x;
  wire  GEN_3_control_w;
  wire  GEN_3_control_r;
  wire [38:0] GEN_3_address;
  wire [3:0] GEN_4_control_ttype;
  wire  GEN_4_control_dmode;
  wire [5:0] GEN_4_control_maskmax;
  wire [39:0] GEN_4_control_reserved;
  wire  GEN_4_control_action;
  wire  GEN_4_control_chain;
  wire [1:0] GEN_4_control_zero;
  wire [1:0] GEN_4_control_tmatch;
  wire  GEN_4_control_m;
  wire  GEN_4_control_h;
  wire  GEN_4_control_s;
  wire  GEN_4_control_u;
  wire  GEN_4_control_x;
  wire  GEN_4_control_w;
  wire  GEN_4_control_r;
  wire [38:0] GEN_4_address;
  wire [1:0] T_5890;
  wire [3:0] GEN_5_control_ttype;
  wire  GEN_5_control_dmode;
  wire [5:0] GEN_5_control_maskmax;
  wire [39:0] GEN_5_control_reserved;
  wire  GEN_5_control_action;
  wire  GEN_5_control_chain;
  wire [1:0] GEN_5_control_zero;
  wire [1:0] GEN_5_control_tmatch;
  wire  GEN_5_control_m;
  wire  GEN_5_control_h;
  wire  GEN_5_control_s;
  wire  GEN_5_control_u;
  wire  GEN_5_control_x;
  wire  GEN_5_control_w;
  wire  GEN_5_control_r;
  wire [38:0] GEN_5_address;
  wire [3:0] GEN_6_control_ttype;
  wire  GEN_6_control_dmode;
  wire [5:0] GEN_6_control_maskmax;
  wire [39:0] GEN_6_control_reserved;
  wire  GEN_6_control_action;
  wire  GEN_6_control_chain;
  wire [1:0] GEN_6_control_zero;
  wire [1:0] GEN_6_control_tmatch;
  wire  GEN_6_control_m;
  wire  GEN_6_control_h;
  wire  GEN_6_control_s;
  wire  GEN_6_control_u;
  wire  GEN_6_control_x;
  wire  GEN_6_control_w;
  wire  GEN_6_control_r;
  wire [38:0] GEN_6_address;
  wire [1:0] T_5891;
  wire [3:0] T_5892;
  wire [6:0] T_5893;
  wire [3:0] GEN_7_control_ttype;
  wire  GEN_7_control_dmode;
  wire [5:0] GEN_7_control_maskmax;
  wire [39:0] GEN_7_control_reserved;
  wire  GEN_7_control_action;
  wire  GEN_7_control_chain;
  wire [1:0] GEN_7_control_zero;
  wire [1:0] GEN_7_control_tmatch;
  wire  GEN_7_control_m;
  wire  GEN_7_control_h;
  wire  GEN_7_control_s;
  wire  GEN_7_control_u;
  wire  GEN_7_control_x;
  wire  GEN_7_control_w;
  wire  GEN_7_control_r;
  wire [38:0] GEN_7_address;
  wire [3:0] GEN_8_control_ttype;
  wire  GEN_8_control_dmode;
  wire [5:0] GEN_8_control_maskmax;
  wire [39:0] GEN_8_control_reserved;
  wire  GEN_8_control_action;
  wire  GEN_8_control_chain;
  wire [1:0] GEN_8_control_zero;
  wire [1:0] GEN_8_control_tmatch;
  wire  GEN_8_control_m;
  wire  GEN_8_control_h;
  wire  GEN_8_control_s;
  wire  GEN_8_control_u;
  wire  GEN_8_control_x;
  wire  GEN_8_control_w;
  wire  GEN_8_control_r;
  wire [38:0] GEN_8_address;
  wire [3:0] T_5894;
  wire [3:0] GEN_9_control_ttype;
  wire  GEN_9_control_dmode;
  wire [5:0] GEN_9_control_maskmax;
  wire [39:0] GEN_9_control_reserved;
  wire  GEN_9_control_action;
  wire  GEN_9_control_chain;
  wire [1:0] GEN_9_control_zero;
  wire [1:0] GEN_9_control_tmatch;
  wire  GEN_9_control_m;
  wire  GEN_9_control_h;
  wire  GEN_9_control_s;
  wire  GEN_9_control_u;
  wire  GEN_9_control_x;
  wire  GEN_9_control_w;
  wire  GEN_9_control_r;
  wire [38:0] GEN_9_address;
  wire [3:0] GEN_10_control_ttype;
  wire  GEN_10_control_dmode;
  wire [5:0] GEN_10_control_maskmax;
  wire [39:0] GEN_10_control_reserved;
  wire  GEN_10_control_action;
  wire  GEN_10_control_chain;
  wire [1:0] GEN_10_control_zero;
  wire [1:0] GEN_10_control_tmatch;
  wire  GEN_10_control_m;
  wire  GEN_10_control_h;
  wire  GEN_10_control_s;
  wire  GEN_10_control_u;
  wire  GEN_10_control_x;
  wire  GEN_10_control_w;
  wire  GEN_10_control_r;
  wire [38:0] GEN_10_address;
  wire [1:0] T_5895;
  wire [5:0] T_5896;
  wire [3:0] GEN_11_control_ttype;
  wire  GEN_11_control_dmode;
  wire [5:0] GEN_11_control_maskmax;
  wire [39:0] GEN_11_control_reserved;
  wire  GEN_11_control_action;
  wire  GEN_11_control_chain;
  wire [1:0] GEN_11_control_zero;
  wire [1:0] GEN_11_control_tmatch;
  wire  GEN_11_control_m;
  wire  GEN_11_control_h;
  wire  GEN_11_control_s;
  wire  GEN_11_control_u;
  wire  GEN_11_control_x;
  wire  GEN_11_control_w;
  wire  GEN_11_control_r;
  wire [38:0] GEN_11_address;
  wire [3:0] GEN_12_control_ttype;
  wire  GEN_12_control_dmode;
  wire [5:0] GEN_12_control_maskmax;
  wire [39:0] GEN_12_control_reserved;
  wire  GEN_12_control_action;
  wire  GEN_12_control_chain;
  wire [1:0] GEN_12_control_zero;
  wire [1:0] GEN_12_control_tmatch;
  wire  GEN_12_control_m;
  wire  GEN_12_control_h;
  wire  GEN_12_control_s;
  wire  GEN_12_control_u;
  wire  GEN_12_control_x;
  wire  GEN_12_control_w;
  wire  GEN_12_control_r;
  wire [38:0] GEN_12_address;
  wire [45:0] T_5897;
  wire [3:0] GEN_13_control_ttype;
  wire  GEN_13_control_dmode;
  wire [5:0] GEN_13_control_maskmax;
  wire [39:0] GEN_13_control_reserved;
  wire  GEN_13_control_action;
  wire  GEN_13_control_chain;
  wire [1:0] GEN_13_control_zero;
  wire [1:0] GEN_13_control_tmatch;
  wire  GEN_13_control_m;
  wire  GEN_13_control_h;
  wire  GEN_13_control_s;
  wire  GEN_13_control_u;
  wire  GEN_13_control_x;
  wire  GEN_13_control_w;
  wire  GEN_13_control_r;
  wire [38:0] GEN_13_address;
  wire [3:0] GEN_14_control_ttype;
  wire  GEN_14_control_dmode;
  wire [5:0] GEN_14_control_maskmax;
  wire [39:0] GEN_14_control_reserved;
  wire  GEN_14_control_action;
  wire  GEN_14_control_chain;
  wire [1:0] GEN_14_control_zero;
  wire [1:0] GEN_14_control_tmatch;
  wire  GEN_14_control_m;
  wire  GEN_14_control_h;
  wire  GEN_14_control_s;
  wire  GEN_14_control_u;
  wire  GEN_14_control_x;
  wire  GEN_14_control_w;
  wire  GEN_14_control_r;
  wire [38:0] GEN_14_address;
  wire [4:0] T_5898;
  wire [50:0] T_5899;
  wire [56:0] T_5900;
  wire [63:0] T_5901;
  wire [3:0] GEN_15_control_ttype;
  wire  GEN_15_control_dmode;
  wire [5:0] GEN_15_control_maskmax;
  wire [39:0] GEN_15_control_reserved;
  wire  GEN_15_control_action;
  wire  GEN_15_control_chain;
  wire [1:0] GEN_15_control_zero;
  wire [1:0] GEN_15_control_tmatch;
  wire  GEN_15_control_m;
  wire  GEN_15_control_h;
  wire  GEN_15_control_s;
  wire  GEN_15_control_u;
  wire  GEN_15_control_x;
  wire  GEN_15_control_w;
  wire  GEN_15_control_r;
  wire [38:0] GEN_15_address;
  wire  T_5919;
  wire [24:0] T_5923;
  wire [3:0] GEN_16_control_ttype;
  wire  GEN_16_control_dmode;
  wire [5:0] GEN_16_control_maskmax;
  wire [39:0] GEN_16_control_reserved;
  wire  GEN_16_control_action;
  wire  GEN_16_control_chain;
  wire [1:0] GEN_16_control_zero;
  wire [1:0] GEN_16_control_tmatch;
  wire  GEN_16_control_m;
  wire  GEN_16_control_h;
  wire  GEN_16_control_s;
  wire  GEN_16_control_u;
  wire  GEN_16_control_x;
  wire  GEN_16_control_w;
  wire  GEN_16_control_r;
  wire [38:0] GEN_16_address;
  wire [63:0] T_5924;
  wire  T_5929;
  wire [23:0] T_5933;
  wire [63:0] T_5934;
  wire  T_5935;
  wire [23:0] T_5939;
  wire [63:0] T_5940;
  wire [2:0] T_5941;
  wire [1:0] T_5942;
  wire [4:0] T_5943;
  wire [3:0] T_5944;
  wire [1:0] T_5945;
  wire [5:0] T_5946;
  wire [10:0] T_5947;
  wire [1:0] T_5948;
  wire [1:0] T_5949;
  wire [3:0] T_5950;
  wire [12:0] T_5951;
  wire [2:0] T_5952;
  wire [3:0] T_5953;
  wire [16:0] T_5954;
  wire [20:0] T_5955;
  wire [31:0] T_5956;
  wire [7:0] T_5957;
  wire [63:0] T_5960;
  wire [63:0] T_5961;
  wire  T_5962_debug;
  wire [1:0] T_5962_prv;
  wire  T_5962_sd;
  wire [30:0] T_5962_zero3;
  wire  T_5962_sd_rv32;
  wire [1:0] T_5962_zero2;
  wire [4:0] T_5962_vm;
  wire [3:0] T_5962_zero1;
  wire  T_5962_mxr;
  wire  T_5962_pum;
  wire  T_5962_mprv;
  wire [1:0] T_5962_xs;
  wire [1:0] T_5962_fs;
  wire [1:0] T_5962_mpp;
  wire [1:0] T_5962_hpp;
  wire  T_5962_spp;
  wire  T_5962_mpie;
  wire  T_5962_hpie;
  wire  T_5962_spie;
  wire  T_5962_upie;
  wire  T_5962_mie;
  wire  T_5962_hie;
  wire  T_5962_sie;
  wire  T_5962_uie;
  wire [1:0] T_5995;
  wire [2:0] T_5996;
  wire [1:0] T_5997;
  wire [2:0] T_5998;
  wire [5:0] T_5999;
  wire [1:0] T_6000;
  wire [2:0] T_6001;
  wire [3:0] T_6002;
  wire [5:0] T_6003;
  wire [8:0] T_6004;
  wire [14:0] T_6005;
  wire [1:0] T_6006;
  wire [3:0] T_6007;
  wire [8:0] T_6008;
  wire [9:0] T_6009;
  wire [13:0] T_6010;
  wire [31:0] T_6011;
  wire [33:0] T_6012;
  wire [2:0] T_6013;
  wire [3:0] T_6014;
  wire [37:0] T_6015;
  wire [51:0] T_6016;
  wire [66:0] T_6017;
  wire [63:0] T_6018;
  wire  T_6019;
  wire [23:0] T_6023;
  wire [63:0] T_6024;
  wire [44:0] T_6025;
  wire  T_6026;
  wire [23:0] T_6030;
  wire [63:0] T_6031;
  wire  T_6032;
  wire [24:0] T_6036;
  wire [63:0] T_6037;
  wire  T_6039;
  wire  T_6041;
  wire  T_6043;
  wire  T_6045;
  wire  T_6047;
  wire  T_6049;
  wire  T_6051;
  wire  T_6053;
  wire  T_6055;
  wire  T_6057;
  wire  T_6059;
  wire  T_6061;
  wire  T_6063;
  wire  T_6065;
  wire  T_6067;
  wire  T_6069;
  wire  T_6071;
  wire  T_6073;
  wire  T_6075;
  wire  T_6077;
  wire  T_6079;
  wire  T_6081;
  wire  T_6083;
  wire  T_6085;
  wire  T_6087;
  wire  T_6089;
  wire  T_6091;
  wire  T_6093;
  wire  T_6095;
  wire  T_6097;
  wire  T_6099;
  wire  T_6101;
  wire  T_6103;
  wire  T_6105;
  wire  T_6107;
  wire  T_6109;
  wire  T_6111;
  wire  T_6113;
  wire  T_6115;
  wire  T_6117;
  wire  T_6119;
  wire  T_6121;
  wire  T_6123;
  wire  T_6125;
  wire  T_6127;
  wire  T_6129;
  wire  T_6131;
  wire  T_6133;
  wire  T_6135;
  wire  T_6137;
  wire  T_6139;
  wire  T_6141;
  wire  T_6143;
  wire  T_6145;
  wire  T_6147;
  wire  T_6149;
  wire  T_6151;
  wire  T_6153;
  wire  T_6155;
  wire  T_6157;
  wire  T_6159;
  wire  T_6161;
  wire  T_6163;
  wire  T_6165;
  wire  T_6167;
  wire  T_6169;
  wire  T_6171;
  wire  T_6173;
  wire  T_6175;
  wire  T_6177;
  wire  T_6179;
  wire  T_6181;
  wire  T_6183;
  wire  T_6185;
  wire  T_6187;
  wire  T_6189;
  wire  T_6191;
  wire  T_6193;
  wire  T_6195;
  wire  T_6197;
  wire  T_6199;
  wire  T_6201;
  wire  T_6203;
  wire  T_6205;
  wire  T_6207;
  wire  T_6209;
  wire  T_6211;
  wire  T_6213;
  wire  T_6215;
  wire  T_6217;
  wire  T_6219;
  wire  T_6221;
  wire  T_6223;
  wire  T_6225;
  wire  T_6227;
  wire  T_6229;
  wire  T_6231;
  wire  T_6233;
  wire  T_6235;
  wire  T_6237;
  wire  T_6239;
  wire  T_6241;
  wire  T_6243;
  wire  T_6245;
  wire  T_6247;
  wire  T_6249;
  wire  T_6251;
  wire  T_6253;
  wire  T_6255;
  wire  T_6257;
  wire  T_6259;
  wire  T_6261;
  wire  T_6263;
  wire  T_6265;
  wire  T_6267;
  wire  T_6269;
  wire  T_6271;
  wire  T_6273;
  wire  T_6275;
  wire  T_6277;
  wire  T_6279;
  wire  T_6281;
  wire  T_6283;
  wire  T_6285;
  wire  T_6287;
  wire  T_6289;
  wire  T_6290;
  wire  T_6291;
  wire  T_6292;
  wire  T_6293;
  wire  T_6294;
  wire  T_6295;
  wire  T_6296;
  wire  T_6297;
  wire  T_6298;
  wire  T_6299;
  wire  T_6300;
  wire  T_6301;
  wire  T_6302;
  wire  T_6303;
  wire  T_6304;
  wire  T_6305;
  wire  T_6306;
  wire  T_6307;
  wire  T_6308;
  wire  T_6309;
  wire  T_6310;
  wire  T_6311;
  wire  T_6312;
  wire  T_6313;
  wire  T_6314;
  wire  T_6315;
  wire  T_6316;
  wire  T_6317;
  wire  T_6318;
  wire  T_6319;
  wire  T_6320;
  wire  T_6321;
  wire  T_6322;
  wire  T_6323;
  wire  T_6324;
  wire  T_6325;
  wire  T_6326;
  wire  T_6327;
  wire  T_6328;
  wire  T_6329;
  wire  T_6330;
  wire  T_6331;
  wire  T_6332;
  wire  T_6333;
  wire  T_6334;
  wire  T_6335;
  wire  T_6336;
  wire  T_6337;
  wire  T_6338;
  wire  T_6339;
  wire  T_6340;
  wire  T_6341;
  wire  T_6342;
  wire  T_6343;
  wire  T_6344;
  wire  T_6345;
  wire  T_6346;
  wire  T_6347;
  wire  T_6348;
  wire  T_6349;
  wire  T_6350;
  wire  T_6351;
  wire  T_6352;
  wire  T_6353;
  wire  T_6354;
  wire  T_6355;
  wire  T_6356;
  wire  T_6357;
  wire  T_6358;
  wire  T_6359;
  wire  T_6360;
  wire  T_6361;
  wire  T_6362;
  wire  T_6363;
  wire  T_6364;
  wire  T_6365;
  wire  T_6366;
  wire  T_6367;
  wire  T_6368;
  wire  T_6369;
  wire  T_6370;
  wire  T_6371;
  wire  T_6372;
  wire  T_6373;
  wire  T_6374;
  wire  T_6375;
  wire  T_6376;
  wire  T_6377;
  wire  T_6378;
  wire  T_6379;
  wire  T_6380;
  wire  T_6381;
  wire  T_6382;
  wire  T_6383;
  wire  T_6384;
  wire  T_6385;
  wire  T_6386;
  wire  T_6387;
  wire  T_6388;
  wire  T_6389;
  wire  T_6390;
  wire  T_6391;
  wire  T_6392;
  wire  T_6393;
  wire  T_6394;
  wire  T_6395;
  wire  T_6396;
  wire  T_6397;
  wire  T_6398;
  wire  T_6399;
  wire  T_6400;
  wire  T_6401;
  wire  T_6402;
  wire  T_6403;
  wire  T_6404;
  wire  T_6405;
  wire  T_6406;
  wire  T_6407;
  wire  T_6408;
  wire  T_6409;
  wire  T_6410;
  wire  T_6411;
  wire  T_6412;
  wire  T_6413;
  wire  addr_valid;
  wire  T_6414;
  wire  fp_csr;
  wire  T_6416;
  wire  T_6418;
  wire  hpm_csr;
  wire  T_6421;
  wire [4:0] T_6424;
  wire [31:0] T_6425;
  wire  T_6426;
  wire  T_6427;
  wire  T_6428;
  wire  T_6430;
  wire [31:0] T_6432;
  wire  T_6433;
  wire  T_6434;
  wire  hpm_en;
  wire [1:0] csr_addr_priv;
  wire [11:0] T_6437;
  wire  T_6439;
  wire  T_6441;
  wire  T_6442;
  wire  T_6443;
  wire  priv_sufficient;
  wire [1:0] T_6444;
  wire [1:0] T_6445;
  wire  read_only;
  wire  T_6447;
  wire  T_6449;
  wire  wen;
  wire  T_6450;
  wire  T_6451;
  wire  T_6452;
  wire [63:0] T_6454;
  wire  T_6455;
  wire [63:0] T_6457;
  wire [63:0] T_6458;
  wire [63:0] T_6461;
  wire [63:0] T_6462;
  wire [63:0] wdata;
  wire  do_system_insn;
  wire [2:0] T_6464;
  wire [7:0] opcode;
  wire  T_6465;
  wire  insn_call;
  wire  T_6466;
  wire  insn_break;
  wire  T_6467;
  wire  insn_ret;
  wire  T_6468;
  wire  insn_sfence_vm;
  wire  T_6469;
  wire  insn_wfi;
  wire  T_6470;
  wire  T_6472;
  wire  T_6474;
  wire  T_6475;
  wire  T_6477;
  wire  T_6478;
  wire  T_6479;
  wire  T_6481;
  wire  T_6483;
  wire  T_6484;
  wire  T_6485;
  wire  T_6486;
  wire  T_6487;
  wire  T_6490;
  wire  T_6491;
  wire  T_6492;
  wire  T_6493;
  wire  GEN_314;
  wire  T_6496;
  wire  GEN_315;
  wire  T_6499;
  wire [3:0] GEN_4;
  wire [4:0] T_6501;
  wire [3:0] T_6502;
  wire [1:0] T_6505;
  wire [3:0] T_6506;
  wire [63:0] cause;
  wire [5:0] cause_lsbs;
  wire  T_6507;
  wire  T_6509;
  wire  causeIsDebugInt;
  wire  T_6512;
  wire  causeIsDebugTrigger;
  wire  T_6518;
  wire [1:0] T_6519;
  wire [1:0] T_6520;
  wire [3:0] T_6521;
  wire [3:0] T_6522;
  wire  T_6523;
  wire  causeIsDebugBreak;
  wire  T_6525;
  wire  T_6526;
  wire  T_6527;
  wire  T_6528;
  wire [63:0] T_6534;
  wire  T_6535;
  wire [63:0] T_6536;
  wire  T_6537;
  wire  T_6538;
  wire  delegate;
  wire [11:0] debugTVec;
  wire [39:0] T_6542;
  wire [39:0] T_6543;
  wire [39:0] tvec;
  wire  T_6545;
  wire  T_6547;
  wire [39:0] T_6549;
  wire [39:0] epc;
  wire [39:0] T_6550;
  wire  T_6553;
  wire [1:0] T_6554;
  wire  T_6556;
  wire [1:0] T_6557;
  wire  T_6559;
  wire  T_6560;
  wire [39:0] T_6561;
  wire [39:0] T_6563;
  wire [39:0] T_6564;
  wire [63:0] T_6565;
  wire  T_6566;
  wire  T_6574;
  wire  T_6575;
  wire  T_6576;
  wire  T_6577;
  wire  T_6578;
  wire  T_6579;
  wire  T_6580;
  wire  T_6581;
  wire  T_6582;
  wire  T_6583;
  wire  T_6584;
  wire  T_6585;
  wire  T_6586;
  wire [1:0] T_6592;
  wire [1:0] T_6593;
  wire [2:0] T_6594;
  wire  GEN_316;
  wire [39:0] GEN_317;
  wire [2:0] GEN_318;
  wire [1:0] GEN_319;
  wire  T_6596;
  wire  T_6597;
  wire [39:0] GEN_320;
  wire [39:0] GEN_321;
  wire [63:0] GEN_322;
  wire [39:0] GEN_323;
  wire  GEN_324;
  wire [1:0] GEN_325;
  wire  GEN_326;
  wire [1:0] GEN_327;
  wire  T_6603;
  wire  T_6604;
  wire [39:0] GEN_328;
  wire [39:0] GEN_329;
  wire [63:0] GEN_330;
  wire [39:0] GEN_331;
  wire  GEN_332;
  wire [1:0] GEN_333;
  wire  GEN_334;
  wire [1:0] GEN_335;
  wire  GEN_336;
  wire [39:0] GEN_337;
  wire [2:0] GEN_338;
  wire [1:0] GEN_339;
  wire [39:0] GEN_340;
  wire [63:0] GEN_341;
  wire [39:0] GEN_342;
  wire  GEN_343;
  wire [1:0] GEN_344;
  wire  GEN_345;
  wire [1:0] GEN_346;
  wire [39:0] GEN_347;
  wire [63:0] GEN_348;
  wire [39:0] GEN_349;
  wire  GEN_350;
  wire [1:0] GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire [1:0] GEN_356;
  wire [1:0] GEN_357;
  wire  T_6616;
  wire  T_6617;
  wire [1:0] GEN_358;
  wire  GEN_359;
  wire  T_6623;
  wire  T_6624;
  wire  GEN_360;
  wire  T_6626;
  wire  T_6629;
  wire  T_6630;
  wire  GEN_361;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire [1:0] GEN_365;
  wire [1:0] GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire [1:0] GEN_369;
  wire [1:0] GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire [1:0] GEN_374;
  wire [1:0] T_6637;
  wire [1:0] GEN_5;
  wire [2:0] T_6638;
  wire  T_6640;
  wire  T_6641;
  wire  T_6643;
  wire  T_6645;
  wire [63:0] T_6647;
  wire [63:0] T_6649;
  wire [63:0] T_6657;
  wire [63:0] T_6659;
  wire [63:0] T_6661;
  wire [63:0] T_6663;
  wire [31:0] T_6665;
  wire [12:0] T_6667;
  wire [63:0] T_6669;
  wire [63:0] T_6671;
  wire [63:0] T_6673;
  wire [63:0] T_6675;
  wire [63:0] T_6677;
  wire [63:0] T_6679;
  wire [63:0] T_6681;
  wire  T_6683;
  wire [31:0] T_6685;
  wire [39:0] T_6687;
  wire [63:0] T_6689;
  wire [4:0] T_6691;
  wire [2:0] T_6693;
  wire [7:0] T_6695;
  wire [63:0] T_6871;
  wire [63:0] T_6873;
  wire [63:0] T_6875;
  wire [63:0] T_6877;
  wire [63:0] T_6879;
  wire [63:0] T_6881;
  wire [44:0] T_6883;
  wire [63:0] T_6885;
  wire [63:0] T_6887;
  wire [31:0] T_6889;
  wire [31:0] T_6891;
  wire [63:0] T_6893;
  wire [63:0] T_6895;
  wire [63:0] GEN_6;
  wire [63:0] T_6897;
  wire [63:0] T_6898;
  wire [63:0] T_6902;
  wire [63:0] T_6903;
  wire [63:0] T_6904;
  wire [63:0] T_6905;
  wire [63:0] GEN_7;
  wire [63:0] T_6906;
  wire [63:0] GEN_8;
  wire [63:0] T_6907;
  wire [63:0] T_6908;
  wire [63:0] T_6909;
  wire [63:0] T_6910;
  wire [63:0] T_6911;
  wire [63:0] T_6912;
  wire [63:0] T_6913;
  wire [63:0] T_6914;
  wire [63:0] GEN_9;
  wire [63:0] T_6915;
  wire [63:0] GEN_10;
  wire [63:0] T_6916;
  wire [63:0] GEN_11;
  wire [63:0] T_6917;
  wire [63:0] T_6918;
  wire [63:0] GEN_12;
  wire [63:0] T_6919;
  wire [63:0] GEN_13;
  wire [63:0] T_6920;
  wire [63:0] GEN_14;
  wire [63:0] T_6921;
  wire [63:0] T_7009;
  wire [63:0] T_7010;
  wire [63:0] T_7011;
  wire [63:0] T_7012;
  wire [63:0] T_7013;
  wire [63:0] T_7014;
  wire [63:0] GEN_15;
  wire [63:0] T_7015;
  wire [63:0] T_7016;
  wire [63:0] T_7017;
  wire [63:0] GEN_16;
  wire [63:0] T_7018;
  wire [63:0] GEN_17;
  wire [63:0] T_7019;
  wire [63:0] T_7020;
  wire [63:0] T_7021;
  wire [63:0] T_7022;
  wire [4:0] T_7023;
  wire [4:0] GEN_375;
  wire  T_7074_debug;
  wire [1:0] T_7074_prv;
  wire  T_7074_sd;
  wire [30:0] T_7074_zero3;
  wire  T_7074_sd_rv32;
  wire [1:0] T_7074_zero2;
  wire [4:0] T_7074_vm;
  wire [3:0] T_7074_zero1;
  wire  T_7074_mxr;
  wire  T_7074_pum;
  wire  T_7074_mprv;
  wire [1:0] T_7074_xs;
  wire [1:0] T_7074_fs;
  wire [1:0] T_7074_mpp;
  wire [1:0] T_7074_hpp;
  wire  T_7074_spp;
  wire  T_7074_mpie;
  wire  T_7074_hpie;
  wire  T_7074_spie;
  wire  T_7074_upie;
  wire  T_7074_mie;
  wire  T_7074_hie;
  wire  T_7074_sie;
  wire  T_7074_uie;
  wire [66:0] T_7100;
  wire  T_7101;
  wire  T_7102;
  wire  T_7103;
  wire  T_7104;
  wire  T_7105;
  wire  T_7106;
  wire  T_7107;
  wire  T_7108;
  wire  T_7109;
  wire [1:0] T_7110;
  wire [1:0] T_7111;
  wire [1:0] T_7112;
  wire [1:0] T_7113;
  wire  T_7114;
  wire  T_7115;
  wire  T_7116;
  wire [3:0] T_7117;
  wire [4:0] T_7118;
  wire [1:0] T_7119;
  wire  T_7120;
  wire [30:0] T_7121;
  wire  T_7122;
  wire [1:0] T_7123;
  wire  T_7124;
  wire  T_7126;
  wire [4:0] GEN_376;
  wire  T_7129;
  wire [4:0] GEN_377;
  wire  T_7132;
  wire [1:0] T_7136;
  wire  GEN_403;
  wire  GEN_404;
  wire  GEN_405;
  wire [1:0] GEN_406;
  wire  GEN_407;
  wire  GEN_408;
  wire [1:0] GEN_409;
  wire  GEN_410;
  wire  GEN_411;
  wire [4:0] GEN_412;
  wire [1:0] GEN_413;
  wire  T_7165_rocc;
  wire  T_7165_meip;
  wire  T_7165_heip;
  wire  T_7165_seip;
  wire  T_7165_ueip;
  wire  T_7165_mtip;
  wire  T_7165_htip;
  wire  T_7165_stip;
  wire  T_7165_utip;
  wire  T_7165_msip;
  wire  T_7165_hsip;
  wire  T_7165_ssip;
  wire  T_7165_usip;
  wire  T_7179;
  wire  T_7180;
  wire  T_7181;
  wire  T_7182;
  wire  T_7183;
  wire  T_7184;
  wire  T_7185;
  wire  T_7186;
  wire  T_7187;
  wire  T_7188;
  wire  T_7189;
  wire  T_7190;
  wire  T_7191;
  wire  GEN_427;
  wire  GEN_428;
  wire [63:0] GEN_934;
  wire [63:0] T_7192;
  wire [63:0] GEN_429;
  wire [63:0] T_7193;
  wire [63:0] T_7195;
  wire [63:0] T_7196;
  wire [63:0] GEN_430;
  wire [63:0] GEN_431;
  wire [61:0] T_7197;
  wire [63:0] GEN_935;
  wire [63:0] T_7198;
  wire [63:0] GEN_432;
  wire [63:0] T_7200;
  wire [63:0] GEN_433;
  wire [39:0] T_7201;
  wire [39:0] GEN_434;
  wire [57:0] T_7202;
  wire [63:0] GEN_435;
  wire [57:0] GEN_436;
  wire [63:0] GEN_437;
  wire [57:0] GEN_438;
  wire [63:0] GEN_439;
  wire [63:0] GEN_440;
  wire [58:0] T_7204;
  wire [63:0] GEN_441;
  wire [63:0] GEN_442;
  wire [1:0] T_7241_xdebugver;
  wire  T_7241_ndreset;
  wire  T_7241_fullreset;
  wire [11:0] T_7241_zero3;
  wire  T_7241_ebreakm;
  wire  T_7241_ebreakh;
  wire  T_7241_ebreaks;
  wire  T_7241_ebreaku;
  wire  T_7241_zero2;
  wire  T_7241_stopcycle;
  wire  T_7241_stoptime;
  wire [2:0] T_7241_cause;
  wire  T_7241_debugint;
  wire  T_7241_zero1;
  wire  T_7241_halt;
  wire  T_7241_step;
  wire [1:0] T_7241_prv;
  wire [1:0] T_7259;
  wire [2:0] T_7264;
  wire  T_7269;
  wire  T_7270;
  wire  T_7271;
  wire [11:0] T_7272;
  wire  T_7273;
  wire  T_7274;
  wire [1:0] T_7275;
  wire  GEN_460;
  wire  GEN_461;
  wire  GEN_462;
  wire  GEN_463;
  wire  GEN_464;
  wire [1:0] GEN_465;
  wire [63:0] GEN_466;
  wire [63:0] GEN_467;
  wire  T_7330_debug;
  wire [1:0] T_7330_prv;
  wire  T_7330_sd;
  wire [30:0] T_7330_zero3;
  wire  T_7330_sd_rv32;
  wire [1:0] T_7330_zero2;
  wire [4:0] T_7330_vm;
  wire [3:0] T_7330_zero1;
  wire  T_7330_mxr;
  wire  T_7330_pum;
  wire  T_7330_mprv;
  wire [1:0] T_7330_xs;
  wire [1:0] T_7330_fs;
  wire [1:0] T_7330_mpp;
  wire [1:0] T_7330_hpp;
  wire  T_7330_spp;
  wire  T_7330_mpie;
  wire  T_7330_hpie;
  wire  T_7330_spie;
  wire  T_7330_upie;
  wire  T_7330_mie;
  wire  T_7330_hie;
  wire  T_7330_sie;
  wire  T_7330_uie;
  wire [66:0] T_7356;
  wire  T_7357;
  wire  T_7358;
  wire  T_7359;
  wire  T_7360;
  wire  T_7361;
  wire  T_7362;
  wire  T_7363;
  wire  T_7364;
  wire  T_7365;
  wire [1:0] T_7366;
  wire [1:0] T_7367;
  wire [1:0] T_7368;
  wire [1:0] T_7369;
  wire  T_7370;
  wire  T_7371;
  wire  T_7372;
  wire [3:0] T_7373;
  wire [4:0] T_7374;
  wire [1:0] T_7375;
  wire  T_7376;
  wire [30:0] T_7377;
  wire  T_7378;
  wire [1:0] T_7379;
  wire  T_7380;
  wire  T_7382;
  wire [1:0] T_7386;
  wire  GEN_493;
  wire  GEN_494;
  wire [1:0] GEN_495;
  wire  GEN_496;
  wire [1:0] GEN_497;
  wire  T_7415_rocc;
  wire  T_7415_meip;
  wire  T_7415_heip;
  wire  T_7415_seip;
  wire  T_7415_ueip;
  wire  T_7415_mtip;
  wire  T_7415_htip;
  wire  T_7415_stip;
  wire  T_7415_utip;
  wire  T_7415_msip;
  wire  T_7415_hsip;
  wire  T_7415_ssip;
  wire  T_7415_usip;
  wire  GEN_511;
  wire [63:0] T_7443;
  wire [63:0] T_7444;
  wire [63:0] T_7445;
  wire [63:0] GEN_512;
  wire [63:0] GEN_513;
  wire [19:0] T_7446;
  wire [37:0] GEN_514;
  wire [63:0] GEN_515;
  wire [63:0] GEN_516;
  wire [63:0] GEN_517;
  wire [39:0] GEN_518;
  wire [63:0] GEN_937;
  wire [63:0] T_7456;
  wire [63:0] GEN_519;
  wire [63:0] T_7457;
  wire [63:0] GEN_520;
  wire [63:0] T_7459;
  wire [63:0] GEN_521;
  wire [63:0] GEN_522;
  wire [3:0] GEN_17_control_ttype;
  wire  GEN_17_control_dmode;
  wire [5:0] GEN_17_control_maskmax;
  wire [39:0] GEN_17_control_reserved;
  wire  GEN_17_control_action;
  wire  GEN_17_control_chain;
  wire [1:0] GEN_17_control_zero;
  wire [1:0] GEN_17_control_tmatch;
  wire  GEN_17_control_m;
  wire  GEN_17_control_h;
  wire  GEN_17_control_s;
  wire  GEN_17_control_u;
  wire  GEN_17_control_x;
  wire  GEN_17_control_w;
  wire  GEN_17_control_r;
  wire [38:0] GEN_17_address;
  wire  T_7480;
  wire  T_7481;
  wire [3:0] T_7514_ttype;
  wire  T_7514_dmode;
  wire [5:0] T_7514_maskmax;
  wire [39:0] T_7514_reserved;
  wire  T_7514_action;
  wire  T_7514_chain;
  wire [1:0] T_7514_zero;
  wire [1:0] T_7514_tmatch;
  wire  T_7514_m;
  wire  T_7514_h;
  wire  T_7514_s;
  wire  T_7514_u;
  wire  T_7514_x;
  wire  T_7514_w;
  wire  T_7514_r;
  wire [1:0] T_7537;
  wire [1:0] T_7538;
  wire [39:0] T_7541;
  wire [5:0] T_7542;
  wire  T_7543;
  wire [3:0] T_7544;
  wire  T_7545;
  wire [3:0] GEN_18;
  wire  GEN_19;
  wire  GEN_542;
  wire [5:0] GEN_20;
  wire [39:0] GEN_21;
  wire  GEN_22;
  wire  GEN_548;
  wire  GEN_23;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_554;
  wire  GEN_26;
  wire  GEN_556;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_560;
  wire  GEN_29;
  wire  GEN_562;
  wire  GEN_30;
  wire  GEN_564;
  wire  GEN_31;
  wire  GEN_566;
  wire  GEN_32;
  wire  GEN_568;
  wire  GEN_33;
  wire  GEN_570;
  wire  T_7546;
  wire  GEN_34;
  wire  GEN_572;
  wire  GEN_593;
  wire  GEN_602;
  wire [1:0] GEN_611;
  wire  GEN_614;
  wire  GEN_620;
  wire  GEN_623;
  wire  GEN_626;
  wire  GEN_629;
  wire  GEN_632;
  wire [38:0] GEN_35;
  wire [38:0] GEN_636;
  wire [38:0] GEN_639;
  wire  GEN_660;
  wire  GEN_669;
  wire [1:0] GEN_678;
  wire  GEN_681;
  wire  GEN_687;
  wire  GEN_690;
  wire  GEN_693;
  wire  GEN_696;
  wire  GEN_699;
  wire [38:0] GEN_704;
  wire  GEN_731;
  wire  GEN_732;
  wire  GEN_733;
  wire [1:0] GEN_734;
  wire  GEN_735;
  wire  GEN_736;
  wire [1:0] GEN_737;
  wire  GEN_738;
  wire  GEN_739;
  wire [4:0] GEN_740;
  wire [1:0] GEN_741;
  wire  GEN_755;
  wire  GEN_756;
  wire [63:0] GEN_757;
  wire [63:0] GEN_758;
  wire [63:0] GEN_759;
  wire [63:0] GEN_760;
  wire [63:0] GEN_761;
  wire [39:0] GEN_762;
  wire [63:0] GEN_763;
  wire [57:0] GEN_764;
  wire [63:0] GEN_765;
  wire [57:0] GEN_766;
  wire [63:0] GEN_767;
  wire [63:0] GEN_768;
  wire  GEN_786;
  wire  GEN_787;
  wire  GEN_788;
  wire  GEN_789;
  wire  GEN_790;
  wire [1:0] GEN_791;
  wire [63:0] GEN_792;
  wire [63:0] GEN_793;
  wire [63:0] GEN_832;
  wire [37:0] GEN_833;
  wire [63:0] GEN_834;
  wire [63:0] GEN_835;
  wire [63:0] GEN_836;
  wire [39:0] GEN_837;
  wire [63:0] GEN_838;
  wire [63:0] GEN_839;
  wire [63:0] GEN_840;
  wire [63:0] GEN_841;
  wire  GEN_878;
  wire  GEN_887;
  wire [1:0] GEN_896;
  wire  GEN_899;
  wire  GEN_905;
  wire  GEN_908;
  wire  GEN_911;
  wire  GEN_914;
  wire  GEN_917;
  wire [38:0] GEN_922;
  wire  GEN_924;
  wire  GEN_925;
  wire  GEN_926;
  wire  GEN_927;
  wire  GEN_928;
  wire [3:0] T_7607_control_ttype;
  wire  T_7607_control_dmode;
  wire [5:0] T_7607_control_maskmax;
  wire [39:0] T_7607_control_reserved;
  wire  T_7607_control_action;
  wire  T_7607_control_chain;
  wire [1:0] T_7607_control_zero;
  wire [1:0] T_7607_control_tmatch;
  wire  T_7607_control_m;
  wire  T_7607_control_h;
  wire  T_7607_control_s;
  wire  T_7607_control_u;
  wire  T_7607_control_x;
  wire  T_7607_control_w;
  wire  T_7607_control_r;
  wire [38:0] T_7607_address;
  wire [102:0] T_7626;
  wire [38:0] T_7627;
  wire  T_7628;
  wire  T_7629;
  wire  T_7630;
  wire  T_7631;
  wire  T_7632;
  wire  T_7633;
  wire  T_7634;
  wire [1:0] T_7635;
  wire [1:0] T_7636;
  wire  T_7637;
  wire  T_7638;
  wire [39:0] T_7639;
  wire [5:0] T_7640;
  wire  T_7641;
  wire [3:0] T_7642;
  wire  GEN_3;
  reg [31:0] GEN_239;
  wire [6:0] GEN_58;
  reg [31:0] GEN_240;
  wire [4:0] GEN_59;
  reg [31:0] GEN_241;
  wire [4:0] GEN_60;
  reg [31:0] GEN_242;
  wire  GEN_61;
  reg [31:0] GEN_243;
  wire  GEN_62;
  reg [31:0] GEN_244;
  wire  GEN_63;
  reg [31:0] GEN_245;
  wire [4:0] GEN_64;
  reg [31:0] GEN_246;
  wire [6:0] GEN_65;
  reg [31:0] GEN_247;
  wire [63:0] GEN_66;
  reg [63:0] GEN_248;
  wire [63:0] GEN_67;
  reg [63:0] GEN_249;
  wire  GEN_68;
  reg [31:0] GEN_250;
  wire [1:0] GEN_69;
  reg [31:0] GEN_251;
  wire  GEN_70;
  reg [31:0] GEN_252;
  wire [30:0] GEN_71;
  reg [31:0] GEN_253;
  wire  GEN_72;
  reg [31:0] GEN_254;
  wire [1:0] GEN_73;
  reg [31:0] GEN_255;
  wire [4:0] GEN_74;
  reg [31:0] GEN_256;
  wire [3:0] GEN_75;
  reg [31:0] GEN_257;
  wire  GEN_76;
  reg [31:0] GEN_258;
  wire  GEN_77;
  reg [31:0] GEN_259;
  wire  GEN_78;
  reg [31:0] GEN_260;
  wire [1:0] GEN_79;
  reg [31:0] GEN_261;
  wire [1:0] GEN_80;
  reg [31:0] GEN_262;
  wire [1:0] GEN_81;
  reg [31:0] GEN_263;
  wire [1:0] GEN_82;
  reg [31:0] GEN_264;
  wire  GEN_83;
  reg [31:0] GEN_265;
  wire  GEN_84;
  reg [31:0] GEN_266;
  wire  GEN_85;
  reg [31:0] GEN_267;
  wire  GEN_86;
  reg [31:0] GEN_268;
  wire  GEN_87;
  reg [31:0] GEN_269;
  wire  GEN_88;
  reg [31:0] GEN_270;
  wire  GEN_89;
  reg [31:0] GEN_271;
  wire  GEN_90;
  reg [31:0] GEN_272;
  wire  GEN_91;
  reg [31:0] GEN_273;
  wire  GEN_92;
  reg [31:0] GEN_274;
  wire  GEN_93;
  reg [31:0] GEN_275;
  wire  GEN_94;
  reg [31:0] GEN_276;
  wire  GEN_95;
  reg [31:0] GEN_277;
  wire [39:0] GEN_96;
  reg [63:0] GEN_278;
  wire [6:0] GEN_97;
  reg [31:0] GEN_279;
  wire [4:0] GEN_98;
  reg [31:0] GEN_280;
  wire [2:0] GEN_99;
  reg [31:0] GEN_281;
  wire [63:0] GEN_100;
  reg [63:0] GEN_282;
  wire  GEN_101;
  reg [31:0] GEN_283;
  wire  GEN_102;
  reg [31:0] GEN_284;
  wire [63:0] GEN_103;
  reg [63:0] GEN_285;
  wire [63:0] GEN_104;
  reg [63:0] GEN_286;
  wire  GEN_105;
  reg [31:0] GEN_287;
  wire  GEN_106;
  reg [31:0] GEN_288;
  wire  GEN_107;
  reg [31:0] GEN_289;
  wire  GEN_108;
  reg [31:0] GEN_290;
  wire  GEN_109;
  reg [31:0] GEN_291;
  wire  GEN_110;
  reg [31:0] GEN_292;
  wire  GEN_111;
  reg [31:0] GEN_293;
  wire  GEN_112;
  reg [31:0] GEN_294;
  wire [2:0] GEN_113;
  reg [31:0] GEN_295;
  wire [1:0] GEN_114;
  reg [31:0] GEN_296;
  wire [2:0] GEN_115;
  reg [31:0] GEN_297;
  wire  GEN_116;
  reg [31:0] GEN_298;
  wire [3:0] GEN_117;
  reg [31:0] GEN_299;
  wire [63:0] GEN_118;
  reg [63:0] GEN_300;
  wire  GEN_119;
  reg [31:0] GEN_301;
  wire  GEN_120;
  reg [31:0] GEN_302;
  wire [64:0] GEN_121;
  reg [95:0] GEN_303;
  wire [4:0] GEN_122;
  reg [31:0] GEN_304;
  wire  GEN_123;
  reg [31:0] GEN_305;
  assign io_rw_rdata = T_7022;
  assign io_csr_stall = reg_wfi;
  assign io_csr_xcpt = T_6493;
  assign io_eret = insn_ret;
  assign io_singleStep = T_6553;
  assign io_status_debug = reg_debug;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = T_6560;
  assign io_status_zero3 = reg_mstatus_zero3;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_vm = reg_mstatus_vm;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_pum = reg_mstatus_pum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr_asid = reg_sptbr_asid;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = T_6550;
  assign io_fatc = insn_sfence_vm;
  assign io_time = T_5589;
  assign io_fcsr_rm = reg_frm;
  assign io_rocc_cmd_valid = GEN_3;
  assign io_rocc_cmd_bits_inst_funct = GEN_58;
  assign io_rocc_cmd_bits_inst_rs2 = GEN_59;
  assign io_rocc_cmd_bits_inst_rs1 = GEN_60;
  assign io_rocc_cmd_bits_inst_xd = GEN_61;
  assign io_rocc_cmd_bits_inst_xs1 = GEN_62;
  assign io_rocc_cmd_bits_inst_xs2 = GEN_63;
  assign io_rocc_cmd_bits_inst_rd = GEN_64;
  assign io_rocc_cmd_bits_inst_opcode = GEN_65;
  assign io_rocc_cmd_bits_rs1 = GEN_66;
  assign io_rocc_cmd_bits_rs2 = GEN_67;
  assign io_rocc_cmd_bits_status_debug = GEN_68;
  assign io_rocc_cmd_bits_status_prv = GEN_69;
  assign io_rocc_cmd_bits_status_sd = GEN_70;
  assign io_rocc_cmd_bits_status_zero3 = GEN_71;
  assign io_rocc_cmd_bits_status_sd_rv32 = GEN_72;
  assign io_rocc_cmd_bits_status_zero2 = GEN_73;
  assign io_rocc_cmd_bits_status_vm = GEN_74;
  assign io_rocc_cmd_bits_status_zero1 = GEN_75;
  assign io_rocc_cmd_bits_status_mxr = GEN_76;
  assign io_rocc_cmd_bits_status_pum = GEN_77;
  assign io_rocc_cmd_bits_status_mprv = GEN_78;
  assign io_rocc_cmd_bits_status_xs = GEN_79;
  assign io_rocc_cmd_bits_status_fs = GEN_80;
  assign io_rocc_cmd_bits_status_mpp = GEN_81;
  assign io_rocc_cmd_bits_status_hpp = GEN_82;
  assign io_rocc_cmd_bits_status_spp = GEN_83;
  assign io_rocc_cmd_bits_status_mpie = GEN_84;
  assign io_rocc_cmd_bits_status_hpie = GEN_85;
  assign io_rocc_cmd_bits_status_spie = GEN_86;
  assign io_rocc_cmd_bits_status_upie = GEN_87;
  assign io_rocc_cmd_bits_status_mie = GEN_88;
  assign io_rocc_cmd_bits_status_hie = GEN_89;
  assign io_rocc_cmd_bits_status_sie = GEN_90;
  assign io_rocc_cmd_bits_status_uie = GEN_91;
  assign io_rocc_resp_ready = GEN_92;
  assign io_rocc_mem_req_ready = GEN_93;
  assign io_rocc_mem_s2_nack = GEN_94;
  assign io_rocc_mem_resp_valid = GEN_95;
  assign io_rocc_mem_resp_bits_addr = GEN_96;
  assign io_rocc_mem_resp_bits_tag = GEN_97;
  assign io_rocc_mem_resp_bits_cmd = GEN_98;
  assign io_rocc_mem_resp_bits_typ = GEN_99;
  assign io_rocc_mem_resp_bits_data = GEN_100;
  assign io_rocc_mem_resp_bits_replay = GEN_101;
  assign io_rocc_mem_resp_bits_has_data = GEN_102;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_103;
  assign io_rocc_mem_resp_bits_store_data = GEN_104;
  assign io_rocc_mem_replay_next = GEN_105;
  assign io_rocc_mem_xcpt_ma_ld = GEN_106;
  assign io_rocc_mem_xcpt_ma_st = GEN_107;
  assign io_rocc_mem_xcpt_pf_ld = GEN_108;
  assign io_rocc_mem_xcpt_pf_st = GEN_109;
  assign io_rocc_mem_ordered = GEN_110;
  assign io_rocc_autl_acquire_ready = GEN_111;
  assign io_rocc_autl_grant_valid = GEN_112;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_113;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_114;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_115;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_116;
  assign io_rocc_autl_grant_bits_g_type = GEN_117;
  assign io_rocc_autl_grant_bits_data = GEN_118;
  assign io_rocc_fpu_req_ready = GEN_119;
  assign io_rocc_fpu_resp_valid = GEN_120;
  assign io_rocc_fpu_resp_bits_data = GEN_121;
  assign io_rocc_fpu_resp_bits_exc = GEN_122;
  assign io_rocc_exception = GEN_123;
  assign io_interrupt = GEN_40;
  assign io_interrupt_cause = GEN_41;
  assign io_bp_0_control_ttype = reg_bp_0_control_ttype;
  assign io_bp_0_control_dmode = reg_bp_0_control_dmode;
  assign io_bp_0_control_maskmax = reg_bp_0_control_maskmax;
  assign io_bp_0_control_reserved = reg_bp_0_control_reserved;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_chain = reg_bp_0_control_chain;
  assign io_bp_0_control_zero = reg_bp_0_control_zero;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_address = reg_bp_0_address;
  assign T_4982_debug = T_5032;
  assign T_4982_prv = T_5031;
  assign T_4982_sd = T_5030;
  assign T_4982_zero3 = T_5029;
  assign T_4982_sd_rv32 = T_5028;
  assign T_4982_zero2 = T_5027;
  assign T_4982_vm = T_5026;
  assign T_4982_zero1 = T_5025;
  assign T_4982_mxr = T_5024;
  assign T_4982_pum = T_5023;
  assign T_4982_mprv = T_5022;
  assign T_4982_xs = T_5021;
  assign T_4982_fs = T_5020;
  assign T_4982_mpp = T_5019;
  assign T_4982_hpp = T_5018;
  assign T_4982_spp = T_5017;
  assign T_4982_mpie = T_5016;
  assign T_4982_hpie = T_5015;
  assign T_4982_spie = T_5014;
  assign T_4982_upie = T_5013;
  assign T_4982_mie = T_5012;
  assign T_4982_hie = T_5011;
  assign T_4982_sie = T_5010;
  assign T_4982_uie = T_5009;
  assign T_5008 = 67'h0;
  assign T_5009 = T_5008[0];
  assign T_5010 = T_5008[1];
  assign T_5011 = T_5008[2];
  assign T_5012 = T_5008[3];
  assign T_5013 = T_5008[4];
  assign T_5014 = T_5008[5];
  assign T_5015 = T_5008[6];
  assign T_5016 = T_5008[7];
  assign T_5017 = T_5008[8];
  assign T_5018 = T_5008[10:9];
  assign T_5019 = T_5008[12:11];
  assign T_5020 = T_5008[14:13];
  assign T_5021 = T_5008[16:15];
  assign T_5022 = T_5008[17];
  assign T_5023 = T_5008[18];
  assign T_5024 = T_5008[19];
  assign T_5025 = T_5008[23:20];
  assign T_5026 = T_5008[28:24];
  assign T_5027 = T_5008[30:29];
  assign T_5028 = T_5008[31];
  assign T_5029 = T_5008[62:32];
  assign T_5030 = T_5008[63];
  assign T_5031 = T_5008[65:64];
  assign T_5032 = T_5008[66];
  assign reset_mstatus_debug = T_4982_debug;
  assign reset_mstatus_prv = 2'h3;
  assign reset_mstatus_sd = T_4982_sd;
  assign reset_mstatus_zero3 = T_4982_zero3;
  assign reset_mstatus_sd_rv32 = T_4982_sd_rv32;
  assign reset_mstatus_zero2 = T_4982_zero2;
  assign reset_mstatus_vm = T_4982_vm;
  assign reset_mstatus_zero1 = T_4982_zero1;
  assign reset_mstatus_mxr = T_4982_mxr;
  assign reset_mstatus_pum = T_4982_pum;
  assign reset_mstatus_mprv = T_4982_mprv;
  assign reset_mstatus_xs = T_4982_xs;
  assign reset_mstatus_fs = T_4982_fs;
  assign reset_mstatus_mpp = 2'h3;
  assign reset_mstatus_hpp = T_4982_hpp;
  assign reset_mstatus_spp = T_4982_spp;
  assign reset_mstatus_mpie = T_4982_mpie;
  assign reset_mstatus_hpie = T_4982_hpie;
  assign reset_mstatus_spie = T_4982_spie;
  assign reset_mstatus_upie = T_4982_upie;
  assign reset_mstatus_mie = T_4982_mie;
  assign reset_mstatus_hie = T_4982_hie;
  assign reset_mstatus_sie = T_4982_sie;
  assign reset_mstatus_uie = T_4982_uie;
  assign new_prv = GEN_370;
  assign T_5084 = new_prv == 2'h2;
  assign T_5086 = T_5084 ? 2'h0 : new_prv;
  assign T_5124_xdebugver = T_5160;
  assign T_5124_ndreset = T_5159;
  assign T_5124_fullreset = T_5158;
  assign T_5124_zero3 = T_5157;
  assign T_5124_ebreakm = T_5156;
  assign T_5124_ebreakh = T_5155;
  assign T_5124_ebreaks = T_5154;
  assign T_5124_ebreaku = T_5153;
  assign T_5124_zero2 = T_5152;
  assign T_5124_stopcycle = T_5151;
  assign T_5124_stoptime = T_5150;
  assign T_5124_cause = T_5149;
  assign T_5124_debugint = T_5148;
  assign T_5124_zero1 = T_5147;
  assign T_5124_halt = T_5146;
  assign T_5124_step = T_5145;
  assign T_5124_prv = T_5144;
  assign T_5143 = 32'h0;
  assign T_5144 = T_5143[1:0];
  assign T_5145 = T_5143[2];
  assign T_5146 = T_5143[3];
  assign T_5147 = T_5143[4];
  assign T_5148 = T_5143[5];
  assign T_5149 = T_5143[8:6];
  assign T_5150 = T_5143[9];
  assign T_5151 = T_5143[10];
  assign T_5152 = T_5143[11];
  assign T_5153 = T_5143[12];
  assign T_5154 = T_5143[13];
  assign T_5155 = T_5143[14];
  assign T_5156 = T_5143[15];
  assign T_5157 = T_5143[27:16];
  assign T_5158 = T_5143[28];
  assign T_5159 = T_5143[29];
  assign T_5160 = T_5143[31:30];
  assign reset_dcsr_xdebugver = 2'h1;
  assign reset_dcsr_ndreset = T_5124_ndreset;
  assign reset_dcsr_fullreset = T_5124_fullreset;
  assign reset_dcsr_zero3 = T_5124_zero3;
  assign reset_dcsr_ebreakm = T_5124_ebreakm;
  assign reset_dcsr_ebreakh = T_5124_ebreakh;
  assign reset_dcsr_ebreaks = T_5124_ebreaks;
  assign reset_dcsr_ebreaku = T_5124_ebreaku;
  assign reset_dcsr_zero2 = T_5124_zero2;
  assign reset_dcsr_stopcycle = T_5124_stopcycle;
  assign reset_dcsr_stoptime = T_5124_stoptime;
  assign reset_dcsr_cause = T_5124_cause;
  assign reset_dcsr_debugint = T_5124_debugint;
  assign reset_dcsr_zero1 = T_5124_zero1;
  assign reset_dcsr_halt = T_5124_halt;
  assign reset_dcsr_step = T_5124_step;
  assign reset_dcsr_prv = 2'h3;
  assign T_5226_rocc = T_5254;
  assign T_5226_meip = T_5253;
  assign T_5226_heip = T_5252;
  assign T_5226_seip = T_5251;
  assign T_5226_ueip = T_5250;
  assign T_5226_mtip = T_5249;
  assign T_5226_htip = T_5248;
  assign T_5226_stip = T_5247;
  assign T_5226_utip = T_5246;
  assign T_5226_msip = T_5245;
  assign T_5226_hsip = T_5244;
  assign T_5226_ssip = T_5243;
  assign T_5226_usip = T_5242;
  assign T_5241 = 13'h0;
  assign T_5242 = T_5241[0];
  assign T_5243 = T_5241[1];
  assign T_5244 = T_5241[2];
  assign T_5245 = T_5241[3];
  assign T_5246 = T_5241[4];
  assign T_5247 = T_5241[5];
  assign T_5248 = T_5241[6];
  assign T_5249 = T_5241[7];
  assign T_5250 = T_5241[8];
  assign T_5251 = T_5241[9];
  assign T_5252 = T_5241[10];
  assign T_5253 = T_5241[11];
  assign T_5254 = T_5241[12];
  assign T_5255_rocc = 1'h0;
  assign T_5255_meip = 1'h1;
  assign T_5255_heip = T_5226_heip;
  assign T_5255_seip = 1'h1;
  assign T_5255_ueip = T_5226_ueip;
  assign T_5255_mtip = 1'h1;
  assign T_5255_htip = T_5226_htip;
  assign T_5255_stip = 1'h1;
  assign T_5255_utip = T_5226_utip;
  assign T_5255_msip = 1'h1;
  assign T_5255_hsip = T_5226_hsip;
  assign T_5255_ssip = 1'h1;
  assign T_5255_usip = T_5226_usip;
  assign T_5276_rocc = T_5255_rocc;
  assign T_5276_meip = 1'h0;
  assign T_5276_heip = T_5255_heip;
  assign T_5276_seip = T_5255_seip;
  assign T_5276_ueip = T_5255_ueip;
  assign T_5276_mtip = 1'h0;
  assign T_5276_htip = T_5255_htip;
  assign T_5276_stip = T_5255_stip;
  assign T_5276_utip = T_5255_utip;
  assign T_5276_msip = 1'h0;
  assign T_5276_hsip = T_5255_hsip;
  assign T_5276_ssip = T_5255_ssip;
  assign T_5276_usip = T_5255_usip;
  assign T_5293 = {T_5255_hsip,T_5255_ssip};
  assign T_5294 = {T_5293,T_5255_usip};
  assign T_5295 = {T_5255_stip,T_5255_utip};
  assign T_5296 = {T_5295,T_5255_msip};
  assign T_5297 = {T_5296,T_5294};
  assign T_5298 = {T_5255_ueip,T_5255_mtip};
  assign T_5299 = {T_5298,T_5255_htip};
  assign T_5300 = {T_5255_heip,T_5255_seip};
  assign T_5301 = {T_5255_rocc,T_5255_meip};
  assign T_5302 = {T_5301,T_5300};
  assign T_5303 = {T_5302,T_5299};
  assign supported_interrupts = {T_5303,T_5297};
  assign T_5304 = {T_5276_hsip,T_5276_ssip};
  assign T_5305 = {T_5304,T_5276_usip};
  assign T_5306 = {T_5276_stip,T_5276_utip};
  assign T_5307 = {T_5306,T_5276_msip};
  assign T_5308 = {T_5307,T_5305};
  assign T_5309 = {T_5276_ueip,T_5276_mtip};
  assign T_5310 = {T_5309,T_5276_htip};
  assign T_5311 = {T_5276_heip,T_5276_seip};
  assign T_5312 = {T_5276_rocc,T_5276_meip};
  assign T_5313 = {T_5312,T_5311};
  assign T_5314 = {T_5313,T_5310};
  assign delegable_interrupts = {T_5314,T_5308};
  assign exception = io_exception | io_csr_xcpt;
  assign T_5320 = io_retire | exception;
  assign GEN_36 = T_5320 ? 1'h1 : reg_singleStepped;
  assign T_5323 = io_singleStep == 1'h0;
  assign GEN_37 = T_5323 ? 1'h0 : GEN_36;
  assign T_5334 = reg_singleStepped == 1'h0;
  assign T_5336 = io_retire == 1'h0;
  assign T_5337 = T_5334 | T_5336;
  assign T_5338 = T_5337 | reset;
  assign T_5340 = T_5338 == 1'h0;
  assign GEN_0 = {{5'd0}, io_retire};
  assign T_5571 = T_5570 + GEN_0;
  assign T_5574 = T_5571[6];
  assign T_5576 = T_5573 + 58'h1;
  assign T_5577 = T_5576[57:0];
  assign GEN_38 = T_5574 ? T_5577 : T_5573;
  assign T_5578 = {T_5573,T_5570};
  assign T_5582 = T_5581 + 6'h1;
  assign T_5585 = T_5582[6];
  assign T_5587 = T_5584 + 58'h1;
  assign T_5588 = T_5587[57:0];
  assign GEN_39 = T_5585 ? T_5588 : T_5584;
  assign T_5589 = {T_5584,T_5581};
  assign mip_rocc = io_rocc_interrupt;
  assign mip_meip = reg_mip_meip;
  assign mip_heip = reg_mip_heip;
  assign mip_seip = reg_mip_seip;
  assign mip_ueip = reg_mip_ueip;
  assign mip_mtip = reg_mip_mtip;
  assign mip_htip = reg_mip_htip;
  assign mip_stip = reg_mip_stip;
  assign mip_utip = reg_mip_utip;
  assign mip_msip = reg_mip_msip;
  assign mip_hsip = reg_mip_hsip;
  assign mip_ssip = reg_mip_ssip;
  assign mip_usip = reg_mip_usip;
  assign T_5603 = {mip_hsip,mip_ssip};
  assign T_5604 = {T_5603,mip_usip};
  assign T_5605 = {mip_stip,mip_utip};
  assign T_5606 = {T_5605,mip_msip};
  assign T_5607 = {T_5606,T_5604};
  assign T_5608 = {mip_ueip,mip_mtip};
  assign T_5609 = {T_5608,mip_htip};
  assign T_5610 = {mip_heip,mip_seip};
  assign T_5611 = {mip_rocc,mip_meip};
  assign T_5612 = {T_5611,T_5610};
  assign T_5613 = {T_5612,T_5609};
  assign T_5614 = {T_5613,T_5607};
  assign read_mip = T_5614 & supported_interrupts;
  assign GEN_1 = {{51'd0}, read_mip};
  assign pending_interrupts = GEN_1 & reg_mie;
  assign T_5616 = reg_debug == 1'h0;
  assign T_5618 = reg_mstatus_prv < 2'h3;
  assign T_5620 = reg_mstatus_prv == 2'h3;
  assign T_5621 = T_5620 & reg_mstatus_mie;
  assign T_5622 = T_5618 | T_5621;
  assign T_5623 = T_5616 & T_5622;
  assign T_5624 = ~ reg_mideleg;
  assign T_5625 = pending_interrupts & T_5624;
  assign m_interrupts = T_5623 ? T_5625 : 64'h0;
  assign T_5630 = reg_mstatus_prv < 2'h1;
  assign T_5632 = reg_mstatus_prv == 2'h1;
  assign T_5633 = T_5632 & reg_mstatus_sie;
  assign T_5634 = T_5630 | T_5633;
  assign T_5635 = T_5616 & T_5634;
  assign T_5636 = pending_interrupts & reg_mideleg;
  assign s_interrupts = T_5635 ? T_5636 : 64'h0;
  assign all_interrupts = m_interrupts | s_interrupts;
  assign T_5639 = all_interrupts[0];
  assign T_5640 = all_interrupts[1];
  assign T_5641 = all_interrupts[2];
  assign T_5642 = all_interrupts[3];
  assign T_5643 = all_interrupts[4];
  assign T_5644 = all_interrupts[5];
  assign T_5645 = all_interrupts[6];
  assign T_5646 = all_interrupts[7];
  assign T_5647 = all_interrupts[8];
  assign T_5648 = all_interrupts[9];
  assign T_5649 = all_interrupts[10];
  assign T_5650 = all_interrupts[11];
  assign T_5651 = all_interrupts[12];
  assign T_5652 = all_interrupts[13];
  assign T_5653 = all_interrupts[14];
  assign T_5654 = all_interrupts[15];
  assign T_5655 = all_interrupts[16];
  assign T_5656 = all_interrupts[17];
  assign T_5657 = all_interrupts[18];
  assign T_5658 = all_interrupts[19];
  assign T_5659 = all_interrupts[20];
  assign T_5660 = all_interrupts[21];
  assign T_5661 = all_interrupts[22];
  assign T_5662 = all_interrupts[23];
  assign T_5663 = all_interrupts[24];
  assign T_5664 = all_interrupts[25];
  assign T_5665 = all_interrupts[26];
  assign T_5666 = all_interrupts[27];
  assign T_5667 = all_interrupts[28];
  assign T_5668 = all_interrupts[29];
  assign T_5669 = all_interrupts[30];
  assign T_5670 = all_interrupts[31];
  assign T_5671 = all_interrupts[32];
  assign T_5672 = all_interrupts[33];
  assign T_5673 = all_interrupts[34];
  assign T_5674 = all_interrupts[35];
  assign T_5675 = all_interrupts[36];
  assign T_5676 = all_interrupts[37];
  assign T_5677 = all_interrupts[38];
  assign T_5678 = all_interrupts[39];
  assign T_5679 = all_interrupts[40];
  assign T_5680 = all_interrupts[41];
  assign T_5681 = all_interrupts[42];
  assign T_5682 = all_interrupts[43];
  assign T_5683 = all_interrupts[44];
  assign T_5684 = all_interrupts[45];
  assign T_5685 = all_interrupts[46];
  assign T_5686 = all_interrupts[47];
  assign T_5687 = all_interrupts[48];
  assign T_5688 = all_interrupts[49];
  assign T_5689 = all_interrupts[50];
  assign T_5690 = all_interrupts[51];
  assign T_5691 = all_interrupts[52];
  assign T_5692 = all_interrupts[53];
  assign T_5693 = all_interrupts[54];
  assign T_5694 = all_interrupts[55];
  assign T_5695 = all_interrupts[56];
  assign T_5696 = all_interrupts[57];
  assign T_5697 = all_interrupts[58];
  assign T_5698 = all_interrupts[59];
  assign T_5699 = all_interrupts[60];
  assign T_5700 = all_interrupts[61];
  assign T_5701 = all_interrupts[62];
  assign T_5767 = T_5701 ? 6'h3e : 6'h3f;
  assign T_5768 = T_5700 ? 6'h3d : T_5767;
  assign T_5769 = T_5699 ? 6'h3c : T_5768;
  assign T_5770 = T_5698 ? 6'h3b : T_5769;
  assign T_5771 = T_5697 ? 6'h3a : T_5770;
  assign T_5772 = T_5696 ? 6'h39 : T_5771;
  assign T_5773 = T_5695 ? 6'h38 : T_5772;
  assign T_5774 = T_5694 ? 6'h37 : T_5773;
  assign T_5775 = T_5693 ? 6'h36 : T_5774;
  assign T_5776 = T_5692 ? 6'h35 : T_5775;
  assign T_5777 = T_5691 ? 6'h34 : T_5776;
  assign T_5778 = T_5690 ? 6'h33 : T_5777;
  assign T_5779 = T_5689 ? 6'h32 : T_5778;
  assign T_5780 = T_5688 ? 6'h31 : T_5779;
  assign T_5781 = T_5687 ? 6'h30 : T_5780;
  assign T_5782 = T_5686 ? 6'h2f : T_5781;
  assign T_5783 = T_5685 ? 6'h2e : T_5782;
  assign T_5784 = T_5684 ? 6'h2d : T_5783;
  assign T_5785 = T_5683 ? 6'h2c : T_5784;
  assign T_5786 = T_5682 ? 6'h2b : T_5785;
  assign T_5787 = T_5681 ? 6'h2a : T_5786;
  assign T_5788 = T_5680 ? 6'h29 : T_5787;
  assign T_5789 = T_5679 ? 6'h28 : T_5788;
  assign T_5790 = T_5678 ? 6'h27 : T_5789;
  assign T_5791 = T_5677 ? 6'h26 : T_5790;
  assign T_5792 = T_5676 ? 6'h25 : T_5791;
  assign T_5793 = T_5675 ? 6'h24 : T_5792;
  assign T_5794 = T_5674 ? 6'h23 : T_5793;
  assign T_5795 = T_5673 ? 6'h22 : T_5794;
  assign T_5796 = T_5672 ? 6'h21 : T_5795;
  assign T_5797 = T_5671 ? 6'h20 : T_5796;
  assign T_5798 = T_5670 ? 6'h1f : T_5797;
  assign T_5799 = T_5669 ? 6'h1e : T_5798;
  assign T_5800 = T_5668 ? 6'h1d : T_5799;
  assign T_5801 = T_5667 ? 6'h1c : T_5800;
  assign T_5802 = T_5666 ? 6'h1b : T_5801;
  assign T_5803 = T_5665 ? 6'h1a : T_5802;
  assign T_5804 = T_5664 ? 6'h19 : T_5803;
  assign T_5805 = T_5663 ? 6'h18 : T_5804;
  assign T_5806 = T_5662 ? 6'h17 : T_5805;
  assign T_5807 = T_5661 ? 6'h16 : T_5806;
  assign T_5808 = T_5660 ? 6'h15 : T_5807;
  assign T_5809 = T_5659 ? 6'h14 : T_5808;
  assign T_5810 = T_5658 ? 6'h13 : T_5809;
  assign T_5811 = T_5657 ? 6'h12 : T_5810;
  assign T_5812 = T_5656 ? 6'h11 : T_5811;
  assign T_5813 = T_5655 ? 6'h10 : T_5812;
  assign T_5814 = T_5654 ? 6'hf : T_5813;
  assign T_5815 = T_5653 ? 6'he : T_5814;
  assign T_5816 = T_5652 ? 6'hd : T_5815;
  assign T_5817 = T_5651 ? 6'hc : T_5816;
  assign T_5818 = T_5650 ? 6'hb : T_5817;
  assign T_5819 = T_5649 ? 6'ha : T_5818;
  assign T_5820 = T_5648 ? 6'h9 : T_5819;
  assign T_5821 = T_5647 ? 6'h8 : T_5820;
  assign T_5822 = T_5646 ? 6'h7 : T_5821;
  assign T_5823 = T_5645 ? 6'h6 : T_5822;
  assign T_5824 = T_5644 ? 6'h5 : T_5823;
  assign T_5825 = T_5643 ? 6'h4 : T_5824;
  assign T_5826 = T_5642 ? 6'h3 : T_5825;
  assign T_5827 = T_5641 ? 6'h2 : T_5826;
  assign T_5828 = T_5640 ? 6'h1 : T_5827;
  assign T_5829 = T_5639 ? 6'h0 : T_5828;
  assign GEN_2 = {{58'd0}, T_5829};
  assign T_5830 = 64'h8000000000000000 + GEN_2;
  assign interruptCause = T_5830[63:0];
  assign T_5832 = all_interrupts != 64'h0;
  assign T_5835 = T_5832 & T_5323;
  assign T_5836 = T_5835 | reg_singleStepped;
  assign T_5841 = reg_dcsr_debugint & T_5616;
  assign GEN_40 = T_5841 ? 1'h1 : T_5836;
  assign GEN_41 = T_5841 ? 64'h800000000000000d : interruptCause;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T_5844 = io_rw_cmd != 3'h0;
  assign T_5846 = system_insn == 1'h0;
  assign cpu_ren = T_5844 & T_5846;
  assign T_5847 = io_rw_cmd != 3'h5;
  assign cpu_wen = cpu_ren & T_5847;
  assign T_5848 = {io_status_hie,io_status_sie};
  assign T_5849 = {T_5848,io_status_uie};
  assign T_5850 = {io_status_spie,io_status_upie};
  assign T_5851 = {T_5850,io_status_mie};
  assign T_5852 = {T_5851,T_5849};
  assign T_5853 = {io_status_spp,io_status_mpie};
  assign T_5854 = {T_5853,io_status_hpie};
  assign T_5855 = {io_status_fs,io_status_mpp};
  assign T_5856 = {T_5855,io_status_hpp};
  assign T_5857 = {T_5856,T_5854};
  assign T_5858 = {T_5857,T_5852};
  assign T_5859 = {io_status_pum,io_status_mprv};
  assign T_5860 = {T_5859,io_status_xs};
  assign T_5861 = {io_status_vm,io_status_zero1};
  assign T_5862 = {T_5861,io_status_mxr};
  assign T_5863 = {T_5862,T_5860};
  assign T_5864 = {io_status_zero3,io_status_sd_rv32};
  assign T_5865 = {T_5864,io_status_zero2};
  assign T_5866 = {io_status_debug,io_status_prv};
  assign T_5867 = {T_5866,io_status_sd};
  assign T_5868 = {T_5867,T_5865};
  assign T_5869 = {T_5868,T_5863};
  assign T_5870 = {T_5869,T_5858};
  assign read_mstatus = T_5870[63:0];
  assign GEN_0_control_ttype = GEN_42;
  assign GEN_0_control_dmode = GEN_43;
  assign GEN_0_control_maskmax = GEN_44;
  assign GEN_0_control_reserved = GEN_45;
  assign GEN_0_control_action = GEN_46;
  assign GEN_0_control_chain = GEN_47;
  assign GEN_0_control_zero = GEN_48;
  assign GEN_0_control_tmatch = GEN_49;
  assign GEN_0_control_m = GEN_50;
  assign GEN_0_control_h = GEN_51;
  assign GEN_0_control_s = GEN_52;
  assign GEN_0_control_u = GEN_53;
  assign GEN_0_control_x = GEN_54;
  assign GEN_0_control_w = GEN_55;
  assign GEN_0_control_r = GEN_56;
  assign GEN_0_address = GEN_57;
  assign GEN_42 = reg_tselect ? reg_bp_1_control_ttype : reg_bp_0_control_ttype;
  assign GEN_43 = reg_tselect ? reg_bp_1_control_dmode : reg_bp_0_control_dmode;
  assign GEN_44 = reg_tselect ? reg_bp_1_control_maskmax : reg_bp_0_control_maskmax;
  assign GEN_45 = reg_tselect ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign GEN_46 = reg_tselect ? reg_bp_1_control_action : reg_bp_0_control_action;
  assign GEN_47 = reg_tselect ? reg_bp_1_control_chain : reg_bp_0_control_chain;
  assign GEN_48 = reg_tselect ? reg_bp_1_control_zero : reg_bp_0_control_zero;
  assign GEN_49 = reg_tselect ? reg_bp_1_control_tmatch : reg_bp_0_control_tmatch;
  assign GEN_50 = reg_tselect ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign GEN_51 = reg_tselect ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign GEN_52 = reg_tselect ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign GEN_53 = reg_tselect ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign GEN_54 = reg_tselect ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign GEN_55 = reg_tselect ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign GEN_56 = reg_tselect ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign GEN_57 = reg_tselect ? reg_bp_1_address : reg_bp_0_address;
  assign GEN_1_control_ttype = GEN_42;
  assign GEN_1_control_dmode = GEN_43;
  assign GEN_1_control_maskmax = GEN_44;
  assign GEN_1_control_reserved = GEN_45;
  assign GEN_1_control_action = GEN_46;
  assign GEN_1_control_chain = GEN_47;
  assign GEN_1_control_zero = GEN_48;
  assign GEN_1_control_tmatch = GEN_49;
  assign GEN_1_control_m = GEN_50;
  assign GEN_1_control_h = GEN_51;
  assign GEN_1_control_s = GEN_52;
  assign GEN_1_control_u = GEN_53;
  assign GEN_1_control_x = GEN_54;
  assign GEN_1_control_w = GEN_55;
  assign GEN_1_control_r = GEN_56;
  assign GEN_1_address = GEN_57;
  assign T_5888 = {GEN_0_control_x,GEN_1_control_w};
  assign GEN_2_control_ttype = GEN_42;
  assign GEN_2_control_dmode = GEN_43;
  assign GEN_2_control_maskmax = GEN_44;
  assign GEN_2_control_reserved = GEN_45;
  assign GEN_2_control_action = GEN_46;
  assign GEN_2_control_chain = GEN_47;
  assign GEN_2_control_zero = GEN_48;
  assign GEN_2_control_tmatch = GEN_49;
  assign GEN_2_control_m = GEN_50;
  assign GEN_2_control_h = GEN_51;
  assign GEN_2_control_s = GEN_52;
  assign GEN_2_control_u = GEN_53;
  assign GEN_2_control_x = GEN_54;
  assign GEN_2_control_w = GEN_55;
  assign GEN_2_control_r = GEN_56;
  assign GEN_2_address = GEN_57;
  assign T_5889 = {T_5888,GEN_2_control_r};
  assign GEN_3_control_ttype = GEN_42;
  assign GEN_3_control_dmode = GEN_43;
  assign GEN_3_control_maskmax = GEN_44;
  assign GEN_3_control_reserved = GEN_45;
  assign GEN_3_control_action = GEN_46;
  assign GEN_3_control_chain = GEN_47;
  assign GEN_3_control_zero = GEN_48;
  assign GEN_3_control_tmatch = GEN_49;
  assign GEN_3_control_m = GEN_50;
  assign GEN_3_control_h = GEN_51;
  assign GEN_3_control_s = GEN_52;
  assign GEN_3_control_u = GEN_53;
  assign GEN_3_control_x = GEN_54;
  assign GEN_3_control_w = GEN_55;
  assign GEN_3_control_r = GEN_56;
  assign GEN_3_address = GEN_57;
  assign GEN_4_control_ttype = GEN_42;
  assign GEN_4_control_dmode = GEN_43;
  assign GEN_4_control_maskmax = GEN_44;
  assign GEN_4_control_reserved = GEN_45;
  assign GEN_4_control_action = GEN_46;
  assign GEN_4_control_chain = GEN_47;
  assign GEN_4_control_zero = GEN_48;
  assign GEN_4_control_tmatch = GEN_49;
  assign GEN_4_control_m = GEN_50;
  assign GEN_4_control_h = GEN_51;
  assign GEN_4_control_s = GEN_52;
  assign GEN_4_control_u = GEN_53;
  assign GEN_4_control_x = GEN_54;
  assign GEN_4_control_w = GEN_55;
  assign GEN_4_control_r = GEN_56;
  assign GEN_4_address = GEN_57;
  assign T_5890 = {GEN_3_control_s,GEN_4_control_u};
  assign GEN_5_control_ttype = GEN_42;
  assign GEN_5_control_dmode = GEN_43;
  assign GEN_5_control_maskmax = GEN_44;
  assign GEN_5_control_reserved = GEN_45;
  assign GEN_5_control_action = GEN_46;
  assign GEN_5_control_chain = GEN_47;
  assign GEN_5_control_zero = GEN_48;
  assign GEN_5_control_tmatch = GEN_49;
  assign GEN_5_control_m = GEN_50;
  assign GEN_5_control_h = GEN_51;
  assign GEN_5_control_s = GEN_52;
  assign GEN_5_control_u = GEN_53;
  assign GEN_5_control_x = GEN_54;
  assign GEN_5_control_w = GEN_55;
  assign GEN_5_control_r = GEN_56;
  assign GEN_5_address = GEN_57;
  assign GEN_6_control_ttype = GEN_42;
  assign GEN_6_control_dmode = GEN_43;
  assign GEN_6_control_maskmax = GEN_44;
  assign GEN_6_control_reserved = GEN_45;
  assign GEN_6_control_action = GEN_46;
  assign GEN_6_control_chain = GEN_47;
  assign GEN_6_control_zero = GEN_48;
  assign GEN_6_control_tmatch = GEN_49;
  assign GEN_6_control_m = GEN_50;
  assign GEN_6_control_h = GEN_51;
  assign GEN_6_control_s = GEN_52;
  assign GEN_6_control_u = GEN_53;
  assign GEN_6_control_x = GEN_54;
  assign GEN_6_control_w = GEN_55;
  assign GEN_6_control_r = GEN_56;
  assign GEN_6_address = GEN_57;
  assign T_5891 = {GEN_5_control_m,GEN_6_control_h};
  assign T_5892 = {T_5891,T_5890};
  assign T_5893 = {T_5892,T_5889};
  assign GEN_7_control_ttype = GEN_42;
  assign GEN_7_control_dmode = GEN_43;
  assign GEN_7_control_maskmax = GEN_44;
  assign GEN_7_control_reserved = GEN_45;
  assign GEN_7_control_action = GEN_46;
  assign GEN_7_control_chain = GEN_47;
  assign GEN_7_control_zero = GEN_48;
  assign GEN_7_control_tmatch = GEN_49;
  assign GEN_7_control_m = GEN_50;
  assign GEN_7_control_h = GEN_51;
  assign GEN_7_control_s = GEN_52;
  assign GEN_7_control_u = GEN_53;
  assign GEN_7_control_x = GEN_54;
  assign GEN_7_control_w = GEN_55;
  assign GEN_7_control_r = GEN_56;
  assign GEN_7_address = GEN_57;
  assign GEN_8_control_ttype = GEN_42;
  assign GEN_8_control_dmode = GEN_43;
  assign GEN_8_control_maskmax = GEN_44;
  assign GEN_8_control_reserved = GEN_45;
  assign GEN_8_control_action = GEN_46;
  assign GEN_8_control_chain = GEN_47;
  assign GEN_8_control_zero = GEN_48;
  assign GEN_8_control_tmatch = GEN_49;
  assign GEN_8_control_m = GEN_50;
  assign GEN_8_control_h = GEN_51;
  assign GEN_8_control_s = GEN_52;
  assign GEN_8_control_u = GEN_53;
  assign GEN_8_control_x = GEN_54;
  assign GEN_8_control_w = GEN_55;
  assign GEN_8_control_r = GEN_56;
  assign GEN_8_address = GEN_57;
  assign T_5894 = {GEN_7_control_zero,GEN_8_control_tmatch};
  assign GEN_9_control_ttype = GEN_42;
  assign GEN_9_control_dmode = GEN_43;
  assign GEN_9_control_maskmax = GEN_44;
  assign GEN_9_control_reserved = GEN_45;
  assign GEN_9_control_action = GEN_46;
  assign GEN_9_control_chain = GEN_47;
  assign GEN_9_control_zero = GEN_48;
  assign GEN_9_control_tmatch = GEN_49;
  assign GEN_9_control_m = GEN_50;
  assign GEN_9_control_h = GEN_51;
  assign GEN_9_control_s = GEN_52;
  assign GEN_9_control_u = GEN_53;
  assign GEN_9_control_x = GEN_54;
  assign GEN_9_control_w = GEN_55;
  assign GEN_9_control_r = GEN_56;
  assign GEN_9_address = GEN_57;
  assign GEN_10_control_ttype = GEN_42;
  assign GEN_10_control_dmode = GEN_43;
  assign GEN_10_control_maskmax = GEN_44;
  assign GEN_10_control_reserved = GEN_45;
  assign GEN_10_control_action = GEN_46;
  assign GEN_10_control_chain = GEN_47;
  assign GEN_10_control_zero = GEN_48;
  assign GEN_10_control_tmatch = GEN_49;
  assign GEN_10_control_m = GEN_50;
  assign GEN_10_control_h = GEN_51;
  assign GEN_10_control_s = GEN_52;
  assign GEN_10_control_u = GEN_53;
  assign GEN_10_control_x = GEN_54;
  assign GEN_10_control_w = GEN_55;
  assign GEN_10_control_r = GEN_56;
  assign GEN_10_address = GEN_57;
  assign T_5895 = {GEN_9_control_action,GEN_10_control_chain};
  assign T_5896 = {T_5895,T_5894};
  assign GEN_11_control_ttype = GEN_42;
  assign GEN_11_control_dmode = GEN_43;
  assign GEN_11_control_maskmax = GEN_44;
  assign GEN_11_control_reserved = GEN_45;
  assign GEN_11_control_action = GEN_46;
  assign GEN_11_control_chain = GEN_47;
  assign GEN_11_control_zero = GEN_48;
  assign GEN_11_control_tmatch = GEN_49;
  assign GEN_11_control_m = GEN_50;
  assign GEN_11_control_h = GEN_51;
  assign GEN_11_control_s = GEN_52;
  assign GEN_11_control_u = GEN_53;
  assign GEN_11_control_x = GEN_54;
  assign GEN_11_control_w = GEN_55;
  assign GEN_11_control_r = GEN_56;
  assign GEN_11_address = GEN_57;
  assign GEN_12_control_ttype = GEN_42;
  assign GEN_12_control_dmode = GEN_43;
  assign GEN_12_control_maskmax = GEN_44;
  assign GEN_12_control_reserved = GEN_45;
  assign GEN_12_control_action = GEN_46;
  assign GEN_12_control_chain = GEN_47;
  assign GEN_12_control_zero = GEN_48;
  assign GEN_12_control_tmatch = GEN_49;
  assign GEN_12_control_m = GEN_50;
  assign GEN_12_control_h = GEN_51;
  assign GEN_12_control_s = GEN_52;
  assign GEN_12_control_u = GEN_53;
  assign GEN_12_control_x = GEN_54;
  assign GEN_12_control_w = GEN_55;
  assign GEN_12_control_r = GEN_56;
  assign GEN_12_address = GEN_57;
  assign T_5897 = {GEN_11_control_maskmax,GEN_12_control_reserved};
  assign GEN_13_control_ttype = GEN_42;
  assign GEN_13_control_dmode = GEN_43;
  assign GEN_13_control_maskmax = GEN_44;
  assign GEN_13_control_reserved = GEN_45;
  assign GEN_13_control_action = GEN_46;
  assign GEN_13_control_chain = GEN_47;
  assign GEN_13_control_zero = GEN_48;
  assign GEN_13_control_tmatch = GEN_49;
  assign GEN_13_control_m = GEN_50;
  assign GEN_13_control_h = GEN_51;
  assign GEN_13_control_s = GEN_52;
  assign GEN_13_control_u = GEN_53;
  assign GEN_13_control_x = GEN_54;
  assign GEN_13_control_w = GEN_55;
  assign GEN_13_control_r = GEN_56;
  assign GEN_13_address = GEN_57;
  assign GEN_14_control_ttype = GEN_42;
  assign GEN_14_control_dmode = GEN_43;
  assign GEN_14_control_maskmax = GEN_44;
  assign GEN_14_control_reserved = GEN_45;
  assign GEN_14_control_action = GEN_46;
  assign GEN_14_control_chain = GEN_47;
  assign GEN_14_control_zero = GEN_48;
  assign GEN_14_control_tmatch = GEN_49;
  assign GEN_14_control_m = GEN_50;
  assign GEN_14_control_h = GEN_51;
  assign GEN_14_control_s = GEN_52;
  assign GEN_14_control_u = GEN_53;
  assign GEN_14_control_x = GEN_54;
  assign GEN_14_control_w = GEN_55;
  assign GEN_14_control_r = GEN_56;
  assign GEN_14_address = GEN_57;
  assign T_5898 = {GEN_13_control_ttype,GEN_14_control_dmode};
  assign T_5899 = {T_5898,T_5897};
  assign T_5900 = {T_5899,T_5896};
  assign T_5901 = {T_5900,T_5893};
  assign GEN_15_control_ttype = GEN_42;
  assign GEN_15_control_dmode = GEN_43;
  assign GEN_15_control_maskmax = GEN_44;
  assign GEN_15_control_reserved = GEN_45;
  assign GEN_15_control_action = GEN_46;
  assign GEN_15_control_chain = GEN_47;
  assign GEN_15_control_zero = GEN_48;
  assign GEN_15_control_tmatch = GEN_49;
  assign GEN_15_control_m = GEN_50;
  assign GEN_15_control_h = GEN_51;
  assign GEN_15_control_s = GEN_52;
  assign GEN_15_control_u = GEN_53;
  assign GEN_15_control_x = GEN_54;
  assign GEN_15_control_w = GEN_55;
  assign GEN_15_control_r = GEN_56;
  assign GEN_15_address = GEN_57;
  assign T_5919 = GEN_15_address[38];
  assign T_5923 = T_5919 ? 25'h1ffffff : 25'h0;
  assign GEN_16_control_ttype = GEN_42;
  assign GEN_16_control_dmode = GEN_43;
  assign GEN_16_control_maskmax = GEN_44;
  assign GEN_16_control_reserved = GEN_45;
  assign GEN_16_control_action = GEN_46;
  assign GEN_16_control_chain = GEN_47;
  assign GEN_16_control_zero = GEN_48;
  assign GEN_16_control_tmatch = GEN_49;
  assign GEN_16_control_m = GEN_50;
  assign GEN_16_control_h = GEN_51;
  assign GEN_16_control_s = GEN_52;
  assign GEN_16_control_u = GEN_53;
  assign GEN_16_control_x = GEN_54;
  assign GEN_16_control_w = GEN_55;
  assign GEN_16_control_r = GEN_56;
  assign GEN_16_address = GEN_57;
  assign T_5924 = {T_5923,GEN_16_address};
  assign T_5929 = reg_mepc[39];
  assign T_5933 = T_5929 ? 24'hffffff : 24'h0;
  assign T_5934 = {T_5933,reg_mepc};
  assign T_5935 = reg_mbadaddr[39];
  assign T_5939 = T_5935 ? 24'hffffff : 24'h0;
  assign T_5940 = {T_5939,reg_mbadaddr};
  assign T_5941 = {reg_dcsr_step,reg_dcsr_prv};
  assign T_5942 = {reg_dcsr_zero1,reg_dcsr_halt};
  assign T_5943 = {T_5942,T_5941};
  assign T_5944 = {reg_dcsr_cause,reg_dcsr_debugint};
  assign T_5945 = {reg_dcsr_stopcycle,reg_dcsr_stoptime};
  assign T_5946 = {T_5945,T_5944};
  assign T_5947 = {T_5946,T_5943};
  assign T_5948 = {reg_dcsr_ebreaku,reg_dcsr_zero2};
  assign T_5949 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign T_5950 = {T_5949,T_5948};
  assign T_5951 = {reg_dcsr_zero3,reg_dcsr_ebreakm};
  assign T_5952 = {reg_dcsr_xdebugver,reg_dcsr_ndreset};
  assign T_5953 = {T_5952,reg_dcsr_fullreset};
  assign T_5954 = {T_5953,T_5951};
  assign T_5955 = {T_5954,T_5950};
  assign T_5956 = {T_5955,T_5947};
  assign T_5957 = {reg_frm,reg_fflags};
  assign T_5960 = reg_mie & reg_mideleg;
  assign T_5961 = GEN_1 & reg_mideleg;
  assign T_5962_debug = io_status_debug;
  assign T_5962_prv = io_status_prv;
  assign T_5962_sd = io_status_sd;
  assign T_5962_zero3 = io_status_zero3;
  assign T_5962_sd_rv32 = io_status_sd_rv32;
  assign T_5962_zero2 = io_status_zero2;
  assign T_5962_vm = 5'h0;
  assign T_5962_zero1 = io_status_zero1;
  assign T_5962_mxr = io_status_mxr;
  assign T_5962_pum = io_status_pum;
  assign T_5962_mprv = 1'h0;
  assign T_5962_xs = io_status_xs;
  assign T_5962_fs = io_status_fs;
  assign T_5962_mpp = 2'h0;
  assign T_5962_hpp = 2'h0;
  assign T_5962_spp = io_status_spp;
  assign T_5962_mpie = 1'h0;
  assign T_5962_hpie = 1'h0;
  assign T_5962_spie = io_status_spie;
  assign T_5962_upie = io_status_upie;
  assign T_5962_mie = 1'h0;
  assign T_5962_hie = 1'h0;
  assign T_5962_sie = io_status_sie;
  assign T_5962_uie = io_status_uie;
  assign T_5995 = {T_5962_hie,T_5962_sie};
  assign T_5996 = {T_5995,T_5962_uie};
  assign T_5997 = {T_5962_spie,T_5962_upie};
  assign T_5998 = {T_5997,T_5962_mie};
  assign T_5999 = {T_5998,T_5996};
  assign T_6000 = {T_5962_spp,T_5962_mpie};
  assign T_6001 = {T_6000,T_5962_hpie};
  assign T_6002 = {T_5962_fs,T_5962_mpp};
  assign T_6003 = {T_6002,T_5962_hpp};
  assign T_6004 = {T_6003,T_6001};
  assign T_6005 = {T_6004,T_5999};
  assign T_6006 = {T_5962_pum,T_5962_mprv};
  assign T_6007 = {T_6006,T_5962_xs};
  assign T_6008 = {T_5962_vm,T_5962_zero1};
  assign T_6009 = {T_6008,T_5962_mxr};
  assign T_6010 = {T_6009,T_6007};
  assign T_6011 = {T_5962_zero3,T_5962_sd_rv32};
  assign T_6012 = {T_6011,T_5962_zero2};
  assign T_6013 = {T_5962_debug,T_5962_prv};
  assign T_6014 = {T_6013,T_5962_sd};
  assign T_6015 = {T_6014,T_6012};
  assign T_6016 = {T_6015,T_6010};
  assign T_6017 = {T_6016,T_6005};
  assign T_6018 = T_6017[63:0];
  assign T_6019 = reg_sbadaddr[39];
  assign T_6023 = T_6019 ? 24'hffffff : 24'h0;
  assign T_6024 = {T_6023,reg_sbadaddr};
  assign T_6025 = {reg_sptbr_asid,reg_sptbr_ppn};
  assign T_6026 = reg_sepc[39];
  assign T_6030 = T_6026 ? 24'hffffff : 24'h0;
  assign T_6031 = {T_6030,reg_sepc};
  assign T_6032 = reg_stvec[38];
  assign T_6036 = T_6032 ? 25'h1ffffff : 25'h0;
  assign T_6037 = {T_6036,reg_stvec};
  assign T_6039 = io_rw_addr == 12'h7a0;
  assign T_6041 = io_rw_addr == 12'h7a1;
  assign T_6043 = io_rw_addr == 12'h7a2;
  assign T_6045 = io_rw_addr == 12'hf13;
  assign T_6047 = io_rw_addr == 12'hf12;
  assign T_6049 = io_rw_addr == 12'hf11;
  assign T_6051 = io_rw_addr == 12'hb00;
  assign T_6053 = io_rw_addr == 12'hb02;
  assign T_6055 = io_rw_addr == 12'h301;
  assign T_6057 = io_rw_addr == 12'h300;
  assign T_6059 = io_rw_addr == 12'h305;
  assign T_6061 = io_rw_addr == 12'h344;
  assign T_6063 = io_rw_addr == 12'h304;
  assign T_6065 = io_rw_addr == 12'h303;
  assign T_6067 = io_rw_addr == 12'h302;
  assign T_6069 = io_rw_addr == 12'h340;
  assign T_6071 = io_rw_addr == 12'h341;
  assign T_6073 = io_rw_addr == 12'h343;
  assign T_6075 = io_rw_addr == 12'h342;
  assign T_6077 = io_rw_addr == 12'hf14;
  assign T_6079 = io_rw_addr == 12'h7b0;
  assign T_6081 = io_rw_addr == 12'h7b1;
  assign T_6083 = io_rw_addr == 12'h7b2;
  assign T_6085 = io_rw_addr == 12'h1;
  assign T_6087 = io_rw_addr == 12'h2;
  assign T_6089 = io_rw_addr == 12'h3;
  assign T_6091 = io_rw_addr == 12'h323;
  assign T_6093 = io_rw_addr == 12'hb03;
  assign T_6095 = io_rw_addr == 12'hc03;
  assign T_6097 = io_rw_addr == 12'h324;
  assign T_6099 = io_rw_addr == 12'hb04;
  assign T_6101 = io_rw_addr == 12'hc04;
  assign T_6103 = io_rw_addr == 12'h325;
  assign T_6105 = io_rw_addr == 12'hb05;
  assign T_6107 = io_rw_addr == 12'hc05;
  assign T_6109 = io_rw_addr == 12'h326;
  assign T_6111 = io_rw_addr == 12'hb06;
  assign T_6113 = io_rw_addr == 12'hc06;
  assign T_6115 = io_rw_addr == 12'h327;
  assign T_6117 = io_rw_addr == 12'hb07;
  assign T_6119 = io_rw_addr == 12'hc07;
  assign T_6121 = io_rw_addr == 12'h328;
  assign T_6123 = io_rw_addr == 12'hb08;
  assign T_6125 = io_rw_addr == 12'hc08;
  assign T_6127 = io_rw_addr == 12'h329;
  assign T_6129 = io_rw_addr == 12'hb09;
  assign T_6131 = io_rw_addr == 12'hc09;
  assign T_6133 = io_rw_addr == 12'h32a;
  assign T_6135 = io_rw_addr == 12'hb0a;
  assign T_6137 = io_rw_addr == 12'hc0a;
  assign T_6139 = io_rw_addr == 12'h32b;
  assign T_6141 = io_rw_addr == 12'hb0b;
  assign T_6143 = io_rw_addr == 12'hc0b;
  assign T_6145 = io_rw_addr == 12'h32c;
  assign T_6147 = io_rw_addr == 12'hb0c;
  assign T_6149 = io_rw_addr == 12'hc0c;
  assign T_6151 = io_rw_addr == 12'h32d;
  assign T_6153 = io_rw_addr == 12'hb0d;
  assign T_6155 = io_rw_addr == 12'hc0d;
  assign T_6157 = io_rw_addr == 12'h32e;
  assign T_6159 = io_rw_addr == 12'hb0e;
  assign T_6161 = io_rw_addr == 12'hc0e;
  assign T_6163 = io_rw_addr == 12'h32f;
  assign T_6165 = io_rw_addr == 12'hb0f;
  assign T_6167 = io_rw_addr == 12'hc0f;
  assign T_6169 = io_rw_addr == 12'h330;
  assign T_6171 = io_rw_addr == 12'hb10;
  assign T_6173 = io_rw_addr == 12'hc10;
  assign T_6175 = io_rw_addr == 12'h331;
  assign T_6177 = io_rw_addr == 12'hb11;
  assign T_6179 = io_rw_addr == 12'hc11;
  assign T_6181 = io_rw_addr == 12'h332;
  assign T_6183 = io_rw_addr == 12'hb12;
  assign T_6185 = io_rw_addr == 12'hc12;
  assign T_6187 = io_rw_addr == 12'h333;
  assign T_6189 = io_rw_addr == 12'hb13;
  assign T_6191 = io_rw_addr == 12'hc13;
  assign T_6193 = io_rw_addr == 12'h334;
  assign T_6195 = io_rw_addr == 12'hb14;
  assign T_6197 = io_rw_addr == 12'hc14;
  assign T_6199 = io_rw_addr == 12'h335;
  assign T_6201 = io_rw_addr == 12'hb15;
  assign T_6203 = io_rw_addr == 12'hc15;
  assign T_6205 = io_rw_addr == 12'h336;
  assign T_6207 = io_rw_addr == 12'hb16;
  assign T_6209 = io_rw_addr == 12'hc16;
  assign T_6211 = io_rw_addr == 12'h337;
  assign T_6213 = io_rw_addr == 12'hb17;
  assign T_6215 = io_rw_addr == 12'hc17;
  assign T_6217 = io_rw_addr == 12'h338;
  assign T_6219 = io_rw_addr == 12'hb18;
  assign T_6221 = io_rw_addr == 12'hc18;
  assign T_6223 = io_rw_addr == 12'h339;
  assign T_6225 = io_rw_addr == 12'hb19;
  assign T_6227 = io_rw_addr == 12'hc19;
  assign T_6229 = io_rw_addr == 12'h33a;
  assign T_6231 = io_rw_addr == 12'hb1a;
  assign T_6233 = io_rw_addr == 12'hc1a;
  assign T_6235 = io_rw_addr == 12'h33b;
  assign T_6237 = io_rw_addr == 12'hb1b;
  assign T_6239 = io_rw_addr == 12'hc1b;
  assign T_6241 = io_rw_addr == 12'h33c;
  assign T_6243 = io_rw_addr == 12'hb1c;
  assign T_6245 = io_rw_addr == 12'hc1c;
  assign T_6247 = io_rw_addr == 12'h33d;
  assign T_6249 = io_rw_addr == 12'hb1d;
  assign T_6251 = io_rw_addr == 12'hc1d;
  assign T_6253 = io_rw_addr == 12'h33e;
  assign T_6255 = io_rw_addr == 12'hb1e;
  assign T_6257 = io_rw_addr == 12'hc1e;
  assign T_6259 = io_rw_addr == 12'h33f;
  assign T_6261 = io_rw_addr == 12'hb1f;
  assign T_6263 = io_rw_addr == 12'hc1f;
  assign T_6265 = io_rw_addr == 12'h100;
  assign T_6267 = io_rw_addr == 12'h144;
  assign T_6269 = io_rw_addr == 12'h104;
  assign T_6271 = io_rw_addr == 12'h140;
  assign T_6273 = io_rw_addr == 12'h142;
  assign T_6275 = io_rw_addr == 12'h143;
  assign T_6277 = io_rw_addr == 12'h180;
  assign T_6279 = io_rw_addr == 12'h141;
  assign T_6281 = io_rw_addr == 12'h105;
  assign T_6283 = io_rw_addr == 12'h321;
  assign T_6285 = io_rw_addr == 12'h320;
  assign T_6287 = io_rw_addr == 12'hc00;
  assign T_6289 = io_rw_addr == 12'hc02;
  assign T_6290 = T_6039 | T_6041;
  assign T_6291 = T_6290 | T_6043;
  assign T_6292 = T_6291 | T_6045;
  assign T_6293 = T_6292 | T_6047;
  assign T_6294 = T_6293 | T_6049;
  assign T_6295 = T_6294 | T_6051;
  assign T_6296 = T_6295 | T_6053;
  assign T_6297 = T_6296 | T_6055;
  assign T_6298 = T_6297 | T_6057;
  assign T_6299 = T_6298 | T_6059;
  assign T_6300 = T_6299 | T_6061;
  assign T_6301 = T_6300 | T_6063;
  assign T_6302 = T_6301 | T_6065;
  assign T_6303 = T_6302 | T_6067;
  assign T_6304 = T_6303 | T_6069;
  assign T_6305 = T_6304 | T_6071;
  assign T_6306 = T_6305 | T_6073;
  assign T_6307 = T_6306 | T_6075;
  assign T_6308 = T_6307 | T_6077;
  assign T_6309 = T_6308 | T_6079;
  assign T_6310 = T_6309 | T_6081;
  assign T_6311 = T_6310 | T_6083;
  assign T_6312 = T_6311 | T_6085;
  assign T_6313 = T_6312 | T_6087;
  assign T_6314 = T_6313 | T_6089;
  assign T_6315 = T_6314 | T_6091;
  assign T_6316 = T_6315 | T_6093;
  assign T_6317 = T_6316 | T_6095;
  assign T_6318 = T_6317 | T_6097;
  assign T_6319 = T_6318 | T_6099;
  assign T_6320 = T_6319 | T_6101;
  assign T_6321 = T_6320 | T_6103;
  assign T_6322 = T_6321 | T_6105;
  assign T_6323 = T_6322 | T_6107;
  assign T_6324 = T_6323 | T_6109;
  assign T_6325 = T_6324 | T_6111;
  assign T_6326 = T_6325 | T_6113;
  assign T_6327 = T_6326 | T_6115;
  assign T_6328 = T_6327 | T_6117;
  assign T_6329 = T_6328 | T_6119;
  assign T_6330 = T_6329 | T_6121;
  assign T_6331 = T_6330 | T_6123;
  assign T_6332 = T_6331 | T_6125;
  assign T_6333 = T_6332 | T_6127;
  assign T_6334 = T_6333 | T_6129;
  assign T_6335 = T_6334 | T_6131;
  assign T_6336 = T_6335 | T_6133;
  assign T_6337 = T_6336 | T_6135;
  assign T_6338 = T_6337 | T_6137;
  assign T_6339 = T_6338 | T_6139;
  assign T_6340 = T_6339 | T_6141;
  assign T_6341 = T_6340 | T_6143;
  assign T_6342 = T_6341 | T_6145;
  assign T_6343 = T_6342 | T_6147;
  assign T_6344 = T_6343 | T_6149;
  assign T_6345 = T_6344 | T_6151;
  assign T_6346 = T_6345 | T_6153;
  assign T_6347 = T_6346 | T_6155;
  assign T_6348 = T_6347 | T_6157;
  assign T_6349 = T_6348 | T_6159;
  assign T_6350 = T_6349 | T_6161;
  assign T_6351 = T_6350 | T_6163;
  assign T_6352 = T_6351 | T_6165;
  assign T_6353 = T_6352 | T_6167;
  assign T_6354 = T_6353 | T_6169;
  assign T_6355 = T_6354 | T_6171;
  assign T_6356 = T_6355 | T_6173;
  assign T_6357 = T_6356 | T_6175;
  assign T_6358 = T_6357 | T_6177;
  assign T_6359 = T_6358 | T_6179;
  assign T_6360 = T_6359 | T_6181;
  assign T_6361 = T_6360 | T_6183;
  assign T_6362 = T_6361 | T_6185;
  assign T_6363 = T_6362 | T_6187;
  assign T_6364 = T_6363 | T_6189;
  assign T_6365 = T_6364 | T_6191;
  assign T_6366 = T_6365 | T_6193;
  assign T_6367 = T_6366 | T_6195;
  assign T_6368 = T_6367 | T_6197;
  assign T_6369 = T_6368 | T_6199;
  assign T_6370 = T_6369 | T_6201;
  assign T_6371 = T_6370 | T_6203;
  assign T_6372 = T_6371 | T_6205;
  assign T_6373 = T_6372 | T_6207;
  assign T_6374 = T_6373 | T_6209;
  assign T_6375 = T_6374 | T_6211;
  assign T_6376 = T_6375 | T_6213;
  assign T_6377 = T_6376 | T_6215;
  assign T_6378 = T_6377 | T_6217;
  assign T_6379 = T_6378 | T_6219;
  assign T_6380 = T_6379 | T_6221;
  assign T_6381 = T_6380 | T_6223;
  assign T_6382 = T_6381 | T_6225;
  assign T_6383 = T_6382 | T_6227;
  assign T_6384 = T_6383 | T_6229;
  assign T_6385 = T_6384 | T_6231;
  assign T_6386 = T_6385 | T_6233;
  assign T_6387 = T_6386 | T_6235;
  assign T_6388 = T_6387 | T_6237;
  assign T_6389 = T_6388 | T_6239;
  assign T_6390 = T_6389 | T_6241;
  assign T_6391 = T_6390 | T_6243;
  assign T_6392 = T_6391 | T_6245;
  assign T_6393 = T_6392 | T_6247;
  assign T_6394 = T_6393 | T_6249;
  assign T_6395 = T_6394 | T_6251;
  assign T_6396 = T_6395 | T_6253;
  assign T_6397 = T_6396 | T_6255;
  assign T_6398 = T_6397 | T_6257;
  assign T_6399 = T_6398 | T_6259;
  assign T_6400 = T_6399 | T_6261;
  assign T_6401 = T_6400 | T_6263;
  assign T_6402 = T_6401 | T_6265;
  assign T_6403 = T_6402 | T_6267;
  assign T_6404 = T_6403 | T_6269;
  assign T_6405 = T_6404 | T_6271;
  assign T_6406 = T_6405 | T_6273;
  assign T_6407 = T_6406 | T_6275;
  assign T_6408 = T_6407 | T_6277;
  assign T_6409 = T_6408 | T_6279;
  assign T_6410 = T_6409 | T_6281;
  assign T_6411 = T_6410 | T_6283;
  assign T_6412 = T_6411 | T_6285;
  assign T_6413 = T_6412 | T_6287;
  assign addr_valid = T_6413 | T_6289;
  assign T_6414 = T_6085 | T_6087;
  assign fp_csr = T_6414 | T_6089;
  assign T_6416 = io_rw_addr >= 12'hc00;
  assign T_6418 = io_rw_addr < 12'hc20;
  assign hpm_csr = T_6416 & T_6418;
  assign T_6421 = reg_debug | T_5620;
  assign T_6424 = io_rw_addr[4:0];
  assign T_6425 = reg_mscounteren >> T_6424;
  assign T_6426 = T_6425[0];
  assign T_6427 = T_5632 & T_6426;
  assign T_6428 = T_6421 | T_6427;
  assign T_6430 = reg_mstatus_prv == 2'h0;
  assign T_6432 = reg_mucounteren >> T_6424;
  assign T_6433 = T_6432[0];
  assign T_6434 = T_6430 & T_6433;
  assign hpm_en = T_6428 | T_6434;
  assign csr_addr_priv = io_rw_addr[9:8];
  assign T_6437 = io_rw_addr & 12'h90;
  assign T_6439 = T_6437 == 12'h90;
  assign T_6441 = T_6439 == 1'h0;
  assign T_6442 = reg_mstatus_prv >= csr_addr_priv;
  assign T_6443 = T_6441 & T_6442;
  assign priv_sufficient = reg_debug | T_6443;
  assign T_6444 = io_rw_addr[11:10];
  assign T_6445 = ~ T_6444;
  assign read_only = T_6445 == 2'h0;
  assign T_6447 = cpu_wen & priv_sufficient;
  assign T_6449 = read_only == 1'h0;
  assign wen = T_6447 & T_6449;
  assign T_6450 = io_rw_cmd == 3'h2;
  assign T_6451 = io_rw_cmd == 3'h3;
  assign T_6452 = T_6450 | T_6451;
  assign T_6454 = T_6452 ? io_rw_rdata : 64'h0;
  assign T_6455 = io_rw_cmd != 3'h3;
  assign T_6457 = T_6455 ? io_rw_wdata : 64'h0;
  assign T_6458 = T_6454 | T_6457;
  assign T_6461 = T_6451 ? io_rw_wdata : 64'h0;
  assign T_6462 = ~ T_6461;
  assign wdata = T_6458 & T_6462;
  assign do_system_insn = priv_sufficient & system_insn;
  assign T_6464 = io_rw_addr[2:0];
  assign opcode = 8'h1 << T_6464;
  assign T_6465 = opcode[0];
  assign insn_call = do_system_insn & T_6465;
  assign T_6466 = opcode[1];
  assign insn_break = do_system_insn & T_6466;
  assign T_6467 = opcode[2];
  assign insn_ret = do_system_insn & T_6467;
  assign T_6468 = opcode[4];
  assign insn_sfence_vm = do_system_insn & T_6468;
  assign T_6469 = opcode[5];
  assign insn_wfi = do_system_insn & T_6469;
  assign T_6470 = cpu_wen & read_only;
  assign T_6472 = priv_sufficient == 1'h0;
  assign T_6474 = addr_valid == 1'h0;
  assign T_6475 = T_6472 | T_6474;
  assign T_6477 = hpm_en == 1'h0;
  assign T_6478 = hpm_csr & T_6477;
  assign T_6479 = T_6475 | T_6478;
  assign T_6481 = io_status_fs != 2'h0;
  assign T_6483 = T_6481 == 1'h0;
  assign T_6484 = fp_csr & T_6483;
  assign T_6485 = T_6479 | T_6484;
  assign T_6486 = cpu_ren & T_6485;
  assign T_6487 = T_6470 | T_6486;
  assign T_6490 = system_insn & T_6472;
  assign T_6491 = T_6487 | T_6490;
  assign T_6492 = T_6491 | insn_call;
  assign T_6493 = T_6492 | insn_break;
  assign GEN_314 = insn_wfi ? 1'h1 : reg_wfi;
  assign T_6496 = pending_interrupts != 64'h0;
  assign GEN_315 = T_6496 ? 1'h0 : GEN_314;
  assign T_6499 = io_csr_xcpt == 1'h0;
  assign GEN_4 = {{2'd0}, reg_mstatus_prv};
  assign T_6501 = GEN_4 + 4'h8;
  assign T_6502 = T_6501[3:0];
  assign T_6505 = insn_break ? 2'h3 : 2'h2;
  assign T_6506 = insn_call ? T_6502 : {{2'd0}, T_6505};
  assign cause = T_6499 ? io_cause : {{60'd0}, T_6506};
  assign cause_lsbs = cause[5:0];
  assign T_6507 = cause[63];
  assign T_6509 = cause_lsbs == 6'hd;
  assign causeIsDebugInt = T_6507 & T_6509;
  assign T_6512 = T_6507 == 1'h0;
  assign causeIsDebugTrigger = T_6512 & T_6509;
  assign T_6518 = T_6512 & insn_break;
  assign T_6519 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign T_6520 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign T_6521 = {T_6520,T_6519};
  assign T_6522 = T_6521 >> reg_mstatus_prv;
  assign T_6523 = T_6522[0];
  assign causeIsDebugBreak = T_6518 & T_6523;
  assign T_6525 = reg_singleStepped | causeIsDebugInt;
  assign T_6526 = T_6525 | causeIsDebugTrigger;
  assign T_6527 = T_6526 | causeIsDebugBreak;
  assign T_6528 = T_6527 | reg_debug;
  assign T_6534 = reg_mideleg >> cause_lsbs;
  assign T_6535 = T_6534[0];
  assign T_6536 = reg_medeleg >> cause_lsbs;
  assign T_6537 = T_6536[0];
  assign T_6538 = T_6507 ? T_6535 : T_6537;
  assign delegate = T_5618 & T_6538;
  assign debugTVec = reg_debug ? 12'h808 : 12'h800;
  assign T_6542 = {T_6032,reg_stvec};
  assign T_6543 = delegate ? T_6542 : {{8'd0}, reg_mtvec};
  assign tvec = T_6528 ? {{28'd0}, debugTVec} : T_6543;
  assign T_6545 = csr_addr_priv[1];
  assign T_6547 = T_6545 == 1'h0;
  assign T_6549 = T_6547 ? reg_sepc : reg_mepc;
  assign epc = T_6439 ? reg_dpc : T_6549;
  assign T_6550 = exception ? tvec : epc;
  assign T_6553 = reg_dcsr_step & T_5616;
  assign T_6554 = ~ io_status_fs;
  assign T_6556 = T_6554 == 2'h0;
  assign T_6557 = ~ io_status_xs;
  assign T_6559 = T_6557 == 2'h0;
  assign T_6560 = T_6556 | T_6559;
  assign T_6561 = ~ io_pc;
  assign T_6563 = T_6561 | 40'h1;
  assign T_6564 = ~ T_6563;
  assign T_6565 = read_mstatus >> reg_mstatus_prv;
  assign T_6566 = T_6565[0];
  assign T_6574 = cause == 64'h3;
  assign T_6575 = cause == 64'h4;
  assign T_6576 = cause == 64'h6;
  assign T_6577 = cause == 64'h0;
  assign T_6578 = cause == 64'h5;
  assign T_6579 = cause == 64'h7;
  assign T_6580 = cause == 64'h1;
  assign T_6581 = T_6574 | T_6575;
  assign T_6582 = T_6581 | T_6576;
  assign T_6583 = T_6582 | T_6577;
  assign T_6584 = T_6583 | T_6578;
  assign T_6585 = T_6584 | T_6579;
  assign T_6586 = T_6585 | T_6580;
  assign T_6592 = causeIsDebugTrigger ? 2'h2 : 2'h1;
  assign T_6593 = causeIsDebugInt ? 2'h3 : T_6592;
  assign T_6594 = reg_singleStepped ? 3'h4 : {{1'd0}, T_6593};
  assign GEN_316 = T_6528 ? 1'h1 : reg_debug;
  assign GEN_317 = T_6528 ? T_6564 : reg_dpc;
  assign GEN_318 = T_6528 ? T_6594 : reg_dcsr_cause;
  assign GEN_319 = T_6528 ? reg_mstatus_prv : reg_dcsr_prv;
  assign T_6596 = T_6528 == 1'h0;
  assign T_6597 = T_6596 & delegate;
  assign GEN_320 = T_6586 ? io_badaddr : reg_sbadaddr;
  assign GEN_321 = T_6597 ? T_6564 : reg_sepc;
  assign GEN_322 = T_6597 ? cause : reg_scause;
  assign GEN_323 = T_6597 ? GEN_320 : reg_sbadaddr;
  assign GEN_324 = T_6597 ? T_6566 : reg_mstatus_spie;
  assign GEN_325 = T_6597 ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp};
  assign GEN_326 = T_6597 ? 1'h0 : reg_mstatus_sie;
  assign GEN_327 = T_6597 ? 2'h1 : reg_mstatus_prv;
  assign T_6603 = delegate == 1'h0;
  assign T_6604 = T_6596 & T_6603;
  assign GEN_328 = T_6586 ? io_badaddr : reg_mbadaddr;
  assign GEN_329 = T_6604 ? T_6564 : reg_mepc;
  assign GEN_330 = T_6604 ? cause : reg_mcause;
  assign GEN_331 = T_6604 ? GEN_328 : reg_mbadaddr;
  assign GEN_332 = T_6604 ? T_6566 : reg_mstatus_mpie;
  assign GEN_333 = T_6604 ? reg_mstatus_prv : reg_mstatus_mpp;
  assign GEN_334 = T_6604 ? 1'h0 : reg_mstatus_mie;
  assign GEN_335 = T_6604 ? 2'h3 : GEN_327;
  assign GEN_336 = exception ? GEN_316 : reg_debug;
  assign GEN_337 = exception ? GEN_317 : reg_dpc;
  assign GEN_338 = exception ? GEN_318 : reg_dcsr_cause;
  assign GEN_339 = exception ? GEN_319 : reg_dcsr_prv;
  assign GEN_340 = exception ? GEN_321 : reg_sepc;
  assign GEN_341 = exception ? GEN_322 : reg_scause;
  assign GEN_342 = exception ? GEN_323 : reg_sbadaddr;
  assign GEN_343 = exception ? GEN_324 : reg_mstatus_spie;
  assign GEN_344 = exception ? GEN_325 : {{1'd0}, reg_mstatus_spp};
  assign GEN_345 = exception ? GEN_326 : reg_mstatus_sie;
  assign GEN_346 = exception ? GEN_335 : reg_mstatus_prv;
  assign GEN_347 = exception ? GEN_329 : reg_mepc;
  assign GEN_348 = exception ? GEN_330 : reg_mcause;
  assign GEN_349 = exception ? GEN_331 : reg_mbadaddr;
  assign GEN_350 = exception ? GEN_332 : reg_mstatus_mpie;
  assign GEN_351 = exception ? GEN_333 : reg_mstatus_mpp;
  assign GEN_352 = exception ? GEN_334 : reg_mstatus_mie;
  assign GEN_353 = reg_mstatus_spp ? reg_mstatus_spie : GEN_345;
  assign GEN_354 = T_6547 ? GEN_353 : GEN_345;
  assign GEN_355 = T_6547 ? 1'h0 : GEN_343;
  assign GEN_356 = T_6547 ? 2'h0 : GEN_344;
  assign GEN_357 = T_6547 ? {{1'd0}, reg_mstatus_spp} : GEN_346;
  assign T_6616 = T_6547 == 1'h0;
  assign T_6617 = T_6616 & T_6439;
  assign GEN_358 = T_6617 ? reg_dcsr_prv : GEN_357;
  assign GEN_359 = T_6617 ? 1'h0 : GEN_336;
  assign T_6623 = T_6616 & T_6441;
  assign T_6624 = reg_mstatus_mpp[1];
  assign GEN_360 = T_6624 ? reg_mstatus_mpie : GEN_352;
  assign T_6626 = reg_mstatus_mpp[0];
  assign T_6629 = T_6624 == 1'h0;
  assign T_6630 = T_6629 & T_6626;
  assign GEN_361 = T_6630 ? reg_mstatus_mpie : GEN_354;
  assign GEN_362 = T_6623 ? GEN_360 : GEN_352;
  assign GEN_363 = T_6623 ? GEN_361 : GEN_354;
  assign GEN_364 = T_6623 ? 1'h0 : GEN_350;
  assign GEN_365 = T_6623 ? 2'h0 : GEN_351;
  assign GEN_366 = T_6623 ? reg_mstatus_mpp : GEN_358;
  assign GEN_367 = insn_ret ? GEN_363 : GEN_345;
  assign GEN_368 = insn_ret ? GEN_355 : GEN_343;
  assign GEN_369 = insn_ret ? GEN_356 : GEN_344;
  assign GEN_370 = insn_ret ? GEN_366 : GEN_346;
  assign GEN_371 = insn_ret ? GEN_359 : GEN_336;
  assign GEN_372 = insn_ret ? GEN_362 : GEN_352;
  assign GEN_373 = insn_ret ? GEN_364 : GEN_350;
  assign GEN_374 = insn_ret ? GEN_365 : GEN_351;
  assign T_6637 = io_exception + io_csr_xcpt;
  assign GEN_5 = {{1'd0}, insn_ret};
  assign T_6638 = GEN_5 + T_6637;
  assign T_6640 = T_6638 <= 3'h1;
  assign T_6641 = T_6640 | reset;
  assign T_6643 = T_6641 == 1'h0;
  assign T_6645 = T_6039 ? reg_tselect : 1'h0;
  assign T_6647 = T_6041 ? T_5901 : 64'h0;
  assign T_6649 = T_6043 ? T_5924 : 64'h0;
  assign T_6657 = T_6051 ? T_5589 : 64'h0;
  assign T_6659 = T_6053 ? T_5578 : 64'h0;
  assign T_6661 = T_6055 ? 64'h8000000000141129 : 64'h0;
  assign T_6663 = T_6057 ? read_mstatus : 64'h0;
  assign T_6665 = T_6059 ? reg_mtvec : 32'h0;
  assign T_6667 = T_6061 ? read_mip : 13'h0;
  assign T_6669 = T_6063 ? reg_mie : 64'h0;
  assign T_6671 = T_6065 ? reg_mideleg : 64'h0;
  assign T_6673 = T_6067 ? reg_medeleg : 64'h0;
  assign T_6675 = T_6069 ? reg_mscratch : 64'h0;
  assign T_6677 = T_6071 ? T_5934 : 64'h0;
  assign T_6679 = T_6073 ? T_5940 : 64'h0;
  assign T_6681 = T_6075 ? reg_mcause : 64'h0;
  assign T_6683 = T_6077 ? io_prci_id : 1'h0;
  assign T_6685 = T_6079 ? T_5956 : 32'h0;
  assign T_6687 = T_6081 ? reg_dpc : 40'h0;
  assign T_6689 = T_6083 ? reg_dscratch : 64'h0;
  assign T_6691 = T_6085 ? reg_fflags : 5'h0;
  assign T_6693 = T_6087 ? reg_frm : 3'h0;
  assign T_6695 = T_6089 ? T_5957 : 8'h0;
  assign T_6871 = T_6265 ? T_6018 : 64'h0;
  assign T_6873 = T_6267 ? T_5961 : 64'h0;
  assign T_6875 = T_6269 ? T_5960 : 64'h0;
  assign T_6877 = T_6271 ? reg_sscratch : 64'h0;
  assign T_6879 = T_6273 ? reg_scause : 64'h0;
  assign T_6881 = T_6275 ? T_6024 : 64'h0;
  assign T_6883 = T_6277 ? T_6025 : 45'h0;
  assign T_6885 = T_6279 ? T_6031 : 64'h0;
  assign T_6887 = T_6281 ? T_6037 : 64'h0;
  assign T_6889 = T_6283 ? reg_mscounteren : 32'h0;
  assign T_6891 = T_6285 ? reg_mucounteren : 32'h0;
  assign T_6893 = T_6287 ? T_5589 : 64'h0;
  assign T_6895 = T_6289 ? T_5578 : 64'h0;
  assign GEN_6 = {{63'd0}, T_6645};
  assign T_6897 = GEN_6 | T_6647;
  assign T_6898 = T_6897 | T_6649;
  assign T_6902 = T_6898 | T_6657;
  assign T_6903 = T_6902 | T_6659;
  assign T_6904 = T_6903 | T_6661;
  assign T_6905 = T_6904 | T_6663;
  assign GEN_7 = {{32'd0}, T_6665};
  assign T_6906 = T_6905 | GEN_7;
  assign GEN_8 = {{51'd0}, T_6667};
  assign T_6907 = T_6906 | GEN_8;
  assign T_6908 = T_6907 | T_6669;
  assign T_6909 = T_6908 | T_6671;
  assign T_6910 = T_6909 | T_6673;
  assign T_6911 = T_6910 | T_6675;
  assign T_6912 = T_6911 | T_6677;
  assign T_6913 = T_6912 | T_6679;
  assign T_6914 = T_6913 | T_6681;
  assign GEN_9 = {{63'd0}, T_6683};
  assign T_6915 = T_6914 | GEN_9;
  assign GEN_10 = {{32'd0}, T_6685};
  assign T_6916 = T_6915 | GEN_10;
  assign GEN_11 = {{24'd0}, T_6687};
  assign T_6917 = T_6916 | GEN_11;
  assign T_6918 = T_6917 | T_6689;
  assign GEN_12 = {{59'd0}, T_6691};
  assign T_6919 = T_6918 | GEN_12;
  assign GEN_13 = {{61'd0}, T_6693};
  assign T_6920 = T_6919 | GEN_13;
  assign GEN_14 = {{56'd0}, T_6695};
  assign T_6921 = T_6920 | GEN_14;
  assign T_7009 = T_6921 | T_6871;
  assign T_7010 = T_7009 | T_6873;
  assign T_7011 = T_7010 | T_6875;
  assign T_7012 = T_7011 | T_6877;
  assign T_7013 = T_7012 | T_6879;
  assign T_7014 = T_7013 | T_6881;
  assign GEN_15 = {{19'd0}, T_6883};
  assign T_7015 = T_7014 | GEN_15;
  assign T_7016 = T_7015 | T_6885;
  assign T_7017 = T_7016 | T_6887;
  assign GEN_16 = {{32'd0}, T_6889};
  assign T_7018 = T_7017 | GEN_16;
  assign GEN_17 = {{32'd0}, T_6891};
  assign T_7019 = T_7018 | GEN_17;
  assign T_7020 = T_7019 | T_6893;
  assign T_7021 = T_7020 | T_6895;
  assign T_7022 = T_7021;
  assign T_7023 = reg_fflags | io_fcsr_flags_bits;
  assign GEN_375 = io_fcsr_flags_valid ? T_7023 : reg_fflags;
  assign T_7074_debug = T_7124;
  assign T_7074_prv = T_7123;
  assign T_7074_sd = T_7122;
  assign T_7074_zero3 = T_7121;
  assign T_7074_sd_rv32 = T_7120;
  assign T_7074_zero2 = T_7119;
  assign T_7074_vm = T_7118;
  assign T_7074_zero1 = T_7117;
  assign T_7074_mxr = T_7116;
  assign T_7074_pum = T_7115;
  assign T_7074_mprv = T_7114;
  assign T_7074_xs = T_7113;
  assign T_7074_fs = T_7112;
  assign T_7074_mpp = T_7111;
  assign T_7074_hpp = T_7110;
  assign T_7074_spp = T_7109;
  assign T_7074_mpie = T_7108;
  assign T_7074_hpie = T_7107;
  assign T_7074_spie = T_7106;
  assign T_7074_upie = T_7105;
  assign T_7074_mie = T_7104;
  assign T_7074_hie = T_7103;
  assign T_7074_sie = T_7102;
  assign T_7074_uie = T_7101;
  assign T_7100 = {{3'd0}, wdata};
  assign T_7101 = T_7100[0];
  assign T_7102 = T_7100[1];
  assign T_7103 = T_7100[2];
  assign T_7104 = T_7100[3];
  assign T_7105 = T_7100[4];
  assign T_7106 = T_7100[5];
  assign T_7107 = T_7100[6];
  assign T_7108 = T_7100[7];
  assign T_7109 = T_7100[8];
  assign T_7110 = T_7100[10:9];
  assign T_7111 = T_7100[12:11];
  assign T_7112 = T_7100[14:13];
  assign T_7113 = T_7100[16:15];
  assign T_7114 = T_7100[17];
  assign T_7115 = T_7100[18];
  assign T_7116 = T_7100[19];
  assign T_7117 = T_7100[23:20];
  assign T_7118 = T_7100[28:24];
  assign T_7119 = T_7100[30:29];
  assign T_7120 = T_7100[31];
  assign T_7121 = T_7100[62:32];
  assign T_7122 = T_7100[63];
  assign T_7123 = T_7100[65:64];
  assign T_7124 = T_7100[66];
  assign T_7126 = T_7074_vm == 5'h0;
  assign GEN_376 = T_7126 ? 5'h0 : reg_mstatus_vm;
  assign T_7129 = T_7074_vm == 5'h9;
  assign GEN_377 = T_7129 ? 5'h9 : GEN_376;
  assign T_7132 = T_7074_fs != 2'h0;
  assign T_7136 = T_7132 ? 2'h3 : 2'h0;
  assign GEN_403 = T_6057 ? T_7074_mie : GEN_372;
  assign GEN_404 = T_6057 ? T_7074_mpie : GEN_373;
  assign GEN_405 = T_6057 ? T_7074_mprv : reg_mstatus_mprv;
  assign GEN_406 = T_6057 ? T_7074_mpp : GEN_374;
  assign GEN_407 = T_6057 ? T_7074_mxr : reg_mstatus_mxr;
  assign GEN_408 = T_6057 ? T_7074_pum : reg_mstatus_pum;
  assign GEN_409 = T_6057 ? {{1'd0}, T_7074_spp} : GEN_369;
  assign GEN_410 = T_6057 ? T_7074_spie : GEN_368;
  assign GEN_411 = T_6057 ? T_7074_sie : GEN_367;
  assign GEN_412 = T_6057 ? GEN_377 : reg_mstatus_vm;
  assign GEN_413 = T_6057 ? T_7136 : reg_mstatus_fs;
  assign T_7165_rocc = T_7191;
  assign T_7165_meip = T_7190;
  assign T_7165_heip = T_7189;
  assign T_7165_seip = T_7188;
  assign T_7165_ueip = T_7187;
  assign T_7165_mtip = T_7186;
  assign T_7165_htip = T_7185;
  assign T_7165_stip = T_7184;
  assign T_7165_utip = T_7183;
  assign T_7165_msip = T_7182;
  assign T_7165_hsip = T_7181;
  assign T_7165_ssip = T_7180;
  assign T_7165_usip = T_7179;
  assign T_7179 = wdata[0];
  assign T_7180 = wdata[1];
  assign T_7181 = wdata[2];
  assign T_7182 = wdata[3];
  assign T_7183 = wdata[4];
  assign T_7184 = wdata[5];
  assign T_7185 = wdata[6];
  assign T_7186 = wdata[7];
  assign T_7187 = wdata[8];
  assign T_7188 = wdata[9];
  assign T_7189 = wdata[10];
  assign T_7190 = wdata[11];
  assign T_7191 = wdata[12];
  assign GEN_427 = T_6061 ? T_7165_ssip : reg_mip_ssip;
  assign GEN_428 = T_6061 ? T_7165_stip : reg_mip_stip;
  assign GEN_934 = {{51'd0}, supported_interrupts};
  assign T_7192 = wdata & GEN_934;
  assign GEN_429 = T_6063 ? T_7192 : reg_mie;
  assign T_7193 = ~ wdata;
  assign T_7195 = T_7193 | 64'h1;
  assign T_7196 = ~ T_7195;
  assign GEN_430 = T_6071 ? T_7196 : {{24'd0}, GEN_347};
  assign GEN_431 = T_6069 ? wdata : reg_mscratch;
  assign T_7197 = wdata[63:2];
  assign GEN_935 = {{2'd0}, T_7197};
  assign T_7198 = GEN_935 << 2;
  assign GEN_432 = T_6059 ? T_7198 : {{32'd0}, reg_mtvec};
  assign T_7200 = wdata & 64'h800000000000001f;
  assign GEN_433 = T_6075 ? T_7200 : GEN_348;
  assign T_7201 = wdata[39:0];
  assign GEN_434 = T_6073 ? T_7201 : GEN_349;
  assign T_7202 = wdata[63:6];
  assign GEN_435 = T_6051 ? wdata : {{57'd0}, T_5582};
  assign GEN_436 = T_6051 ? T_7202 : GEN_39;
  assign GEN_437 = T_6053 ? wdata : {{57'd0}, T_5571};
  assign GEN_438 = T_6053 ? T_7202 : GEN_38;
  assign GEN_439 = T_6085 ? wdata : {{59'd0}, GEN_375};
  assign GEN_440 = T_6087 ? wdata : {{61'd0}, reg_frm};
  assign T_7204 = wdata[63:5];
  assign GEN_441 = T_6089 ? wdata : GEN_439;
  assign GEN_442 = T_6089 ? {{5'd0}, T_7204} : GEN_440;
  assign T_7241_xdebugver = T_7275;
  assign T_7241_ndreset = T_7274;
  assign T_7241_fullreset = T_7273;
  assign T_7241_zero3 = T_7272;
  assign T_7241_ebreakm = T_7271;
  assign T_7241_ebreakh = T_7270;
  assign T_7241_ebreaks = T_7269;
  assign T_7241_ebreaku = T_7191;
  assign T_7241_zero2 = T_7190;
  assign T_7241_stopcycle = T_7189;
  assign T_7241_stoptime = T_7188;
  assign T_7241_cause = T_7264;
  assign T_7241_debugint = T_7184;
  assign T_7241_zero1 = T_7183;
  assign T_7241_halt = T_7182;
  assign T_7241_step = T_7181;
  assign T_7241_prv = T_7259;
  assign T_7259 = wdata[1:0];
  assign T_7264 = wdata[8:6];
  assign T_7269 = wdata[13];
  assign T_7270 = wdata[14];
  assign T_7271 = wdata[15];
  assign T_7272 = wdata[27:16];
  assign T_7273 = wdata[28];
  assign T_7274 = wdata[29];
  assign T_7275 = wdata[31:30];
  assign GEN_460 = T_6079 ? T_7241_halt : reg_dcsr_halt;
  assign GEN_461 = T_6079 ? T_7241_step : reg_dcsr_step;
  assign GEN_462 = T_6079 ? T_7241_ebreakm : reg_dcsr_ebreakm;
  assign GEN_463 = T_6079 ? T_7241_ebreaks : reg_dcsr_ebreaks;
  assign GEN_464 = T_6079 ? T_7241_ebreaku : reg_dcsr_ebreaku;
  assign GEN_465 = T_6079 ? T_7241_prv : GEN_339;
  assign GEN_466 = T_6081 ? T_7196 : {{24'd0}, GEN_337};
  assign GEN_467 = T_6083 ? wdata : reg_dscratch;
  assign T_7330_debug = T_7380;
  assign T_7330_prv = T_7379;
  assign T_7330_sd = T_7378;
  assign T_7330_zero3 = T_7377;
  assign T_7330_sd_rv32 = T_7376;
  assign T_7330_zero2 = T_7375;
  assign T_7330_vm = T_7374;
  assign T_7330_zero1 = T_7373;
  assign T_7330_mxr = T_7372;
  assign T_7330_pum = T_7371;
  assign T_7330_mprv = T_7370;
  assign T_7330_xs = T_7369;
  assign T_7330_fs = T_7368;
  assign T_7330_mpp = T_7367;
  assign T_7330_hpp = T_7366;
  assign T_7330_spp = T_7365;
  assign T_7330_mpie = T_7364;
  assign T_7330_hpie = T_7363;
  assign T_7330_spie = T_7362;
  assign T_7330_upie = T_7361;
  assign T_7330_mie = T_7360;
  assign T_7330_hie = T_7359;
  assign T_7330_sie = T_7358;
  assign T_7330_uie = T_7357;
  assign T_7356 = {{3'd0}, wdata};
  assign T_7357 = T_7356[0];
  assign T_7358 = T_7356[1];
  assign T_7359 = T_7356[2];
  assign T_7360 = T_7356[3];
  assign T_7361 = T_7356[4];
  assign T_7362 = T_7356[5];
  assign T_7363 = T_7356[6];
  assign T_7364 = T_7356[7];
  assign T_7365 = T_7356[8];
  assign T_7366 = T_7356[10:9];
  assign T_7367 = T_7356[12:11];
  assign T_7368 = T_7356[14:13];
  assign T_7369 = T_7356[16:15];
  assign T_7370 = T_7356[17];
  assign T_7371 = T_7356[18];
  assign T_7372 = T_7356[19];
  assign T_7373 = T_7356[23:20];
  assign T_7374 = T_7356[28:24];
  assign T_7375 = T_7356[30:29];
  assign T_7376 = T_7356[31];
  assign T_7377 = T_7356[62:32];
  assign T_7378 = T_7356[63];
  assign T_7379 = T_7356[65:64];
  assign T_7380 = T_7356[66];
  assign T_7382 = T_7330_fs != 2'h0;
  assign T_7386 = T_7382 ? 2'h3 : 2'h0;
  assign GEN_493 = T_6265 ? T_7330_sie : GEN_411;
  assign GEN_494 = T_6265 ? T_7330_spie : GEN_410;
  assign GEN_495 = T_6265 ? {{1'd0}, T_7330_spp} : GEN_409;
  assign GEN_496 = T_6265 ? T_7330_pum : GEN_408;
  assign GEN_497 = T_6265 ? T_7386 : GEN_413;
  assign T_7415_rocc = T_7191;
  assign T_7415_meip = T_7190;
  assign T_7415_heip = T_7189;
  assign T_7415_seip = T_7188;
  assign T_7415_ueip = T_7187;
  assign T_7415_mtip = T_7186;
  assign T_7415_htip = T_7185;
  assign T_7415_stip = T_7184;
  assign T_7415_utip = T_7183;
  assign T_7415_msip = T_7182;
  assign T_7415_hsip = T_7181;
  assign T_7415_ssip = T_7180;
  assign T_7415_usip = T_7179;
  assign GEN_511 = T_6267 ? T_7415_ssip : GEN_427;
  assign T_7443 = reg_mie & T_5624;
  assign T_7444 = wdata & reg_mideleg;
  assign T_7445 = T_7443 | T_7444;
  assign GEN_512 = T_6269 ? T_7445 : GEN_429;
  assign GEN_513 = T_6271 ? wdata : reg_sscratch;
  assign T_7446 = wdata[19:0];
  assign GEN_514 = T_6277 ? {{18'd0}, T_7446} : reg_sptbr_ppn;
  assign GEN_515 = T_6279 ? T_7196 : {{24'd0}, GEN_340};
  assign GEN_516 = T_6281 ? T_7198 : {{25'd0}, reg_stvec};
  assign GEN_517 = T_6273 ? T_7200 : GEN_341;
  assign GEN_518 = T_6275 ? T_7201 : GEN_342;
  assign GEN_937 = {{51'd0}, delegable_interrupts};
  assign T_7456 = wdata & GEN_937;
  assign GEN_519 = T_6065 ? T_7456 : reg_mideleg;
  assign T_7457 = wdata & 64'h1ab;
  assign GEN_520 = T_6067 ? T_7457 : reg_medeleg;
  assign T_7459 = wdata & 64'h7;
  assign GEN_521 = T_6283 ? T_7459 : {{32'd0}, reg_mscounteren};
  assign GEN_522 = T_6285 ? T_7459 : {{32'd0}, reg_mucounteren};
  assign GEN_17_control_ttype = GEN_42;
  assign GEN_17_control_dmode = GEN_43;
  assign GEN_17_control_maskmax = GEN_44;
  assign GEN_17_control_reserved = GEN_45;
  assign GEN_17_control_action = GEN_46;
  assign GEN_17_control_chain = GEN_47;
  assign GEN_17_control_zero = GEN_48;
  assign GEN_17_control_tmatch = GEN_49;
  assign GEN_17_control_m = GEN_50;
  assign GEN_17_control_h = GEN_51;
  assign GEN_17_control_s = GEN_52;
  assign GEN_17_control_u = GEN_53;
  assign GEN_17_control_x = GEN_54;
  assign GEN_17_control_w = GEN_55;
  assign GEN_17_control_r = GEN_56;
  assign GEN_17_address = GEN_57;
  assign T_7480 = GEN_17_control_dmode == 1'h0;
  assign T_7481 = T_7480 | reg_debug;
  assign T_7514_ttype = T_7544;
  assign T_7514_dmode = T_7543;
  assign T_7514_maskmax = T_7542;
  assign T_7514_reserved = T_7541;
  assign T_7514_action = T_7191;
  assign T_7514_chain = T_7190;
  assign T_7514_zero = T_7538;
  assign T_7514_tmatch = T_7537;
  assign T_7514_m = T_7185;
  assign T_7514_h = T_7184;
  assign T_7514_s = T_7183;
  assign T_7514_u = T_7182;
  assign T_7514_x = T_7181;
  assign T_7514_w = T_7180;
  assign T_7514_r = T_7179;
  assign T_7537 = wdata[8:7];
  assign T_7538 = wdata[10:9];
  assign T_7541 = wdata[52:13];
  assign T_7542 = wdata[58:53];
  assign T_7543 = wdata[59];
  assign T_7544 = wdata[63:60];
  assign T_7545 = T_7514_dmode & reg_debug;
  assign GEN_18 = T_7514_ttype;
  assign GEN_19 = T_7514_dmode;
  assign GEN_542 = 1'h0 == reg_tselect ? GEN_19 : reg_bp_0_control_dmode;
  assign GEN_20 = T_7514_maskmax;
  assign GEN_21 = T_7514_reserved;
  assign GEN_22 = T_7514_action;
  assign GEN_548 = 1'h0 == reg_tselect ? GEN_22 : reg_bp_0_control_action;
  assign GEN_23 = T_7514_chain;
  assign GEN_24 = T_7514_zero;
  assign GEN_25 = T_7514_tmatch;
  assign GEN_554 = 1'h0 == reg_tselect ? GEN_25 : reg_bp_0_control_tmatch;
  assign GEN_26 = T_7514_m;
  assign GEN_556 = 1'h0 == reg_tselect ? GEN_26 : reg_bp_0_control_m;
  assign GEN_27 = T_7514_h;
  assign GEN_28 = T_7514_s;
  assign GEN_560 = 1'h0 == reg_tselect ? GEN_28 : reg_bp_0_control_s;
  assign GEN_29 = T_7514_u;
  assign GEN_562 = 1'h0 == reg_tselect ? GEN_29 : reg_bp_0_control_u;
  assign GEN_30 = T_7514_x;
  assign GEN_564 = 1'h0 == reg_tselect ? GEN_30 : reg_bp_0_control_x;
  assign GEN_31 = T_7514_w;
  assign GEN_566 = 1'h0 == reg_tselect ? GEN_31 : reg_bp_0_control_w;
  assign GEN_32 = T_7514_r;
  assign GEN_568 = 1'h0 == reg_tselect ? GEN_32 : reg_bp_0_control_r;
  assign GEN_33 = T_7545;
  assign GEN_570 = 1'h0 == reg_tselect ? GEN_33 : GEN_542;
  assign T_7546 = T_7545 & T_7514_action;
  assign GEN_34 = T_7546;
  assign GEN_572 = 1'h0 == reg_tselect ? GEN_34 : GEN_548;
  assign GEN_593 = T_6041 ? GEN_570 : reg_bp_0_control_dmode;
  assign GEN_602 = T_6041 ? GEN_572 : reg_bp_0_control_action;
  assign GEN_611 = T_6041 ? GEN_554 : reg_bp_0_control_tmatch;
  assign GEN_614 = T_6041 ? GEN_556 : reg_bp_0_control_m;
  assign GEN_620 = T_6041 ? GEN_560 : reg_bp_0_control_s;
  assign GEN_623 = T_6041 ? GEN_562 : reg_bp_0_control_u;
  assign GEN_626 = T_6041 ? GEN_564 : reg_bp_0_control_x;
  assign GEN_629 = T_6041 ? GEN_566 : reg_bp_0_control_w;
  assign GEN_632 = T_6041 ? GEN_568 : reg_bp_0_control_r;
  assign GEN_35 = wdata[38:0];
  assign GEN_636 = 1'h0 == reg_tselect ? GEN_35 : reg_bp_0_address;
  assign GEN_639 = T_6043 ? GEN_636 : reg_bp_0_address;
  assign GEN_660 = T_7481 ? GEN_593 : reg_bp_0_control_dmode;
  assign GEN_669 = T_7481 ? GEN_602 : reg_bp_0_control_action;
  assign GEN_678 = T_7481 ? GEN_611 : reg_bp_0_control_tmatch;
  assign GEN_681 = T_7481 ? GEN_614 : reg_bp_0_control_m;
  assign GEN_687 = T_7481 ? GEN_620 : reg_bp_0_control_s;
  assign GEN_690 = T_7481 ? GEN_623 : reg_bp_0_control_u;
  assign GEN_693 = T_7481 ? GEN_626 : reg_bp_0_control_x;
  assign GEN_696 = T_7481 ? GEN_629 : reg_bp_0_control_w;
  assign GEN_699 = T_7481 ? GEN_632 : reg_bp_0_control_r;
  assign GEN_704 = T_7481 ? GEN_639 : reg_bp_0_address;
  assign GEN_731 = wen ? GEN_403 : GEN_372;
  assign GEN_732 = wen ? GEN_404 : GEN_373;
  assign GEN_733 = wen ? GEN_405 : reg_mstatus_mprv;
  assign GEN_734 = wen ? GEN_406 : GEN_374;
  assign GEN_735 = wen ? GEN_407 : reg_mstatus_mxr;
  assign GEN_736 = wen ? GEN_496 : reg_mstatus_pum;
  assign GEN_737 = wen ? GEN_495 : GEN_369;
  assign GEN_738 = wen ? GEN_494 : GEN_368;
  assign GEN_739 = wen ? GEN_493 : GEN_367;
  assign GEN_740 = wen ? GEN_412 : reg_mstatus_vm;
  assign GEN_741 = wen ? GEN_497 : reg_mstatus_fs;
  assign GEN_755 = wen ? GEN_511 : reg_mip_ssip;
  assign GEN_756 = wen ? GEN_428 : reg_mip_stip;
  assign GEN_757 = wen ? GEN_512 : reg_mie;
  assign GEN_758 = wen ? GEN_430 : {{24'd0}, GEN_347};
  assign GEN_759 = wen ? GEN_431 : reg_mscratch;
  assign GEN_760 = wen ? GEN_432 : {{32'd0}, reg_mtvec};
  assign GEN_761 = wen ? GEN_433 : GEN_348;
  assign GEN_762 = wen ? GEN_434 : GEN_349;
  assign GEN_763 = wen ? GEN_435 : {{57'd0}, T_5582};
  assign GEN_764 = wen ? GEN_436 : GEN_39;
  assign GEN_765 = wen ? GEN_437 : {{57'd0}, T_5571};
  assign GEN_766 = wen ? GEN_438 : GEN_38;
  assign GEN_767 = wen ? GEN_441 : {{59'd0}, GEN_375};
  assign GEN_768 = wen ? GEN_442 : {{61'd0}, reg_frm};
  assign GEN_786 = wen ? GEN_460 : reg_dcsr_halt;
  assign GEN_787 = wen ? GEN_461 : reg_dcsr_step;
  assign GEN_788 = wen ? GEN_462 : reg_dcsr_ebreakm;
  assign GEN_789 = wen ? GEN_463 : reg_dcsr_ebreaks;
  assign GEN_790 = wen ? GEN_464 : reg_dcsr_ebreaku;
  assign GEN_791 = wen ? GEN_465 : GEN_339;
  assign GEN_792 = wen ? GEN_466 : {{24'd0}, GEN_337};
  assign GEN_793 = wen ? GEN_467 : reg_dscratch;
  assign GEN_832 = wen ? GEN_513 : reg_sscratch;
  assign GEN_833 = wen ? GEN_514 : reg_sptbr_ppn;
  assign GEN_834 = wen ? GEN_515 : {{24'd0}, GEN_340};
  assign GEN_835 = wen ? GEN_516 : {{25'd0}, reg_stvec};
  assign GEN_836 = wen ? GEN_517 : GEN_341;
  assign GEN_837 = wen ? GEN_518 : GEN_342;
  assign GEN_838 = wen ? GEN_519 : reg_mideleg;
  assign GEN_839 = wen ? GEN_520 : reg_medeleg;
  assign GEN_840 = wen ? GEN_521 : {{32'd0}, reg_mscounteren};
  assign GEN_841 = wen ? GEN_522 : {{32'd0}, reg_mucounteren};
  assign GEN_878 = wen ? GEN_660 : reg_bp_0_control_dmode;
  assign GEN_887 = wen ? GEN_669 : reg_bp_0_control_action;
  assign GEN_896 = wen ? GEN_678 : reg_bp_0_control_tmatch;
  assign GEN_899 = wen ? GEN_681 : reg_bp_0_control_m;
  assign GEN_905 = wen ? GEN_687 : reg_bp_0_control_s;
  assign GEN_908 = wen ? GEN_690 : reg_bp_0_control_u;
  assign GEN_911 = wen ? GEN_693 : reg_bp_0_control_x;
  assign GEN_914 = wen ? GEN_696 : reg_bp_0_control_w;
  assign GEN_917 = wen ? GEN_699 : reg_bp_0_control_r;
  assign GEN_922 = wen ? GEN_704 : reg_bp_0_address;
  assign GEN_924 = reset ? 1'h0 : GEN_887;
  assign GEN_925 = reset ? 1'h0 : GEN_878;
  assign GEN_926 = reset ? 1'h0 : GEN_917;
  assign GEN_927 = reset ? 1'h0 : GEN_914;
  assign GEN_928 = reset ? 1'h0 : GEN_911;
  assign T_7607_control_ttype = T_7642;
  assign T_7607_control_dmode = T_7641;
  assign T_7607_control_maskmax = T_7640;
  assign T_7607_control_reserved = T_7639;
  assign T_7607_control_action = T_7638;
  assign T_7607_control_chain = T_7637;
  assign T_7607_control_zero = T_7636;
  assign T_7607_control_tmatch = T_7635;
  assign T_7607_control_m = T_7634;
  assign T_7607_control_h = T_7633;
  assign T_7607_control_s = T_7632;
  assign T_7607_control_u = T_7631;
  assign T_7607_control_x = T_7630;
  assign T_7607_control_w = T_7629;
  assign T_7607_control_r = T_7628;
  assign T_7607_address = T_7627;
  assign T_7626 = 103'h0;
  assign T_7627 = T_7626[38:0];
  assign T_7628 = T_7626[39];
  assign T_7629 = T_7626[40];
  assign T_7630 = T_7626[41];
  assign T_7631 = T_7626[42];
  assign T_7632 = T_7626[43];
  assign T_7633 = T_7626[44];
  assign T_7634 = T_7626[45];
  assign T_7635 = T_7626[47:46];
  assign T_7636 = T_7626[49:48];
  assign T_7637 = T_7626[50];
  assign T_7638 = T_7626[51];
  assign T_7639 = T_7626[91:52];
  assign T_7640 = T_7626[97:92];
  assign T_7641 = T_7626[98];
  assign T_7642 = T_7626[102:99];
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_58 = GEN_240[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_241[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_242[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_243[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_244[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_245[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_64 = GEN_246[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_65 = GEN_247[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_66 = GEN_248[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_67 = GEN_249[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_250[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_69 = GEN_251[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_70 = GEN_252[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_71 = GEN_253[30:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_72 = GEN_254[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_73 = GEN_255[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_74 = GEN_256[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_75 = GEN_257[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_76 = GEN_258[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_77 = GEN_259[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_78 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_79 = GEN_261[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_80 = GEN_262[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_81 = GEN_263[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_82 = GEN_264[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_83 = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_84 = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_85 = GEN_267[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_86 = GEN_268[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_87 = GEN_269[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_88 = GEN_270[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_89 = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_90 = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_91 = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_92 = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_93 = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_94 = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_95 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_96 = GEN_278[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_97 = GEN_279[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_98 = GEN_280[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_99 = GEN_281[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_100 = GEN_282[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_101 = GEN_283[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_102 = GEN_284[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_103 = GEN_285[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_104 = GEN_286[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_105 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_106 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_107 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_108 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_109 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_110 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_111 = GEN_293[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_112 = GEN_294[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_113 = GEN_295[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_114 = GEN_296[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_115 = GEN_297[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_116 = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_117 = GEN_299[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_118 = GEN_300[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_119 = GEN_301[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_120 = GEN_302[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_121 = GEN_303[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_122 = GEN_304[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_123 = GEN_305[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_124 = {1{$random}};
  reg_mstatus_debug = GEN_124[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  reg_mstatus_prv = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {1{$random}};
  reg_mstatus_sd = GEN_126[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {1{$random}};
  reg_mstatus_zero3 = GEN_127[30:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {1{$random}};
  reg_mstatus_sd_rv32 = GEN_128[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {1{$random}};
  reg_mstatus_zero2 = GEN_129[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {1{$random}};
  reg_mstatus_vm = GEN_130[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  reg_mstatus_zero1 = GEN_131[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  reg_mstatus_mxr = GEN_132[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  reg_mstatus_pum = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  reg_mstatus_mprv = GEN_134[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  reg_mstatus_xs = GEN_135[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {1{$random}};
  reg_mstatus_fs = GEN_136[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  reg_mstatus_mpp = GEN_137[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  reg_mstatus_hpp = GEN_138[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  reg_mstatus_spp = GEN_139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  reg_mstatus_mpie = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  reg_mstatus_hpie = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  reg_mstatus_spie = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  reg_mstatus_upie = GEN_143[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  reg_mstatus_mie = GEN_144[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  reg_mstatus_hie = GEN_145[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  reg_mstatus_sie = GEN_146[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  reg_mstatus_uie = GEN_147[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {1{$random}};
  reg_dcsr_xdebugver = GEN_148[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  reg_dcsr_ndreset = GEN_149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  reg_dcsr_fullreset = GEN_150[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  reg_dcsr_zero3 = GEN_151[11:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  reg_dcsr_ebreakm = GEN_152[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  reg_dcsr_ebreakh = GEN_153[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  reg_dcsr_ebreaks = GEN_154[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  reg_dcsr_ebreaku = GEN_155[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  reg_dcsr_zero2 = GEN_156[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  reg_dcsr_stopcycle = GEN_157[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  reg_dcsr_stoptime = GEN_158[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  reg_dcsr_cause = GEN_159[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {1{$random}};
  reg_dcsr_debugint = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  reg_dcsr_zero1 = GEN_161[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {1{$random}};
  reg_dcsr_halt = GEN_162[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {1{$random}};
  reg_dcsr_step = GEN_163[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {1{$random}};
  reg_dcsr_prv = GEN_164[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {1{$random}};
  reg_debug = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_166 = {2{$random}};
  reg_dpc = GEN_166[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_167 = {2{$random}};
  reg_dscratch = GEN_167[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_168 = {1{$random}};
  reg_singleStepped = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_169 = {1{$random}};
  reg_tselect = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_170 = {1{$random}};
  reg_bp_0_control_ttype = GEN_170[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_171 = {1{$random}};
  reg_bp_0_control_dmode = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_172 = {1{$random}};
  reg_bp_0_control_maskmax = GEN_172[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_173 = {2{$random}};
  reg_bp_0_control_reserved = GEN_173[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_174 = {1{$random}};
  reg_bp_0_control_action = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_175 = {1{$random}};
  reg_bp_0_control_chain = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_176 = {1{$random}};
  reg_bp_0_control_zero = GEN_176[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_177 = {1{$random}};
  reg_bp_0_control_tmatch = GEN_177[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_178 = {1{$random}};
  reg_bp_0_control_m = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_179 = {1{$random}};
  reg_bp_0_control_h = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_180 = {1{$random}};
  reg_bp_0_control_s = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_181 = {1{$random}};
  reg_bp_0_control_u = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_182 = {1{$random}};
  reg_bp_0_control_x = GEN_182[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_183 = {1{$random}};
  reg_bp_0_control_w = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_184 = {1{$random}};
  reg_bp_0_control_r = GEN_184[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_185 = {2{$random}};
  reg_bp_0_address = GEN_185[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_186 = {1{$random}};
  reg_bp_1_control_ttype = GEN_186[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_187 = {1{$random}};
  reg_bp_1_control_dmode = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_188 = {1{$random}};
  reg_bp_1_control_maskmax = GEN_188[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_189 = {2{$random}};
  reg_bp_1_control_reserved = GEN_189[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_190 = {1{$random}};
  reg_bp_1_control_action = GEN_190[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_191 = {1{$random}};
  reg_bp_1_control_chain = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_192 = {1{$random}};
  reg_bp_1_control_zero = GEN_192[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_193 = {1{$random}};
  reg_bp_1_control_tmatch = GEN_193[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_194 = {1{$random}};
  reg_bp_1_control_m = GEN_194[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_195 = {1{$random}};
  reg_bp_1_control_h = GEN_195[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_196 = {1{$random}};
  reg_bp_1_control_s = GEN_196[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_197 = {1{$random}};
  reg_bp_1_control_u = GEN_197[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_198 = {1{$random}};
  reg_bp_1_control_x = GEN_198[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_199 = {1{$random}};
  reg_bp_1_control_w = GEN_199[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_200 = {1{$random}};
  reg_bp_1_control_r = GEN_200[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_201 = {2{$random}};
  reg_bp_1_address = GEN_201[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_202 = {2{$random}};
  reg_mie = GEN_202[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_203 = {2{$random}};
  reg_mideleg = GEN_203[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_204 = {2{$random}};
  reg_medeleg = GEN_204[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_205 = {1{$random}};
  reg_mip_rocc = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_206 = {1{$random}};
  reg_mip_meip = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_207 = {1{$random}};
  reg_mip_heip = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_208 = {1{$random}};
  reg_mip_seip = GEN_208[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_209 = {1{$random}};
  reg_mip_ueip = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_210 = {1{$random}};
  reg_mip_mtip = GEN_210[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_211 = {1{$random}};
  reg_mip_htip = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_212 = {1{$random}};
  reg_mip_stip = GEN_212[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_213 = {1{$random}};
  reg_mip_utip = GEN_213[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_214 = {1{$random}};
  reg_mip_msip = GEN_214[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_215 = {1{$random}};
  reg_mip_hsip = GEN_215[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_216 = {1{$random}};
  reg_mip_ssip = GEN_216[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_217 = {1{$random}};
  reg_mip_usip = GEN_217[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_218 = {2{$random}};
  reg_mepc = GEN_218[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_219 = {2{$random}};
  reg_mcause = GEN_219[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_220 = {2{$random}};
  reg_mbadaddr = GEN_220[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_221 = {2{$random}};
  reg_mscratch = GEN_221[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_222 = {1{$random}};
  reg_mtvec = GEN_222[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_223 = {1{$random}};
  reg_mucounteren = GEN_223[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_224 = {1{$random}};
  reg_mscounteren = GEN_224[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_225 = {2{$random}};
  reg_sepc = GEN_225[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_226 = {2{$random}};
  reg_scause = GEN_226[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_227 = {2{$random}};
  reg_sbadaddr = GEN_227[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_228 = {2{$random}};
  reg_sscratch = GEN_228[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_229 = {2{$random}};
  reg_stvec = GEN_229[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_230 = {1{$random}};
  reg_sptbr_asid = GEN_230[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_231 = {2{$random}};
  reg_sptbr_ppn = GEN_231[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_232 = {1{$random}};
  reg_wfi = GEN_232[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_233 = {1{$random}};
  reg_fflags = GEN_233[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_234 = {1{$random}};
  reg_frm = GEN_234[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_235 = {1{$random}};
  T_5570 = GEN_235[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_236 = {2{$random}};
  T_5573 = GEN_236[57:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_237 = {1{$random}};
  T_5581 = GEN_237[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_238 = {2{$random}};
  T_5584 = GEN_238[57:0];
  `endif
  GEN_239 = {1{$random}};
  GEN_240 = {1{$random}};
  GEN_241 = {1{$random}};
  GEN_242 = {1{$random}};
  GEN_243 = {1{$random}};
  GEN_244 = {1{$random}};
  GEN_245 = {1{$random}};
  GEN_246 = {1{$random}};
  GEN_247 = {1{$random}};
  GEN_248 = {2{$random}};
  GEN_249 = {2{$random}};
  GEN_250 = {1{$random}};
  GEN_251 = {1{$random}};
  GEN_252 = {1{$random}};
  GEN_253 = {1{$random}};
  GEN_254 = {1{$random}};
  GEN_255 = {1{$random}};
  GEN_256 = {1{$random}};
  GEN_257 = {1{$random}};
  GEN_258 = {1{$random}};
  GEN_259 = {1{$random}};
  GEN_260 = {1{$random}};
  GEN_261 = {1{$random}};
  GEN_262 = {1{$random}};
  GEN_263 = {1{$random}};
  GEN_264 = {1{$random}};
  GEN_265 = {1{$random}};
  GEN_266 = {1{$random}};
  GEN_267 = {1{$random}};
  GEN_268 = {1{$random}};
  GEN_269 = {1{$random}};
  GEN_270 = {1{$random}};
  GEN_271 = {1{$random}};
  GEN_272 = {1{$random}};
  GEN_273 = {1{$random}};
  GEN_274 = {1{$random}};
  GEN_275 = {1{$random}};
  GEN_276 = {1{$random}};
  GEN_277 = {1{$random}};
  GEN_278 = {2{$random}};
  GEN_279 = {1{$random}};
  GEN_280 = {1{$random}};
  GEN_281 = {1{$random}};
  GEN_282 = {2{$random}};
  GEN_283 = {1{$random}};
  GEN_284 = {1{$random}};
  GEN_285 = {2{$random}};
  GEN_286 = {2{$random}};
  GEN_287 = {1{$random}};
  GEN_288 = {1{$random}};
  GEN_289 = {1{$random}};
  GEN_290 = {1{$random}};
  GEN_291 = {1{$random}};
  GEN_292 = {1{$random}};
  GEN_293 = {1{$random}};
  GEN_294 = {1{$random}};
  GEN_295 = {1{$random}};
  GEN_296 = {1{$random}};
  GEN_297 = {1{$random}};
  GEN_298 = {1{$random}};
  GEN_299 = {1{$random}};
  GEN_300 = {2{$random}};
  GEN_301 = {1{$random}};
  GEN_302 = {1{$random}};
  GEN_303 = {3{$random}};
  GEN_304 = {1{$random}};
  GEN_305 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reg_mstatus_debug <= reset_mstatus_debug;
    end
    if(reset) begin
      reg_mstatus_prv <= reset_mstatus_prv;
    end else begin
      if(T_5084) begin
        reg_mstatus_prv <= 2'h0;
      end else begin
        reg_mstatus_prv <= new_prv;
      end
    end
    if(reset) begin
      reg_mstatus_sd <= reset_mstatus_sd;
    end
    if(reset) begin
      reg_mstatus_zero3 <= reset_mstatus_zero3;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= reset_mstatus_sd_rv32;
    end
    if(reset) begin
      reg_mstatus_zero2 <= reset_mstatus_zero2;
    end
    if(reset) begin
      reg_mstatus_vm <= reset_mstatus_vm;
    end else begin
      if(wen) begin
        if(T_6057) begin
          if(T_7129) begin
            reg_mstatus_vm <= 5'h9;
          end else begin
            if(T_7126) begin
              reg_mstatus_vm <= 5'h0;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_zero1 <= reset_mstatus_zero1;
    end
    if(reset) begin
      reg_mstatus_mxr <= reset_mstatus_mxr;
    end else begin
      if(wen) begin
        if(T_6057) begin
          reg_mstatus_mxr <= T_7074_mxr;
        end
      end
    end
    if(reset) begin
      reg_mstatus_pum <= reset_mstatus_pum;
    end else begin
      if(wen) begin
        if(T_6265) begin
          reg_mstatus_pum <= T_7330_pum;
        end else begin
          if(T_6057) begin
            reg_mstatus_pum <= T_7074_pum;
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_mprv <= reset_mstatus_mprv;
    end else begin
      if(wen) begin
        if(T_6057) begin
          reg_mstatus_mprv <= T_7074_mprv;
        end
      end
    end
    if(reset) begin
      reg_mstatus_xs <= reset_mstatus_xs;
    end
    if(reset) begin
      reg_mstatus_fs <= reset_mstatus_fs;
    end else begin
      if(wen) begin
        if(T_6265) begin
          if(T_7382) begin
            reg_mstatus_fs <= 2'h3;
          end else begin
            reg_mstatus_fs <= 2'h0;
          end
        end else begin
          if(T_6057) begin
            if(T_7132) begin
              reg_mstatus_fs <= 2'h3;
            end else begin
              reg_mstatus_fs <= 2'h0;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_mpp <= reset_mstatus_mpp;
    end else begin
      if(wen) begin
        if(T_6057) begin
          reg_mstatus_mpp <= T_7074_mpp;
        end else begin
          if(insn_ret) begin
            if(T_6623) begin
              reg_mstatus_mpp <= 2'h0;
            end else begin
              if(exception) begin
                if(T_6604) begin
                  reg_mstatus_mpp <= reg_mstatus_prv;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6604) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6623) begin
            reg_mstatus_mpp <= 2'h0;
          end else begin
            if(exception) begin
              if(T_6604) begin
                reg_mstatus_mpp <= reg_mstatus_prv;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6604) begin
              reg_mstatus_mpp <= reg_mstatus_prv;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpp <= reset_mstatus_hpp;
    end
    if(reset) begin
      reg_mstatus_spp <= reset_mstatus_spp;
    end else begin
      reg_mstatus_spp <= GEN_737[0];
    end
    if(reset) begin
      reg_mstatus_mpie <= reset_mstatus_mpie;
    end else begin
      if(wen) begin
        if(T_6057) begin
          reg_mstatus_mpie <= T_7074_mpie;
        end else begin
          if(insn_ret) begin
            if(T_6623) begin
              reg_mstatus_mpie <= 1'h0;
            end else begin
              if(exception) begin
                if(T_6604) begin
                  reg_mstatus_mpie <= T_6566;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6604) begin
                reg_mstatus_mpie <= T_6566;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6623) begin
            reg_mstatus_mpie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6604) begin
                reg_mstatus_mpie <= T_6566;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6604) begin
              reg_mstatus_mpie <= T_6566;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpie <= reset_mstatus_hpie;
    end
    if(reset) begin
      reg_mstatus_spie <= reset_mstatus_spie;
    end else begin
      if(wen) begin
        if(T_6265) begin
          reg_mstatus_spie <= T_7330_spie;
        end else begin
          if(T_6057) begin
            reg_mstatus_spie <= T_7074_spie;
          end else begin
            if(insn_ret) begin
              if(T_6547) begin
                reg_mstatus_spie <= 1'h0;
              end else begin
                if(exception) begin
                  if(T_6597) begin
                    reg_mstatus_spie <= T_6566;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6597) begin
                  reg_mstatus_spie <= T_6566;
                end
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6547) begin
            reg_mstatus_spie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6597) begin
                reg_mstatus_spie <= T_6566;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6597) begin
              reg_mstatus_spie <= T_6566;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_upie <= reset_mstatus_upie;
    end
    if(reset) begin
      reg_mstatus_mie <= reset_mstatus_mie;
    end else begin
      if(wen) begin
        if(T_6057) begin
          reg_mstatus_mie <= T_7074_mie;
        end else begin
          if(insn_ret) begin
            if(T_6623) begin
              if(T_6624) begin
                reg_mstatus_mie <= reg_mstatus_mpie;
              end else begin
                if(exception) begin
                  if(T_6604) begin
                    reg_mstatus_mie <= 1'h0;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6604) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6604) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6623) begin
            if(T_6624) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end else begin
              if(exception) begin
                if(T_6604) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            reg_mstatus_mie <= GEN_352;
          end
        end else begin
          reg_mstatus_mie <= GEN_352;
        end
      end
    end
    if(reset) begin
      reg_mstatus_hie <= reset_mstatus_hie;
    end
    if(reset) begin
      reg_mstatus_sie <= reset_mstatus_sie;
    end else begin
      if(wen) begin
        if(T_6265) begin
          reg_mstatus_sie <= T_7330_sie;
        end else begin
          if(T_6057) begin
            reg_mstatus_sie <= T_7074_sie;
          end else begin
            if(insn_ret) begin
              if(T_6623) begin
                if(T_6630) begin
                  reg_mstatus_sie <= reg_mstatus_mpie;
                end else begin
                  if(T_6547) begin
                    if(reg_mstatus_spp) begin
                      reg_mstatus_sie <= reg_mstatus_spie;
                    end else begin
                      if(exception) begin
                        if(T_6597) begin
                          reg_mstatus_sie <= 1'h0;
                        end
                      end
                    end
                  end else begin
                    if(exception) begin
                      if(T_6597) begin
                        reg_mstatus_sie <= 1'h0;
                      end
                    end
                  end
                end
              end else begin
                if(T_6547) begin
                  if(reg_mstatus_spp) begin
                    reg_mstatus_sie <= reg_mstatus_spie;
                  end else begin
                    if(exception) begin
                      if(T_6597) begin
                        reg_mstatus_sie <= 1'h0;
                      end
                    end
                  end
                end else begin
                  if(exception) begin
                    if(T_6597) begin
                      reg_mstatus_sie <= 1'h0;
                    end
                  end
                end
              end
            end else begin
              reg_mstatus_sie <= GEN_345;
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6623) begin
            if(T_6630) begin
              reg_mstatus_sie <= reg_mstatus_mpie;
            end else begin
              if(T_6547) begin
                if(reg_mstatus_spp) begin
                  reg_mstatus_sie <= reg_mstatus_spie;
                end else begin
                  reg_mstatus_sie <= GEN_345;
                end
              end else begin
                reg_mstatus_sie <= GEN_345;
              end
            end
          end else begin
            if(T_6547) begin
              if(reg_mstatus_spp) begin
                reg_mstatus_sie <= reg_mstatus_spie;
              end else begin
                reg_mstatus_sie <= GEN_345;
              end
            end else begin
              reg_mstatus_sie <= GEN_345;
            end
          end
        end else begin
          reg_mstatus_sie <= GEN_345;
        end
      end
    end
    if(reset) begin
      reg_mstatus_uie <= reset_mstatus_uie;
    end
    if(reset) begin
      reg_dcsr_xdebugver <= reset_dcsr_xdebugver;
    end
    if(reset) begin
      reg_dcsr_ndreset <= reset_dcsr_ndreset;
    end
    if(reset) begin
      reg_dcsr_fullreset <= reset_dcsr_fullreset;
    end
    if(reset) begin
      reg_dcsr_zero3 <= reset_dcsr_zero3;
    end
    if(reset) begin
      reg_dcsr_ebreakm <= reset_dcsr_ebreakm;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_ebreakm <= T_7241_ebreakm;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreakh <= reset_dcsr_ebreakh;
    end
    if(reset) begin
      reg_dcsr_ebreaks <= reset_dcsr_ebreaks;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_ebreaks <= T_7241_ebreaks;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreaku <= reset_dcsr_ebreaku;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_ebreaku <= T_7241_ebreaku;
        end
      end
    end
    if(reset) begin
      reg_dcsr_zero2 <= reset_dcsr_zero2;
    end
    if(reset) begin
      reg_dcsr_stopcycle <= reset_dcsr_stopcycle;
    end
    if(reset) begin
      reg_dcsr_stoptime <= reset_dcsr_stoptime;
    end
    if(reset) begin
      reg_dcsr_cause <= reset_dcsr_cause;
    end else begin
      if(exception) begin
        if(T_6528) begin
          if(reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, T_6593};
          end
        end
      end
    end
    if(reset) begin
      reg_dcsr_debugint <= reset_dcsr_debugint;
    end else begin
      reg_dcsr_debugint <= io_prci_interrupts_debug;
    end
    if(reset) begin
      reg_dcsr_zero1 <= reset_dcsr_zero1;
    end
    if(reset) begin
      reg_dcsr_halt <= reset_dcsr_halt;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_halt <= T_7241_halt;
        end
      end
    end
    if(reset) begin
      reg_dcsr_step <= reset_dcsr_step;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_step <= T_7241_step;
        end
      end
    end
    if(reset) begin
      reg_dcsr_prv <= reset_dcsr_prv;
    end else begin
      if(wen) begin
        if(T_6079) begin
          reg_dcsr_prv <= T_7241_prv;
        end else begin
          if(exception) begin
            if(T_6528) begin
              reg_dcsr_prv <= reg_mstatus_prv;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6528) begin
            reg_dcsr_prv <= reg_mstatus_prv;
          end
        end
      end
    end
    if(reset) begin
      reg_debug <= 1'h0;
    end else begin
      if(insn_ret) begin
        if(T_6617) begin
          reg_debug <= 1'h0;
        end else begin
          if(exception) begin
            if(T_6528) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6528) begin
            reg_debug <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_dpc <= GEN_792[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6083) begin
          reg_dscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5323) begin
        reg_singleStepped <= 1'h0;
      end else begin
        if(T_5320) begin
          reg_singleStepped <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_tselect <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_ttype <= 4'h2;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_dmode <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7481) begin
            if(T_6041) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_dmode <= GEN_33;
              end else begin
                if(1'h0 == reg_tselect) begin
                  reg_bp_0_control_dmode <= GEN_19;
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_maskmax <= 6'h4;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_reserved <= 40'h0;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_action <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7481) begin
            if(T_6041) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_action <= GEN_34;
              end else begin
                if(1'h0 == reg_tselect) begin
                  reg_bp_0_control_action <= GEN_22;
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_chain <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_zero <= 2'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7481) begin
          if(T_6041) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_control_tmatch <= GEN_25;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7481) begin
          if(T_6041) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_control_m <= GEN_26;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7481) begin
          if(T_6041) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_control_s <= GEN_28;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7481) begin
          if(T_6041) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_control_u <= GEN_29;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_x <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7481) begin
            if(T_6041) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_x <= GEN_30;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_w <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7481) begin
            if(T_6041) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_w <= GEN_31;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_r <= 1'h0;
      end else begin
        if(wen) begin
          if(T_7481) begin
            if(T_6041) begin
              if(1'h0 == reg_tselect) begin
                reg_bp_0_control_r <= GEN_32;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_7481) begin
          if(T_6043) begin
            if(1'h0 == reg_tselect) begin
              reg_bp_0_address <= GEN_35;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_ttype <= T_7607_control_ttype;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_dmode <= T_7607_control_dmode;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_maskmax <= T_7607_control_maskmax;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_reserved <= T_7607_control_reserved;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_action <= T_7607_control_action;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_chain <= T_7607_control_chain;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_zero <= T_7607_control_zero;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_tmatch <= T_7607_control_tmatch;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_m <= T_7607_control_m;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_h <= T_7607_control_h;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_s <= T_7607_control_s;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_u <= T_7607_control_u;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_x <= T_7607_control_x;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_w <= T_7607_control_w;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_r <= T_7607_control_r;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_address <= T_7607_address;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6269) begin
          reg_mie <= T_7445;
        end else begin
          if(T_6063) begin
            reg_mie <= T_7192;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6065) begin
          reg_mideleg <= T_7456;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6067) begin
          reg_medeleg <= T_7457;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_meip <= io_prci_interrupts_meip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_seip <= io_prci_interrupts_seip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_mtip <= io_prci_interrupts_mtip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6061) begin
          reg_mip_stip <= T_7165_stip;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_msip <= io_prci_interrupts_msip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6267) begin
          reg_mip_ssip <= T_7415_ssip;
        end else begin
          if(T_6061) begin
            reg_mip_ssip <= T_7165_ssip;
          end
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mepc <= GEN_758[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6075) begin
          reg_mcause <= T_7200;
        end else begin
          if(exception) begin
            if(T_6604) begin
              if(T_6499) begin
                reg_mcause <= io_cause;
              end else begin
                reg_mcause <= {{60'd0}, T_6506};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6604) begin
            if(T_6499) begin
              reg_mcause <= io_cause;
            end else begin
              reg_mcause <= {{60'd0}, T_6506};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6073) begin
          reg_mbadaddr <= T_7201;
        end else begin
          if(exception) begin
            if(T_6604) begin
              if(T_6586) begin
                reg_mbadaddr <= io_badaddr;
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6604) begin
            if(T_6586) begin
              reg_mbadaddr <= io_badaddr;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6069) begin
          reg_mscratch <= wdata;
        end
      end
    end
    if(reset) begin
      reg_mtvec <= 32'h1010;
    end else begin
      reg_mtvec <= GEN_760[31:0];
    end
    if(1'h0) begin
    end else begin
      reg_mucounteren <= GEN_841[31:0];
    end
    if(1'h0) begin
    end else begin
      reg_mscounteren <= GEN_840[31:0];
    end
    if(1'h0) begin
    end else begin
      reg_sepc <= GEN_834[39:0];
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6273) begin
          reg_scause <= T_7200;
        end else begin
          if(exception) begin
            if(T_6597) begin
              if(T_6499) begin
                reg_scause <= io_cause;
              end else begin
                reg_scause <= {{60'd0}, T_6506};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6597) begin
            if(T_6499) begin
              reg_scause <= io_cause;
            end else begin
              reg_scause <= {{60'd0}, T_6506};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6275) begin
          reg_sbadaddr <= T_7201;
        end else begin
          if(exception) begin
            if(T_6597) begin
              if(T_6586) begin
                reg_sbadaddr <= io_badaddr;
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6597) begin
            if(T_6586) begin
              reg_sbadaddr <= io_badaddr;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6271) begin
          reg_sscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_stvec <= GEN_835[38:0];
    end
    if(1'h0) begin
    end else begin
      reg_sptbr_asid <= 7'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6277) begin
          reg_sptbr_ppn <= {{18'd0}, T_7446};
        end
      end
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if(T_6496) begin
        reg_wfi <= 1'h0;
      end else begin
        if(insn_wfi) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_fflags <= GEN_767[4:0];
    end
    if(1'h0) begin
    end else begin
      reg_frm <= GEN_768[2:0];
    end
    if(reset) begin
      T_5570 <= 6'h0;
    end else begin
      T_5570 <= GEN_765[5:0];
    end
    if(reset) begin
      T_5573 <= 58'h0;
    end else begin
      if(wen) begin
        if(T_6053) begin
          T_5573 <= T_7202;
        end else begin
          if(T_5574) begin
            T_5573 <= T_5577;
          end
        end
      end else begin
        if(T_5574) begin
          T_5573 <= T_5577;
        end
      end
    end
    if(reset) begin
      T_5581 <= 6'h0;
    end else begin
      T_5581 <= GEN_763[5:0];
    end
    if(reset) begin
      T_5584 <= 58'h0;
    end else begin
      if(wen) begin
        if(T_6051) begin
          T_5584 <= T_7202;
        end else begin
          if(T_5585) begin
            T_5584 <= T_5588;
          end
        end
      end else begin
        if(T_5585) begin
          T_5584 <= T_5588;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:204 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_5340) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:205 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_5340) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6643) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at csr.scala:478 assert(PopCount(insn_ret :: io.exception :: io.csr_xcpt :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_6643) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BreakpointUnit(
  input   clk,
  input   reset,
  input   io_status_debug,
  input  [1:0] io_status_prv,
  input   io_status_sd,
  input  [30:0] io_status_zero3,
  input   io_status_sd_rv32,
  input  [1:0] io_status_zero2,
  input  [4:0] io_status_vm,
  input  [3:0] io_status_zero1,
  input   io_status_mxr,
  input   io_status_pum,
  input   io_status_mprv,
  input  [1:0] io_status_xs,
  input  [1:0] io_status_fs,
  input  [1:0] io_status_mpp,
  input  [1:0] io_status_hpp,
  input   io_status_spp,
  input   io_status_mpie,
  input   io_status_hpie,
  input   io_status_spie,
  input   io_status_upie,
  input   io_status_mie,
  input   io_status_hie,
  input   io_status_sie,
  input   io_status_uie,
  input  [3:0] io_bp_0_control_ttype,
  input   io_bp_0_control_dmode,
  input  [5:0] io_bp_0_control_maskmax,
  input  [39:0] io_bp_0_control_reserved,
  input   io_bp_0_control_action,
  input   io_bp_0_control_chain,
  input  [1:0] io_bp_0_control_zero,
  input  [1:0] io_bp_0_control_tmatch,
  input   io_bp_0_control_m,
  input   io_bp_0_control_h,
  input   io_bp_0_control_s,
  input   io_bp_0_control_u,
  input   io_bp_0_control_x,
  input   io_bp_0_control_w,
  input   io_bp_0_control_r,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output  io_xcpt_if,
  output  io_xcpt_ld,
  output  io_xcpt_st,
  output  io_debug_if,
  output  io_debug_ld,
  output  io_debug_st
);
  wire  T_212;
  wire [1:0] T_213;
  wire [1:0] T_214;
  wire [3:0] T_215;
  wire [3:0] T_216;
  wire  T_217;
  wire  T_218;
  wire  T_220;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire  T_224;
  wire [38:0] T_225;
  wire  T_227;
  wire  T_228;
  wire  T_229;
  wire  T_230;
  wire  T_231;
  wire  T_232;
  wire [1:0] T_233;
  wire [1:0] T_234;
  wire [3:0] T_235;
  wire [38:0] GEN_6;
  wire [38:0] T_236;
  wire [38:0] T_237;
  wire [38:0] T_248;
  wire  T_249;
  wire  T_250;
  wire  T_251;
  wire  T_253;
  wire  T_284;
  wire  T_286;
  wire  T_288;
  wire  T_290;
  wire [38:0] T_291;
  wire [38:0] T_302;
  wire  T_315;
  wire  T_316;
  wire  T_317;
  wire  T_319;
  wire  T_320;
  wire  T_322;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_323;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_326;
  wire  GEN_4;
  wire  GEN_5;
  assign io_xcpt_if = GEN_4;
  assign io_xcpt_ld = GEN_0;
  assign io_xcpt_st = GEN_2;
  assign io_debug_if = GEN_5;
  assign io_debug_ld = GEN_1;
  assign io_debug_st = GEN_3;
  assign T_212 = io_status_debug == 1'h0;
  assign T_213 = {io_bp_0_control_s,io_bp_0_control_u};
  assign T_214 = {io_bp_0_control_m,io_bp_0_control_h};
  assign T_215 = {T_214,T_213};
  assign T_216 = T_215 >> io_status_prv;
  assign T_217 = T_216[0];
  assign T_218 = T_212 & T_217;
  assign T_220 = T_218 & io_bp_0_control_r;
  assign T_221 = io_bp_0_control_tmatch[1];
  assign T_222 = io_ea >= io_bp_0_address;
  assign T_223 = io_bp_0_control_tmatch[0];
  assign T_224 = T_222 ^ T_223;
  assign T_225 = ~ io_ea;
  assign T_227 = io_bp_0_address[0];
  assign T_228 = T_223 & T_227;
  assign T_229 = io_bp_0_address[1];
  assign T_230 = T_228 & T_229;
  assign T_231 = io_bp_0_address[2];
  assign T_232 = T_230 & T_231;
  assign T_233 = {T_228,T_223};
  assign T_234 = {T_232,T_230};
  assign T_235 = {T_234,T_233};
  assign GEN_6 = {{35'd0}, T_235};
  assign T_236 = T_225 | GEN_6;
  assign T_237 = ~ io_bp_0_address;
  assign T_248 = T_237 | GEN_6;
  assign T_249 = T_236 == T_248;
  assign T_250 = T_221 ? T_224 : T_249;
  assign T_251 = T_220 & T_250;
  assign T_253 = T_218 & io_bp_0_control_w;
  assign T_284 = T_253 & T_250;
  assign T_286 = T_218 & io_bp_0_control_x;
  assign T_288 = io_pc >= io_bp_0_address;
  assign T_290 = T_288 ^ T_223;
  assign T_291 = ~ io_pc;
  assign T_302 = T_291 | GEN_6;
  assign T_315 = T_302 == T_248;
  assign T_316 = T_221 ? T_290 : T_315;
  assign T_317 = T_286 & T_316;
  assign T_319 = io_bp_0_control_chain == 1'h0;
  assign T_320 = T_319 & T_251;
  assign T_322 = io_bp_0_control_action == 1'h0;
  assign GEN_0 = T_320 ? T_322 : 1'h0;
  assign GEN_1 = T_320 ? io_bp_0_control_action : 1'h0;
  assign T_323 = T_319 & T_284;
  assign GEN_2 = T_323 ? T_322 : 1'h0;
  assign GEN_3 = T_323 ? io_bp_0_control_action : 1'h0;
  assign T_326 = T_319 & T_317;
  assign GEN_4 = T_326 ? T_322 : 1'h0;
  assign GEN_5 = T_326 ? io_bp_0_control_action : 1'h0;
endmodule
module ALU(
  input   clk,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_7;
  wire [63:0] T_8;
  wire [63:0] in2_inv;
  wire [63:0] in1_xor_in2;
  wire [64:0] T_9;
  wire [63:0] T_10;
  wire [63:0] GEN_1;
  wire [64:0] T_12;
  wire [63:0] T_13;
  wire  T_14;
  wire  T_17;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_30;
  wire  T_32;
  wire  T_33;
  wire [31:0] T_37;
  wire [31:0] T_39;
  wire [31:0] T_40;
  wire  T_41;
  wire  T_43;
  wire [4:0] T_44;
  wire [5:0] shamt;
  wire [31:0] T_45;
  wire [63:0] shin_r;
  wire  T_46;
  wire  T_47;
  wire  T_48;
  wire [31:0] T_53;
  wire [63:0] T_54;
  wire [31:0] T_55;
  wire [63:0] GEN_2;
  wire [63:0] T_56;
  wire [63:0] T_58;
  wire [63:0] T_59;
  wire [47:0] T_63;
  wire [63:0] GEN_3;
  wire [63:0] T_64;
  wire [47:0] T_65;
  wire [63:0] GEN_4;
  wire [63:0] T_66;
  wire [63:0] T_68;
  wire [63:0] T_69;
  wire [55:0] T_73;
  wire [63:0] GEN_5;
  wire [63:0] T_74;
  wire [55:0] T_75;
  wire [63:0] GEN_6;
  wire [63:0] T_76;
  wire [63:0] T_78;
  wire [63:0] T_79;
  wire [59:0] T_83;
  wire [63:0] GEN_7;
  wire [63:0] T_84;
  wire [59:0] T_85;
  wire [63:0] GEN_8;
  wire [63:0] T_86;
  wire [63:0] T_88;
  wire [63:0] T_89;
  wire [61:0] T_93;
  wire [63:0] GEN_9;
  wire [63:0] T_94;
  wire [61:0] T_95;
  wire [63:0] GEN_10;
  wire [63:0] T_96;
  wire [63:0] T_98;
  wire [63:0] T_99;
  wire [62:0] T_103;
  wire [63:0] GEN_11;
  wire [63:0] T_104;
  wire [62:0] T_105;
  wire [63:0] GEN_12;
  wire [63:0] T_106;
  wire [63:0] T_108;
  wire [63:0] T_109;
  wire [63:0] shin;
  wire  T_111;
  wire  T_112;
  wire [64:0] T_113;
  wire [64:0] T_114;
  wire [64:0] T_115;
  wire [63:0] shout_r;
  wire [31:0] T_120;
  wire [63:0] T_121;
  wire [31:0] T_122;
  wire [63:0] GEN_13;
  wire [63:0] T_123;
  wire [63:0] T_125;
  wire [63:0] T_126;
  wire [47:0] T_130;
  wire [63:0] GEN_14;
  wire [63:0] T_131;
  wire [47:0] T_132;
  wire [63:0] GEN_15;
  wire [63:0] T_133;
  wire [63:0] T_135;
  wire [63:0] T_136;
  wire [55:0] T_140;
  wire [63:0] GEN_16;
  wire [63:0] T_141;
  wire [55:0] T_142;
  wire [63:0] GEN_17;
  wire [63:0] T_143;
  wire [63:0] T_145;
  wire [63:0] T_146;
  wire [59:0] T_150;
  wire [63:0] GEN_18;
  wire [63:0] T_151;
  wire [59:0] T_152;
  wire [63:0] GEN_19;
  wire [63:0] T_153;
  wire [63:0] T_155;
  wire [63:0] T_156;
  wire [61:0] T_160;
  wire [63:0] GEN_20;
  wire [63:0] T_161;
  wire [61:0] T_162;
  wire [63:0] GEN_21;
  wire [63:0] T_163;
  wire [63:0] T_165;
  wire [63:0] T_166;
  wire [62:0] T_170;
  wire [63:0] GEN_22;
  wire [63:0] T_171;
  wire [62:0] T_172;
  wire [63:0] GEN_23;
  wire [63:0] T_173;
  wire [63:0] T_175;
  wire [63:0] shout_l;
  wire [63:0] T_180;
  wire  T_181;
  wire [63:0] T_183;
  wire [63:0] shout;
  wire  T_184;
  wire  T_185;
  wire  T_186;
  wire [63:0] T_188;
  wire  T_190;
  wire  T_191;
  wire [63:0] T_192;
  wire [63:0] T_194;
  wire [63:0] logic$;
  wire  T_195;
  wire  T_196;
  wire  T_197;
  wire  T_198;
  wire  T_199;
  wire  T_200;
  wire [63:0] GEN_24;
  wire [63:0] T_201;
  wire [63:0] shift_logic;
  wire  T_202;
  wire  T_203;
  wire  T_204;
  wire [63:0] out;
  wire  T_205;
  wire  T_206;
  wire [31:0] T_210;
  wire [31:0] T_211;
  wire [63:0] T_212;
  wire [63:0] GEN_0;
  assign io_out = GEN_0;
  assign io_adder_out = T_13;
  assign io_cmp_out = T_30;
  assign T_7 = io_fn[3];
  assign T_8 = ~ io_in2;
  assign in2_inv = T_7 ? T_8 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_9 = io_in1 + in2_inv;
  assign T_10 = T_9[63:0];
  assign GEN_1 = {{63'd0}, T_7};
  assign T_12 = T_10 + GEN_1;
  assign T_13 = T_12[63:0];
  assign T_14 = io_fn[0];
  assign T_17 = T_7 == 1'h0;
  assign T_19 = in1_xor_in2 == 64'h0;
  assign T_20 = io_in1[63];
  assign T_21 = io_in2[63];
  assign T_22 = T_20 == T_21;
  assign T_23 = io_adder_out[63];
  assign T_24 = io_fn[1];
  assign T_27 = T_24 ? T_21 : T_20;
  assign T_28 = T_22 ? T_23 : T_27;
  assign T_29 = T_17 ? T_19 : T_28;
  assign T_30 = T_14 ^ T_29;
  assign T_32 = io_in1[31];
  assign T_33 = T_7 & T_32;
  assign T_37 = T_33 ? 32'hffffffff : 32'h0;
  assign T_39 = io_in1[63:32];
  assign T_40 = io_dw ? T_39 : T_37;
  assign T_41 = io_in2[5];
  assign T_43 = T_41 & io_dw;
  assign T_44 = io_in2[4:0];
  assign shamt = {T_43,T_44};
  assign T_45 = io_in1[31:0];
  assign shin_r = {T_40,T_45};
  assign T_46 = io_fn == 4'h5;
  assign T_47 = io_fn == 4'hb;
  assign T_48 = T_46 | T_47;
  assign T_53 = shin_r[63:32];
  assign T_54 = {{32'd0}, T_53};
  assign T_55 = shin_r[31:0];
  assign GEN_2 = {{32'd0}, T_55};
  assign T_56 = GEN_2 << 32;
  assign T_58 = T_56 & 64'hffffffff00000000;
  assign T_59 = T_54 | T_58;
  assign T_63 = T_59[63:16];
  assign GEN_3 = {{16'd0}, T_63};
  assign T_64 = GEN_3 & 64'hffff0000ffff;
  assign T_65 = T_59[47:0];
  assign GEN_4 = {{16'd0}, T_65};
  assign T_66 = GEN_4 << 16;
  assign T_68 = T_66 & 64'hffff0000ffff0000;
  assign T_69 = T_64 | T_68;
  assign T_73 = T_69[63:8];
  assign GEN_5 = {{8'd0}, T_73};
  assign T_74 = GEN_5 & 64'hff00ff00ff00ff;
  assign T_75 = T_69[55:0];
  assign GEN_6 = {{8'd0}, T_75};
  assign T_76 = GEN_6 << 8;
  assign T_78 = T_76 & 64'hff00ff00ff00ff00;
  assign T_79 = T_74 | T_78;
  assign T_83 = T_79[63:4];
  assign GEN_7 = {{4'd0}, T_83};
  assign T_84 = GEN_7 & 64'hf0f0f0f0f0f0f0f;
  assign T_85 = T_79[59:0];
  assign GEN_8 = {{4'd0}, T_85};
  assign T_86 = GEN_8 << 4;
  assign T_88 = T_86 & 64'hf0f0f0f0f0f0f0f0;
  assign T_89 = T_84 | T_88;
  assign T_93 = T_89[63:2];
  assign GEN_9 = {{2'd0}, T_93};
  assign T_94 = GEN_9 & 64'h3333333333333333;
  assign T_95 = T_89[61:0];
  assign GEN_10 = {{2'd0}, T_95};
  assign T_96 = GEN_10 << 2;
  assign T_98 = T_96 & 64'hcccccccccccccccc;
  assign T_99 = T_94 | T_98;
  assign T_103 = T_99[63:1];
  assign GEN_11 = {{1'd0}, T_103};
  assign T_104 = GEN_11 & 64'h5555555555555555;
  assign T_105 = T_99[62:0];
  assign GEN_12 = {{1'd0}, T_105};
  assign T_106 = GEN_12 << 1;
  assign T_108 = T_106 & 64'haaaaaaaaaaaaaaaa;
  assign T_109 = T_104 | T_108;
  assign shin = T_48 ? shin_r : T_109;
  assign T_111 = shin[63];
  assign T_112 = T_7 & T_111;
  assign T_113 = {T_112,shin};
  assign T_114 = $signed(T_113);
  assign T_115 = $signed(T_114) >>> shamt;
  assign shout_r = T_115[63:0];
  assign T_120 = shout_r[63:32];
  assign T_121 = {{32'd0}, T_120};
  assign T_122 = shout_r[31:0];
  assign GEN_13 = {{32'd0}, T_122};
  assign T_123 = GEN_13 << 32;
  assign T_125 = T_123 & 64'hffffffff00000000;
  assign T_126 = T_121 | T_125;
  assign T_130 = T_126[63:16];
  assign GEN_14 = {{16'd0}, T_130};
  assign T_131 = GEN_14 & 64'hffff0000ffff;
  assign T_132 = T_126[47:0];
  assign GEN_15 = {{16'd0}, T_132};
  assign T_133 = GEN_15 << 16;
  assign T_135 = T_133 & 64'hffff0000ffff0000;
  assign T_136 = T_131 | T_135;
  assign T_140 = T_136[63:8];
  assign GEN_16 = {{8'd0}, T_140};
  assign T_141 = GEN_16 & 64'hff00ff00ff00ff;
  assign T_142 = T_136[55:0];
  assign GEN_17 = {{8'd0}, T_142};
  assign T_143 = GEN_17 << 8;
  assign T_145 = T_143 & 64'hff00ff00ff00ff00;
  assign T_146 = T_141 | T_145;
  assign T_150 = T_146[63:4];
  assign GEN_18 = {{4'd0}, T_150};
  assign T_151 = GEN_18 & 64'hf0f0f0f0f0f0f0f;
  assign T_152 = T_146[59:0];
  assign GEN_19 = {{4'd0}, T_152};
  assign T_153 = GEN_19 << 4;
  assign T_155 = T_153 & 64'hf0f0f0f0f0f0f0f0;
  assign T_156 = T_151 | T_155;
  assign T_160 = T_156[63:2];
  assign GEN_20 = {{2'd0}, T_160};
  assign T_161 = GEN_20 & 64'h3333333333333333;
  assign T_162 = T_156[61:0];
  assign GEN_21 = {{2'd0}, T_162};
  assign T_163 = GEN_21 << 2;
  assign T_165 = T_163 & 64'hcccccccccccccccc;
  assign T_166 = T_161 | T_165;
  assign T_170 = T_166[63:1];
  assign GEN_22 = {{1'd0}, T_170};
  assign T_171 = GEN_22 & 64'h5555555555555555;
  assign T_172 = T_166[62:0];
  assign GEN_23 = {{1'd0}, T_172};
  assign T_173 = GEN_23 << 1;
  assign T_175 = T_173 & 64'haaaaaaaaaaaaaaaa;
  assign shout_l = T_171 | T_175;
  assign T_180 = T_48 ? shout_r : 64'h0;
  assign T_181 = io_fn == 4'h1;
  assign T_183 = T_181 ? shout_l : 64'h0;
  assign shout = T_180 | T_183;
  assign T_184 = io_fn == 4'h4;
  assign T_185 = io_fn == 4'h6;
  assign T_186 = T_184 | T_185;
  assign T_188 = T_186 ? in1_xor_in2 : 64'h0;
  assign T_190 = io_fn == 4'h7;
  assign T_191 = T_185 | T_190;
  assign T_192 = io_in1 & io_in2;
  assign T_194 = T_191 ? T_192 : 64'h0;
  assign logic$ = T_188 | T_194;
  assign T_195 = io_fn == 4'h2;
  assign T_196 = io_fn == 4'h3;
  assign T_197 = T_195 | T_196;
  assign T_198 = io_fn >= 4'hc;
  assign T_199 = T_197 | T_198;
  assign T_200 = T_199 & io_cmp_out;
  assign GEN_24 = {{63'd0}, T_200};
  assign T_201 = GEN_24 | logic$;
  assign shift_logic = T_201 | shout;
  assign T_202 = io_fn == 4'h0;
  assign T_203 = io_fn == 4'ha;
  assign T_204 = T_202 | T_203;
  assign out = T_204 ? io_adder_out : shift_logic;
  assign T_205 = io_dw == 1'h0;
  assign T_206 = out[31];
  assign T_210 = T_206 ? 32'hffffffff : 32'h0;
  assign T_211 = out[31:0];
  assign T_212 = {T_210,T_211};
  assign GEN_0 = T_205 ? T_212 : out;
endmodule
module MulDiv(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [3:0] io_req_bits_fn,
  input   io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0] io_req_bits_tag,
  input   io_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] GEN_37;
  reg [3:0] req_fn;
  reg [31:0] GEN_38;
  reg  req_dw;
  reg [31:0] GEN_39;
  reg [63:0] req_in1;
  reg [63:0] GEN_40;
  reg [63:0] req_in2;
  reg [63:0] GEN_41;
  reg [4:0] req_tag;
  reg [31:0] GEN_42;
  reg [6:0] count;
  reg [31:0] GEN_43;
  reg  neg_out;
  reg [31:0] GEN_44;
  reg  isMul;
  reg [31:0] GEN_45;
  reg  isHi;
  reg [31:0] GEN_46;
  reg [64:0] divisor;
  reg [95:0] GEN_47;
  reg [129:0] remainder;
  reg [159:0] GEN_48;
  wire [3:0] T_62;
  wire  T_64;
  wire [3:0] T_66;
  wire  T_68;
  wire  T_71;
  wire [3:0] T_73;
  wire  T_75;
  wire [3:0] T_77;
  wire  T_79;
  wire  T_82;
  wire  T_83;
  wire [3:0] T_85;
  wire  T_87;
  wire [3:0] T_89;
  wire  T_91;
  wire  T_94;
  wire  T_95;
  wire  T_100;
  wire  T_102;
  wire  T_103;
  wire  T_104;
  wire  lhs_sign;
  wire [31:0] T_108;
  wire [31:0] T_109;
  wire [31:0] T_110;
  wire [31:0] T_111;
  wire [63:0] lhs_in;
  wire  T_115;
  wire  T_116;
  wire  T_117;
  wire  rhs_sign;
  wire [31:0] T_121;
  wire [31:0] T_122;
  wire [31:0] T_123;
  wire [31:0] T_124;
  wire [63:0] rhs_in;
  wire [64:0] T_125;
  wire [65:0] T_127;
  wire [64:0] subtractor;
  wire  less;
  wire [63:0] T_128;
  wire [64:0] T_130;
  wire [63:0] negated_remainder;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [129:0] GEN_0;
  wire  T_134;
  wire  T_135;
  wire [64:0] GEN_1;
  wire [129:0] GEN_2;
  wire [64:0] GEN_3;
  wire [2:0] GEN_4;
  wire  T_136;
  wire [129:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_137;
  wire [63:0] T_138;
  wire [2:0] T_139;
  wire [129:0] GEN_7;
  wire [2:0] GEN_8;
  wire  T_140;
  wire  T_141;
  wire [64:0] T_142;
  wire [128:0] T_144;
  wire [63:0] T_145;
  wire [64:0] T_146;
  wire [64:0] T_147;
  wire [64:0] T_148;
  wire [7:0] T_149;
  wire [64:0] GEN_34;
  wire [72:0] T_150;
  wire [72:0] GEN_35;
  wire [73:0] T_151;
  wire [72:0] T_152;
  wire [72:0] T_153;
  wire [55:0] T_154;
  wire [72:0] T_155;
  wire [128:0] T_156;
  wire [10:0] T_159;
  wire [5:0] T_160;
  wire [64:0] T_161;
  wire [63:0] T_162;
  wire  T_165;
  wire  T_168;
  wire  T_169;
  wire  T_171;
  wire  T_172;
  wire [63:0] T_173;
  wire [63:0] T_174;
  wire  T_176;
  wire  T_177;
  wire [11:0] T_181;
  wire [10:0] T_182;
  wire [5:0] T_183;
  wire [128:0] T_184;
  wire [64:0] T_185;
  wire [128:0] T_186;
  wire [63:0] T_187;
  wire [128:0] T_188;
  wire [64:0] T_189;
  wire [63:0] T_191;
  wire [65:0] T_192;
  wire [129:0] T_193;
  wire [7:0] T_195;
  wire [6:0] T_196;
  wire  T_198;
  wire  T_199;
  wire [2:0] T_200;
  wire [2:0] GEN_9;
  wire [129:0] GEN_10;
  wire [6:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_203;
  wire  T_204;
  wire  T_206;
  wire [2:0] T_208;
  wire [2:0] GEN_13;
  wire [63:0] T_212;
  wire [63:0] T_213;
  wire [63:0] T_214;
  wire  T_217;
  wire [127:0] T_218;
  wire [128:0] T_219;
  wire [63:0] T_220;
  wire [31:0] T_221;
  wire [31:0] T_222;
  wire  T_224;
  wire [15:0] T_225;
  wire [15:0] T_226;
  wire  T_228;
  wire [7:0] T_229;
  wire [7:0] T_230;
  wire  T_232;
  wire [3:0] T_233;
  wire [3:0] T_234;
  wire  T_236;
  wire  T_237;
  wire  T_239;
  wire  T_241;
  wire [1:0] T_243;
  wire [1:0] T_244;
  wire  T_245;
  wire  T_247;
  wire  T_249;
  wire [1:0] T_251;
  wire [1:0] T_252;
  wire [1:0] T_253;
  wire [2:0] T_254;
  wire [3:0] T_255;
  wire [3:0] T_256;
  wire  T_258;
  wire  T_259;
  wire  T_261;
  wire  T_263;
  wire [1:0] T_265;
  wire [1:0] T_266;
  wire  T_267;
  wire  T_269;
  wire  T_271;
  wire [1:0] T_273;
  wire [1:0] T_274;
  wire [1:0] T_275;
  wire [2:0] T_276;
  wire [2:0] T_277;
  wire [3:0] T_278;
  wire [7:0] T_279;
  wire [7:0] T_280;
  wire  T_282;
  wire [3:0] T_283;
  wire [3:0] T_284;
  wire  T_286;
  wire  T_287;
  wire  T_289;
  wire  T_291;
  wire [1:0] T_293;
  wire [1:0] T_294;
  wire  T_295;
  wire  T_297;
  wire  T_299;
  wire [1:0] T_301;
  wire [1:0] T_302;
  wire [1:0] T_303;
  wire [2:0] T_304;
  wire [3:0] T_305;
  wire [3:0] T_306;
  wire  T_308;
  wire  T_309;
  wire  T_311;
  wire  T_313;
  wire [1:0] T_315;
  wire [1:0] T_316;
  wire  T_317;
  wire  T_319;
  wire  T_321;
  wire [1:0] T_323;
  wire [1:0] T_324;
  wire [1:0] T_325;
  wire [2:0] T_326;
  wire [2:0] T_327;
  wire [3:0] T_328;
  wire [3:0] T_329;
  wire [4:0] T_330;
  wire [15:0] T_331;
  wire [15:0] T_332;
  wire  T_334;
  wire [7:0] T_335;
  wire [7:0] T_336;
  wire  T_338;
  wire [3:0] T_339;
  wire [3:0] T_340;
  wire  T_342;
  wire  T_343;
  wire  T_345;
  wire  T_347;
  wire [1:0] T_349;
  wire [1:0] T_350;
  wire  T_351;
  wire  T_353;
  wire  T_355;
  wire [1:0] T_357;
  wire [1:0] T_358;
  wire [1:0] T_359;
  wire [2:0] T_360;
  wire [3:0] T_361;
  wire [3:0] T_362;
  wire  T_364;
  wire  T_365;
  wire  T_367;
  wire  T_369;
  wire [1:0] T_371;
  wire [1:0] T_372;
  wire  T_373;
  wire  T_375;
  wire  T_377;
  wire [1:0] T_379;
  wire [1:0] T_380;
  wire [1:0] T_381;
  wire [2:0] T_382;
  wire [2:0] T_383;
  wire [3:0] T_384;
  wire [7:0] T_385;
  wire [7:0] T_386;
  wire  T_388;
  wire [3:0] T_389;
  wire [3:0] T_390;
  wire  T_392;
  wire  T_393;
  wire  T_395;
  wire  T_397;
  wire [1:0] T_399;
  wire [1:0] T_400;
  wire  T_401;
  wire  T_403;
  wire  T_405;
  wire [1:0] T_407;
  wire [1:0] T_408;
  wire [1:0] T_409;
  wire [2:0] T_410;
  wire [3:0] T_411;
  wire [3:0] T_412;
  wire  T_414;
  wire  T_415;
  wire  T_417;
  wire  T_419;
  wire [1:0] T_421;
  wire [1:0] T_422;
  wire  T_423;
  wire  T_425;
  wire  T_427;
  wire [1:0] T_429;
  wire [1:0] T_430;
  wire [1:0] T_431;
  wire [2:0] T_432;
  wire [2:0] T_433;
  wire [3:0] T_434;
  wire [3:0] T_435;
  wire [4:0] T_436;
  wire [4:0] T_437;
  wire [5:0] T_438;
  wire [31:0] T_440;
  wire [31:0] T_441;
  wire  T_443;
  wire [15:0] T_444;
  wire [15:0] T_445;
  wire  T_447;
  wire [7:0] T_448;
  wire [7:0] T_449;
  wire  T_451;
  wire [3:0] T_452;
  wire [3:0] T_453;
  wire  T_455;
  wire  T_456;
  wire  T_458;
  wire  T_460;
  wire [1:0] T_462;
  wire [1:0] T_463;
  wire  T_464;
  wire  T_466;
  wire  T_468;
  wire [1:0] T_470;
  wire [1:0] T_471;
  wire [1:0] T_472;
  wire [2:0] T_473;
  wire [3:0] T_474;
  wire [3:0] T_475;
  wire  T_477;
  wire  T_478;
  wire  T_480;
  wire  T_482;
  wire [1:0] T_484;
  wire [1:0] T_485;
  wire  T_486;
  wire  T_488;
  wire  T_490;
  wire [1:0] T_492;
  wire [1:0] T_493;
  wire [1:0] T_494;
  wire [2:0] T_495;
  wire [2:0] T_496;
  wire [3:0] T_497;
  wire [7:0] T_498;
  wire [7:0] T_499;
  wire  T_501;
  wire [3:0] T_502;
  wire [3:0] T_503;
  wire  T_505;
  wire  T_506;
  wire  T_508;
  wire  T_510;
  wire [1:0] T_512;
  wire [1:0] T_513;
  wire  T_514;
  wire  T_516;
  wire  T_518;
  wire [1:0] T_520;
  wire [1:0] T_521;
  wire [1:0] T_522;
  wire [2:0] T_523;
  wire [3:0] T_524;
  wire [3:0] T_525;
  wire  T_527;
  wire  T_528;
  wire  T_530;
  wire  T_532;
  wire [1:0] T_534;
  wire [1:0] T_535;
  wire  T_536;
  wire  T_538;
  wire  T_540;
  wire [1:0] T_542;
  wire [1:0] T_543;
  wire [1:0] T_544;
  wire [2:0] T_545;
  wire [2:0] T_546;
  wire [3:0] T_547;
  wire [3:0] T_548;
  wire [4:0] T_549;
  wire [15:0] T_550;
  wire [15:0] T_551;
  wire  T_553;
  wire [7:0] T_554;
  wire [7:0] T_555;
  wire  T_557;
  wire [3:0] T_558;
  wire [3:0] T_559;
  wire  T_561;
  wire  T_562;
  wire  T_564;
  wire  T_566;
  wire [1:0] T_568;
  wire [1:0] T_569;
  wire  T_570;
  wire  T_572;
  wire  T_574;
  wire [1:0] T_576;
  wire [1:0] T_577;
  wire [1:0] T_578;
  wire [2:0] T_579;
  wire [3:0] T_580;
  wire [3:0] T_581;
  wire  T_583;
  wire  T_584;
  wire  T_586;
  wire  T_588;
  wire [1:0] T_590;
  wire [1:0] T_591;
  wire  T_592;
  wire  T_594;
  wire  T_596;
  wire [1:0] T_598;
  wire [1:0] T_599;
  wire [1:0] T_600;
  wire [2:0] T_601;
  wire [2:0] T_602;
  wire [3:0] T_603;
  wire [7:0] T_604;
  wire [7:0] T_605;
  wire  T_607;
  wire [3:0] T_608;
  wire [3:0] T_609;
  wire  T_611;
  wire  T_612;
  wire  T_614;
  wire  T_616;
  wire [1:0] T_618;
  wire [1:0] T_619;
  wire  T_620;
  wire  T_622;
  wire  T_624;
  wire [1:0] T_626;
  wire [1:0] T_627;
  wire [1:0] T_628;
  wire [2:0] T_629;
  wire [3:0] T_630;
  wire [3:0] T_631;
  wire  T_633;
  wire  T_634;
  wire  T_636;
  wire  T_638;
  wire [1:0] T_640;
  wire [1:0] T_641;
  wire  T_642;
  wire  T_644;
  wire  T_646;
  wire [1:0] T_648;
  wire [1:0] T_649;
  wire [1:0] T_650;
  wire [2:0] T_651;
  wire [2:0] T_652;
  wire [3:0] T_653;
  wire [3:0] T_654;
  wire [4:0] T_655;
  wire [4:0] T_656;
  wire [5:0] T_657;
  wire [6:0] T_659;
  wire [5:0] T_660;
  wire [6:0] T_661;
  wire [5:0] T_662;
  wire  T_663;
  wire  T_665;
  wire  T_666;
  wire  T_668;
  wire  T_669;
  wire  T_670;
  wire [5:0] T_675;
  wire [126:0] GEN_36;
  wire [126:0] T_677;
  wire [128:0] GEN_14;
  wire [6:0] GEN_15;
  wire  T_682;
  wire  T_685;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [6:0] GEN_18;
  wire [129:0] GEN_19;
  wire  GEN_20;
  wire  T_687;
  wire  T_688;
  wire [2:0] GEN_21;
  wire  T_689;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire [2:0] T_694;
  wire  T_698;
  wire  T_699;
  wire  T_700;
  wire [64:0] T_701;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [6:0] GEN_25;
  wire  GEN_26;
  wire [64:0] GEN_27;
  wire [129:0] GEN_28;
  wire [3:0] GEN_29;
  wire  GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [4:0] GEN_33;
  wire  T_703;
  wire  T_705;
  wire [31:0] T_709;
  wire [31:0] T_710;
  wire [63:0] T_711;
  wire [63:0] T_713;
  wire  T_714;
  wire  T_715;
  assign io_req_ready = T_715;
  assign io_resp_valid = T_714;
  assign io_resp_bits_data = T_713;
  assign io_resp_bits_tag = req_tag;
  assign T_62 = io_req_bits_fn & 4'h4;
  assign T_64 = T_62 == 4'h0;
  assign T_66 = io_req_bits_fn & 4'h8;
  assign T_68 = T_66 == 4'h8;
  assign T_71 = T_64 | T_68;
  assign T_73 = io_req_bits_fn & 4'h5;
  assign T_75 = T_73 == 4'h1;
  assign T_77 = io_req_bits_fn & 4'h2;
  assign T_79 = T_77 == 4'h2;
  assign T_82 = T_75 | T_79;
  assign T_83 = T_82 | T_68;
  assign T_85 = io_req_bits_fn & 4'h9;
  assign T_87 = T_85 == 4'h0;
  assign T_89 = io_req_bits_fn & 4'h3;
  assign T_91 = T_89 == 4'h0;
  assign T_94 = T_87 | T_64;
  assign T_95 = T_94 | T_91;
  assign T_100 = io_req_bits_dw == 1'h0;
  assign T_102 = io_req_bits_in1[31];
  assign T_103 = io_req_bits_in1[63];
  assign T_104 = T_100 ? T_102 : T_103;
  assign lhs_sign = T_95 & T_104;
  assign T_108 = lhs_sign ? 32'hffffffff : 32'h0;
  assign T_109 = io_req_bits_in1[63:32];
  assign T_110 = T_100 ? T_108 : T_109;
  assign T_111 = io_req_bits_in1[31:0];
  assign lhs_in = {T_110,T_111};
  assign T_115 = io_req_bits_in2[31];
  assign T_116 = io_req_bits_in2[63];
  assign T_117 = T_100 ? T_115 : T_116;
  assign rhs_sign = T_94 & T_117;
  assign T_121 = rhs_sign ? 32'hffffffff : 32'h0;
  assign T_122 = io_req_bits_in2[63:32];
  assign T_123 = T_100 ? T_121 : T_122;
  assign T_124 = io_req_bits_in2[31:0];
  assign rhs_in = {T_123,T_124};
  assign T_125 = remainder[128:64];
  assign T_127 = T_125 - divisor;
  assign subtractor = T_127[64:0];
  assign less = subtractor[64];
  assign T_128 = remainder[63:0];
  assign T_130 = 64'h0 - T_128;
  assign negated_remainder = T_130[63:0];
  assign T_131 = state == 3'h1;
  assign T_132 = remainder[63];
  assign T_133 = T_132 | isMul;
  assign GEN_0 = T_133 ? {{66'd0}, negated_remainder} : remainder;
  assign T_134 = divisor[63];
  assign T_135 = T_134 | isMul;
  assign GEN_1 = T_135 ? subtractor : divisor;
  assign GEN_2 = T_131 ? GEN_0 : remainder;
  assign GEN_3 = T_131 ? GEN_1 : divisor;
  assign GEN_4 = T_131 ? 3'h2 : state;
  assign T_136 = state == 3'h4;
  assign GEN_5 = T_136 ? {{66'd0}, negated_remainder} : GEN_2;
  assign GEN_6 = T_136 ? 3'h5 : GEN_4;
  assign T_137 = state == 3'h3;
  assign T_138 = remainder[128:65];
  assign T_139 = neg_out ? 3'h4 : 3'h5;
  assign GEN_7 = T_137 ? {{66'd0}, T_138} : GEN_5;
  assign GEN_8 = T_137 ? T_139 : GEN_6;
  assign T_140 = state == 3'h2;
  assign T_141 = T_140 & isMul;
  assign T_142 = remainder[129:65];
  assign T_144 = {T_142,T_128};
  assign T_145 = T_144[63:0];
  assign T_146 = T_144[128:64];
  assign T_147 = $signed(T_146);
  assign T_148 = $signed(divisor);
  assign T_149 = T_145[7:0];
  assign GEN_34 = {{57'd0}, T_149};
  assign T_150 = $signed(T_148) * $signed({1'b0,GEN_34});
  assign GEN_35 = {{8{T_147[64]}},T_147};
  assign T_151 = $signed(T_150) + $signed(GEN_35);
  assign T_152 = T_151[72:0];
  assign T_153 = $signed(T_152);
  assign T_154 = T_145[63:8];
  assign T_155 = $unsigned(T_153);
  assign T_156 = {T_155,T_154};
  assign T_159 = count * 7'h8;
  assign T_160 = T_159[5:0];
  assign T_161 = $signed(65'sh10000000000000000) >>> T_160;
  assign T_162 = T_161[63:0];
  assign T_165 = count != 7'h7;
  assign T_168 = count != 7'h0;
  assign T_169 = T_165 & T_168;
  assign T_171 = isHi == 1'h0;
  assign T_172 = T_169 & T_171;
  assign T_173 = ~ T_162;
  assign T_174 = T_145 & T_173;
  assign T_176 = T_174 == 64'h0;
  assign T_177 = T_172 & T_176;
  assign T_181 = 11'h40 - T_159;
  assign T_182 = T_181[10:0];
  assign T_183 = T_182[5:0];
  assign T_184 = T_144 >> T_183;
  assign T_185 = T_156[128:64];
  assign T_186 = T_177 ? T_184 : T_156;
  assign T_187 = T_186[63:0];
  assign T_188 = {T_185,T_187};
  assign T_189 = T_188[128:64];
  assign T_191 = T_188[63:0];
  assign T_192 = {T_189,1'h0};
  assign T_193 = {T_192,T_191};
  assign T_195 = count + 7'h1;
  assign T_196 = T_195[6:0];
  assign T_198 = count == 7'h7;
  assign T_199 = T_177 | T_198;
  assign T_200 = isHi ? 3'h3 : 3'h5;
  assign GEN_9 = T_199 ? T_200 : GEN_8;
  assign GEN_10 = T_141 ? T_193 : GEN_7;
  assign GEN_11 = T_141 ? T_196 : count;
  assign GEN_12 = T_141 ? GEN_9 : GEN_8;
  assign T_203 = isMul == 1'h0;
  assign T_204 = T_140 & T_203;
  assign T_206 = count == 7'h40;
  assign T_208 = isHi ? 3'h3 : T_139;
  assign GEN_13 = T_206 ? T_208 : GEN_12;
  assign T_212 = remainder[127:64];
  assign T_213 = subtractor[63:0];
  assign T_214 = less ? T_212 : T_213;
  assign T_217 = less == 1'h0;
  assign T_218 = {T_214,T_128};
  assign T_219 = {T_218,T_217};
  assign T_220 = divisor[63:0];
  assign T_221 = T_220[63:32];
  assign T_222 = T_220[31:0];
  assign T_224 = T_221 != 32'h0;
  assign T_225 = T_221[31:16];
  assign T_226 = T_221[15:0];
  assign T_228 = T_225 != 16'h0;
  assign T_229 = T_225[15:8];
  assign T_230 = T_225[7:0];
  assign T_232 = T_229 != 8'h0;
  assign T_233 = T_229[7:4];
  assign T_234 = T_229[3:0];
  assign T_236 = T_233 != 4'h0;
  assign T_237 = T_233[3];
  assign T_239 = T_233[2];
  assign T_241 = T_233[1];
  assign T_243 = T_239 ? 2'h2 : {{1'd0}, T_241};
  assign T_244 = T_237 ? 2'h3 : T_243;
  assign T_245 = T_234[3];
  assign T_247 = T_234[2];
  assign T_249 = T_234[1];
  assign T_251 = T_247 ? 2'h2 : {{1'd0}, T_249};
  assign T_252 = T_245 ? 2'h3 : T_251;
  assign T_253 = T_236 ? T_244 : T_252;
  assign T_254 = {T_236,T_253};
  assign T_255 = T_230[7:4];
  assign T_256 = T_230[3:0];
  assign T_258 = T_255 != 4'h0;
  assign T_259 = T_255[3];
  assign T_261 = T_255[2];
  assign T_263 = T_255[1];
  assign T_265 = T_261 ? 2'h2 : {{1'd0}, T_263};
  assign T_266 = T_259 ? 2'h3 : T_265;
  assign T_267 = T_256[3];
  assign T_269 = T_256[2];
  assign T_271 = T_256[1];
  assign T_273 = T_269 ? 2'h2 : {{1'd0}, T_271};
  assign T_274 = T_267 ? 2'h3 : T_273;
  assign T_275 = T_258 ? T_266 : T_274;
  assign T_276 = {T_258,T_275};
  assign T_277 = T_232 ? T_254 : T_276;
  assign T_278 = {T_232,T_277};
  assign T_279 = T_226[15:8];
  assign T_280 = T_226[7:0];
  assign T_282 = T_279 != 8'h0;
  assign T_283 = T_279[7:4];
  assign T_284 = T_279[3:0];
  assign T_286 = T_283 != 4'h0;
  assign T_287 = T_283[3];
  assign T_289 = T_283[2];
  assign T_291 = T_283[1];
  assign T_293 = T_289 ? 2'h2 : {{1'd0}, T_291};
  assign T_294 = T_287 ? 2'h3 : T_293;
  assign T_295 = T_284[3];
  assign T_297 = T_284[2];
  assign T_299 = T_284[1];
  assign T_301 = T_297 ? 2'h2 : {{1'd0}, T_299};
  assign T_302 = T_295 ? 2'h3 : T_301;
  assign T_303 = T_286 ? T_294 : T_302;
  assign T_304 = {T_286,T_303};
  assign T_305 = T_280[7:4];
  assign T_306 = T_280[3:0];
  assign T_308 = T_305 != 4'h0;
  assign T_309 = T_305[3];
  assign T_311 = T_305[2];
  assign T_313 = T_305[1];
  assign T_315 = T_311 ? 2'h2 : {{1'd0}, T_313};
  assign T_316 = T_309 ? 2'h3 : T_315;
  assign T_317 = T_306[3];
  assign T_319 = T_306[2];
  assign T_321 = T_306[1];
  assign T_323 = T_319 ? 2'h2 : {{1'd0}, T_321};
  assign T_324 = T_317 ? 2'h3 : T_323;
  assign T_325 = T_308 ? T_316 : T_324;
  assign T_326 = {T_308,T_325};
  assign T_327 = T_282 ? T_304 : T_326;
  assign T_328 = {T_282,T_327};
  assign T_329 = T_228 ? T_278 : T_328;
  assign T_330 = {T_228,T_329};
  assign T_331 = T_222[31:16];
  assign T_332 = T_222[15:0];
  assign T_334 = T_331 != 16'h0;
  assign T_335 = T_331[15:8];
  assign T_336 = T_331[7:0];
  assign T_338 = T_335 != 8'h0;
  assign T_339 = T_335[7:4];
  assign T_340 = T_335[3:0];
  assign T_342 = T_339 != 4'h0;
  assign T_343 = T_339[3];
  assign T_345 = T_339[2];
  assign T_347 = T_339[1];
  assign T_349 = T_345 ? 2'h2 : {{1'd0}, T_347};
  assign T_350 = T_343 ? 2'h3 : T_349;
  assign T_351 = T_340[3];
  assign T_353 = T_340[2];
  assign T_355 = T_340[1];
  assign T_357 = T_353 ? 2'h2 : {{1'd0}, T_355};
  assign T_358 = T_351 ? 2'h3 : T_357;
  assign T_359 = T_342 ? T_350 : T_358;
  assign T_360 = {T_342,T_359};
  assign T_361 = T_336[7:4];
  assign T_362 = T_336[3:0];
  assign T_364 = T_361 != 4'h0;
  assign T_365 = T_361[3];
  assign T_367 = T_361[2];
  assign T_369 = T_361[1];
  assign T_371 = T_367 ? 2'h2 : {{1'd0}, T_369};
  assign T_372 = T_365 ? 2'h3 : T_371;
  assign T_373 = T_362[3];
  assign T_375 = T_362[2];
  assign T_377 = T_362[1];
  assign T_379 = T_375 ? 2'h2 : {{1'd0}, T_377};
  assign T_380 = T_373 ? 2'h3 : T_379;
  assign T_381 = T_364 ? T_372 : T_380;
  assign T_382 = {T_364,T_381};
  assign T_383 = T_338 ? T_360 : T_382;
  assign T_384 = {T_338,T_383};
  assign T_385 = T_332[15:8];
  assign T_386 = T_332[7:0];
  assign T_388 = T_385 != 8'h0;
  assign T_389 = T_385[7:4];
  assign T_390 = T_385[3:0];
  assign T_392 = T_389 != 4'h0;
  assign T_393 = T_389[3];
  assign T_395 = T_389[2];
  assign T_397 = T_389[1];
  assign T_399 = T_395 ? 2'h2 : {{1'd0}, T_397};
  assign T_400 = T_393 ? 2'h3 : T_399;
  assign T_401 = T_390[3];
  assign T_403 = T_390[2];
  assign T_405 = T_390[1];
  assign T_407 = T_403 ? 2'h2 : {{1'd0}, T_405};
  assign T_408 = T_401 ? 2'h3 : T_407;
  assign T_409 = T_392 ? T_400 : T_408;
  assign T_410 = {T_392,T_409};
  assign T_411 = T_386[7:4];
  assign T_412 = T_386[3:0];
  assign T_414 = T_411 != 4'h0;
  assign T_415 = T_411[3];
  assign T_417 = T_411[2];
  assign T_419 = T_411[1];
  assign T_421 = T_417 ? 2'h2 : {{1'd0}, T_419};
  assign T_422 = T_415 ? 2'h3 : T_421;
  assign T_423 = T_412[3];
  assign T_425 = T_412[2];
  assign T_427 = T_412[1];
  assign T_429 = T_425 ? 2'h2 : {{1'd0}, T_427};
  assign T_430 = T_423 ? 2'h3 : T_429;
  assign T_431 = T_414 ? T_422 : T_430;
  assign T_432 = {T_414,T_431};
  assign T_433 = T_388 ? T_410 : T_432;
  assign T_434 = {T_388,T_433};
  assign T_435 = T_334 ? T_384 : T_434;
  assign T_436 = {T_334,T_435};
  assign T_437 = T_224 ? T_330 : T_436;
  assign T_438 = {T_224,T_437};
  assign T_440 = T_128[63:32];
  assign T_441 = T_128[31:0];
  assign T_443 = T_440 != 32'h0;
  assign T_444 = T_440[31:16];
  assign T_445 = T_440[15:0];
  assign T_447 = T_444 != 16'h0;
  assign T_448 = T_444[15:8];
  assign T_449 = T_444[7:0];
  assign T_451 = T_448 != 8'h0;
  assign T_452 = T_448[7:4];
  assign T_453 = T_448[3:0];
  assign T_455 = T_452 != 4'h0;
  assign T_456 = T_452[3];
  assign T_458 = T_452[2];
  assign T_460 = T_452[1];
  assign T_462 = T_458 ? 2'h2 : {{1'd0}, T_460};
  assign T_463 = T_456 ? 2'h3 : T_462;
  assign T_464 = T_453[3];
  assign T_466 = T_453[2];
  assign T_468 = T_453[1];
  assign T_470 = T_466 ? 2'h2 : {{1'd0}, T_468};
  assign T_471 = T_464 ? 2'h3 : T_470;
  assign T_472 = T_455 ? T_463 : T_471;
  assign T_473 = {T_455,T_472};
  assign T_474 = T_449[7:4];
  assign T_475 = T_449[3:0];
  assign T_477 = T_474 != 4'h0;
  assign T_478 = T_474[3];
  assign T_480 = T_474[2];
  assign T_482 = T_474[1];
  assign T_484 = T_480 ? 2'h2 : {{1'd0}, T_482};
  assign T_485 = T_478 ? 2'h3 : T_484;
  assign T_486 = T_475[3];
  assign T_488 = T_475[2];
  assign T_490 = T_475[1];
  assign T_492 = T_488 ? 2'h2 : {{1'd0}, T_490};
  assign T_493 = T_486 ? 2'h3 : T_492;
  assign T_494 = T_477 ? T_485 : T_493;
  assign T_495 = {T_477,T_494};
  assign T_496 = T_451 ? T_473 : T_495;
  assign T_497 = {T_451,T_496};
  assign T_498 = T_445[15:8];
  assign T_499 = T_445[7:0];
  assign T_501 = T_498 != 8'h0;
  assign T_502 = T_498[7:4];
  assign T_503 = T_498[3:0];
  assign T_505 = T_502 != 4'h0;
  assign T_506 = T_502[3];
  assign T_508 = T_502[2];
  assign T_510 = T_502[1];
  assign T_512 = T_508 ? 2'h2 : {{1'd0}, T_510};
  assign T_513 = T_506 ? 2'h3 : T_512;
  assign T_514 = T_503[3];
  assign T_516 = T_503[2];
  assign T_518 = T_503[1];
  assign T_520 = T_516 ? 2'h2 : {{1'd0}, T_518};
  assign T_521 = T_514 ? 2'h3 : T_520;
  assign T_522 = T_505 ? T_513 : T_521;
  assign T_523 = {T_505,T_522};
  assign T_524 = T_499[7:4];
  assign T_525 = T_499[3:0];
  assign T_527 = T_524 != 4'h0;
  assign T_528 = T_524[3];
  assign T_530 = T_524[2];
  assign T_532 = T_524[1];
  assign T_534 = T_530 ? 2'h2 : {{1'd0}, T_532};
  assign T_535 = T_528 ? 2'h3 : T_534;
  assign T_536 = T_525[3];
  assign T_538 = T_525[2];
  assign T_540 = T_525[1];
  assign T_542 = T_538 ? 2'h2 : {{1'd0}, T_540};
  assign T_543 = T_536 ? 2'h3 : T_542;
  assign T_544 = T_527 ? T_535 : T_543;
  assign T_545 = {T_527,T_544};
  assign T_546 = T_501 ? T_523 : T_545;
  assign T_547 = {T_501,T_546};
  assign T_548 = T_447 ? T_497 : T_547;
  assign T_549 = {T_447,T_548};
  assign T_550 = T_441[31:16];
  assign T_551 = T_441[15:0];
  assign T_553 = T_550 != 16'h0;
  assign T_554 = T_550[15:8];
  assign T_555 = T_550[7:0];
  assign T_557 = T_554 != 8'h0;
  assign T_558 = T_554[7:4];
  assign T_559 = T_554[3:0];
  assign T_561 = T_558 != 4'h0;
  assign T_562 = T_558[3];
  assign T_564 = T_558[2];
  assign T_566 = T_558[1];
  assign T_568 = T_564 ? 2'h2 : {{1'd0}, T_566};
  assign T_569 = T_562 ? 2'h3 : T_568;
  assign T_570 = T_559[3];
  assign T_572 = T_559[2];
  assign T_574 = T_559[1];
  assign T_576 = T_572 ? 2'h2 : {{1'd0}, T_574};
  assign T_577 = T_570 ? 2'h3 : T_576;
  assign T_578 = T_561 ? T_569 : T_577;
  assign T_579 = {T_561,T_578};
  assign T_580 = T_555[7:4];
  assign T_581 = T_555[3:0];
  assign T_583 = T_580 != 4'h0;
  assign T_584 = T_580[3];
  assign T_586 = T_580[2];
  assign T_588 = T_580[1];
  assign T_590 = T_586 ? 2'h2 : {{1'd0}, T_588};
  assign T_591 = T_584 ? 2'h3 : T_590;
  assign T_592 = T_581[3];
  assign T_594 = T_581[2];
  assign T_596 = T_581[1];
  assign T_598 = T_594 ? 2'h2 : {{1'd0}, T_596};
  assign T_599 = T_592 ? 2'h3 : T_598;
  assign T_600 = T_583 ? T_591 : T_599;
  assign T_601 = {T_583,T_600};
  assign T_602 = T_557 ? T_579 : T_601;
  assign T_603 = {T_557,T_602};
  assign T_604 = T_551[15:8];
  assign T_605 = T_551[7:0];
  assign T_607 = T_604 != 8'h0;
  assign T_608 = T_604[7:4];
  assign T_609 = T_604[3:0];
  assign T_611 = T_608 != 4'h0;
  assign T_612 = T_608[3];
  assign T_614 = T_608[2];
  assign T_616 = T_608[1];
  assign T_618 = T_614 ? 2'h2 : {{1'd0}, T_616};
  assign T_619 = T_612 ? 2'h3 : T_618;
  assign T_620 = T_609[3];
  assign T_622 = T_609[2];
  assign T_624 = T_609[1];
  assign T_626 = T_622 ? 2'h2 : {{1'd0}, T_624};
  assign T_627 = T_620 ? 2'h3 : T_626;
  assign T_628 = T_611 ? T_619 : T_627;
  assign T_629 = {T_611,T_628};
  assign T_630 = T_605[7:4];
  assign T_631 = T_605[3:0];
  assign T_633 = T_630 != 4'h0;
  assign T_634 = T_630[3];
  assign T_636 = T_630[2];
  assign T_638 = T_630[1];
  assign T_640 = T_636 ? 2'h2 : {{1'd0}, T_638};
  assign T_641 = T_634 ? 2'h3 : T_640;
  assign T_642 = T_631[3];
  assign T_644 = T_631[2];
  assign T_646 = T_631[1];
  assign T_648 = T_644 ? 2'h2 : {{1'd0}, T_646};
  assign T_649 = T_642 ? 2'h3 : T_648;
  assign T_650 = T_633 ? T_641 : T_649;
  assign T_651 = {T_633,T_650};
  assign T_652 = T_607 ? T_629 : T_651;
  assign T_653 = {T_607,T_652};
  assign T_654 = T_553 ? T_603 : T_653;
  assign T_655 = {T_553,T_654};
  assign T_656 = T_443 ? T_549 : T_655;
  assign T_657 = {T_443,T_656};
  assign T_659 = 6'h3f + T_438;
  assign T_660 = T_659[5:0];
  assign T_661 = T_660 - T_657;
  assign T_662 = T_661[5:0];
  assign T_663 = T_438 > T_657;
  assign T_665 = count == 7'h0;
  assign T_666 = T_665 & less;
  assign T_668 = T_662 > 6'h0;
  assign T_669 = T_668 | T_663;
  assign T_670 = T_666 & T_669;
  assign T_675 = T_663 ? 6'h3f : T_662;
  assign GEN_36 = {{63'd0}, T_128};
  assign T_677 = GEN_36 << T_675;
  assign GEN_14 = T_670 ? {{2'd0}, T_677} : T_219;
  assign GEN_15 = T_670 ? {{1'd0}, T_675} : T_196;
  assign T_682 = T_665 & T_217;
  assign T_685 = T_682 & T_171;
  assign GEN_16 = T_685 ? 1'h0 : neg_out;
  assign GEN_17 = T_204 ? GEN_13 : GEN_12;
  assign GEN_18 = T_204 ? GEN_15 : GEN_11;
  assign GEN_19 = T_204 ? {{1'd0}, GEN_14} : GEN_10;
  assign GEN_20 = T_204 ? GEN_16 : neg_out;
  assign T_687 = io_resp_ready & io_resp_valid;
  assign T_688 = T_687 | io_kill;
  assign GEN_21 = T_688 ? 3'h0 : GEN_17;
  assign T_689 = io_req_ready & io_req_valid;
  assign T_691 = T_71 == 1'h0;
  assign T_692 = rhs_sign & T_691;
  assign T_693 = lhs_sign | T_692;
  assign T_694 = T_693 ? 3'h1 : 3'h2;
  assign T_698 = lhs_sign != rhs_sign;
  assign T_699 = T_83 ? lhs_sign : T_698;
  assign T_700 = T_691 & T_699;
  assign T_701 = {rhs_sign,rhs_in};
  assign GEN_22 = T_689 ? T_694 : GEN_21;
  assign GEN_23 = T_689 ? T_71 : isMul;
  assign GEN_24 = T_689 ? T_83 : isHi;
  assign GEN_25 = T_689 ? 7'h0 : GEN_18;
  assign GEN_26 = T_689 ? T_700 : GEN_20;
  assign GEN_27 = T_689 ? T_701 : GEN_3;
  assign GEN_28 = T_689 ? {{66'd0}, lhs_in} : GEN_19;
  assign GEN_29 = T_689 ? io_req_bits_fn : req_fn;
  assign GEN_30 = T_689 ? io_req_bits_dw : req_dw;
  assign GEN_31 = T_689 ? io_req_bits_in1 : req_in1;
  assign GEN_32 = T_689 ? io_req_bits_in2 : req_in2;
  assign GEN_33 = T_689 ? io_req_bits_tag : req_tag;
  assign T_703 = req_dw == 1'h0;
  assign T_705 = remainder[31];
  assign T_709 = T_705 ? 32'hffffffff : 32'h0;
  assign T_710 = remainder[31:0];
  assign T_711 = {T_709,T_710};
  assign T_713 = T_703 ? T_711 : T_128;
  assign T_714 = state == 3'h5;
  assign T_715 = state == 3'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  state = GEN_37[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  req_fn = GEN_38[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  req_dw = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {2{$random}};
  req_in1 = GEN_40[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {2{$random}};
  req_in2 = GEN_41[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  req_tag = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  count = GEN_43[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  neg_out = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  isMul = GEN_45[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  isHi = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {3{$random}};
  divisor = GEN_47[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {5{$random}};
  remainder = GEN_48[129:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_689) begin
        if(T_693) begin
          state <= 3'h1;
        end else begin
          state <= 3'h2;
        end
      end else begin
        if(T_688) begin
          state <= 3'h0;
        end else begin
          if(T_204) begin
            if(T_206) begin
              if(isHi) begin
                state <= 3'h3;
              end else begin
                if(neg_out) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h5;
                end
              end
            end else begin
              if(T_141) begin
                if(T_199) begin
                  if(isHi) begin
                    state <= 3'h3;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_137) begin
                    if(neg_out) begin
                      state <= 3'h4;
                    end else begin
                      state <= 3'h5;
                    end
                  end else begin
                    if(T_136) begin
                      state <= 3'h5;
                    end else begin
                      if(T_131) begin
                        state <= 3'h2;
                      end
                    end
                  end
                end
              end else begin
                if(T_137) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_136) begin
                    state <= 3'h5;
                  end else begin
                    if(T_131) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end
          end else begin
            if(T_141) begin
              if(T_199) begin
                if(isHi) begin
                  state <= 3'h3;
                end else begin
                  state <= 3'h5;
                end
              end else begin
                if(T_137) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_136) begin
                    state <= 3'h5;
                  end else begin
                    if(T_131) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(T_137) begin
                state <= T_139;
              end else begin
                if(T_136) begin
                  state <= 3'h5;
                end else begin
                  if(T_131) begin
                    state <= 3'h2;
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_fn <= io_req_bits_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_dw <= io_req_bits_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_in1 <= io_req_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_in2 <= io_req_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        count <= 7'h0;
      end else begin
        if(T_204) begin
          if(T_670) begin
            count <= {{1'd0}, T_675};
          end else begin
            count <= T_196;
          end
        end else begin
          if(T_141) begin
            count <= T_196;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        neg_out <= T_700;
      end else begin
        if(T_204) begin
          if(T_685) begin
            neg_out <= 1'h0;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        isMul <= T_71;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        isHi <= T_83;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        divisor <= T_701;
      end else begin
        if(T_131) begin
          if(T_135) begin
            divisor <= subtractor;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_689) begin
        remainder <= {{66'd0}, lhs_in};
      end else begin
        if(T_204) begin
          remainder <= {{1'd0}, GEN_14};
        end else begin
          if(T_141) begin
            remainder <= T_193;
          end else begin
            if(T_137) begin
              remainder <= {{66'd0}, T_138};
            end else begin
              if(T_136) begin
                remainder <= {{66'd0}, negated_remainder};
              end else begin
                if(T_131) begin
                  if(T_133) begin
                    remainder <= {{66'd0}, negated_remainder};
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Rocket(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  output  io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output  io_imem_req_bits_speculative,
  output  io_imem_resp_ready,
  input   io_imem_resp_valid,
  input   io_imem_resp_bits_btb_valid,
  input   io_imem_resp_bits_btb_bits_taken,
  input  [1:0] io_imem_resp_bits_btb_bits_mask,
  input   io_imem_resp_bits_btb_bits_bridx,
  input  [38:0] io_imem_resp_bits_btb_bits_target,
  input  [5:0] io_imem_resp_bits_btb_bits_entry,
  input  [6:0] io_imem_resp_bits_btb_bits_bht_history,
  input  [1:0] io_imem_resp_bits_btb_bits_bht_value,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input  [1:0] io_imem_resp_bits_mask,
  input   io_imem_resp_bits_xcpt_if,
  input   io_imem_resp_bits_replay,
  output  io_imem_btb_update_valid,
  output  io_imem_btb_update_bits_prediction_valid,
  output  io_imem_btb_update_bits_prediction_bits_taken,
  output [1:0] io_imem_btb_update_bits_prediction_bits_mask,
  output  io_imem_btb_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_btb_update_bits_prediction_bits_target,
  output [5:0] io_imem_btb_update_bits_prediction_bits_entry,
  output [6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_btb_update_bits_pc,
  output [38:0] io_imem_btb_update_bits_target,
  output  io_imem_btb_update_bits_taken,
  output  io_imem_btb_update_bits_isValid,
  output  io_imem_btb_update_bits_isJump,
  output  io_imem_btb_update_bits_isReturn,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output  io_imem_bht_update_valid,
  output  io_imem_bht_update_bits_prediction_valid,
  output  io_imem_bht_update_bits_prediction_bits_taken,
  output [1:0] io_imem_bht_update_bits_prediction_bits_mask,
  output  io_imem_bht_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_bht_update_bits_prediction_bits_target,
  output [5:0] io_imem_bht_update_bits_prediction_bits_entry,
  output [6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_bht_update_bits_pc,
  output  io_imem_bht_update_bits_taken,
  output  io_imem_bht_update_bits_mispredict,
  output  io_imem_ras_update_valid,
  output  io_imem_ras_update_bits_isCall,
  output  io_imem_ras_update_bits_isReturn,
  output [38:0] io_imem_ras_update_bits_returnAddr,
  output  io_imem_ras_update_bits_prediction_valid,
  output  io_imem_ras_update_bits_prediction_bits_taken,
  output [1:0] io_imem_ras_update_bits_prediction_bits_mask,
  output  io_imem_ras_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_ras_update_bits_prediction_bits_target,
  output [5:0] io_imem_ras_update_bits_prediction_bits_entry,
  output [6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
  output  io_imem_flush_icache,
  output  io_imem_flush_tlb,
  input  [39:0] io_imem_npc,
  input   io_dmem_req_ready,
  output  io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [6:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [2:0] io_dmem_req_bits_typ,
  output  io_dmem_req_bits_phys,
  output [63:0] io_dmem_req_bits_data,
  output  io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data,
  input   io_dmem_s2_nack,
  input   io_dmem_resp_valid,
  input  [39:0] io_dmem_resp_bits_addr,
  input  [6:0] io_dmem_resp_bits_tag,
  input  [4:0] io_dmem_resp_bits_cmd,
  input  [2:0] io_dmem_resp_bits_typ,
  input  [63:0] io_dmem_resp_bits_data,
  input   io_dmem_resp_bits_replay,
  input   io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input  [63:0] io_dmem_resp_bits_store_data,
  input   io_dmem_replay_next,
  input   io_dmem_xcpt_ma_ld,
  input   io_dmem_xcpt_ma_st,
  input   io_dmem_xcpt_pf_ld,
  input   io_dmem_xcpt_pf_st,
  output  io_dmem_invalidate_lr,
  input   io_dmem_ordered,
  output [6:0] io_ptw_ptbr_asid,
  output [37:0] io_ptw_ptbr_ppn,
  output  io_ptw_invalidate,
  output  io_ptw_status_debug,
  output [1:0] io_ptw_status_prv,
  output  io_ptw_status_sd,
  output [30:0] io_ptw_status_zero3,
  output  io_ptw_status_sd_rv32,
  output [1:0] io_ptw_status_zero2,
  output [4:0] io_ptw_status_vm,
  output [3:0] io_ptw_status_zero1,
  output  io_ptw_status_mxr,
  output  io_ptw_status_pum,
  output  io_ptw_status_mprv,
  output [1:0] io_ptw_status_xs,
  output [1:0] io_ptw_status_fs,
  output [1:0] io_ptw_status_mpp,
  output [1:0] io_ptw_status_hpp,
  output  io_ptw_status_spp,
  output  io_ptw_status_mpie,
  output  io_ptw_status_hpie,
  output  io_ptw_status_spie,
  output  io_ptw_status_upie,
  output  io_ptw_status_mie,
  output  io_ptw_status_hie,
  output  io_ptw_status_sie,
  output  io_ptw_status_uie,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input   io_fpu_fcsr_flags_valid,
  input  [4:0] io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output  io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output  io_fpu_valid,
  input   io_fpu_fcsr_rdy,
  input   io_fpu_nack_mem,
  input   io_fpu_illegal_rm,
  output  io_fpu_killx,
  output  io_fpu_killm,
  input  [4:0] io_fpu_dec_cmd,
  input   io_fpu_dec_ldst,
  input   io_fpu_dec_wen,
  input   io_fpu_dec_ren1,
  input   io_fpu_dec_ren2,
  input   io_fpu_dec_ren3,
  input   io_fpu_dec_swap12,
  input   io_fpu_dec_swap23,
  input   io_fpu_dec_single,
  input   io_fpu_dec_fromint,
  input   io_fpu_dec_toint,
  input   io_fpu_dec_fastpipe,
  input   io_fpu_dec_fma,
  input   io_fpu_dec_div,
  input   io_fpu_dec_sqrt,
  input   io_fpu_dec_round,
  input   io_fpu_dec_wflags,
  input   io_fpu_sboard_set,
  input   io_fpu_sboard_clr,
  input  [4:0] io_fpu_sboard_clra,
  input   io_fpu_cp_req_ready,
  output  io_fpu_cp_req_valid,
  output [4:0] io_fpu_cp_req_bits_cmd,
  output  io_fpu_cp_req_bits_ldst,
  output  io_fpu_cp_req_bits_wen,
  output  io_fpu_cp_req_bits_ren1,
  output  io_fpu_cp_req_bits_ren2,
  output  io_fpu_cp_req_bits_ren3,
  output  io_fpu_cp_req_bits_swap12,
  output  io_fpu_cp_req_bits_swap23,
  output  io_fpu_cp_req_bits_single,
  output  io_fpu_cp_req_bits_fromint,
  output  io_fpu_cp_req_bits_toint,
  output  io_fpu_cp_req_bits_fastpipe,
  output  io_fpu_cp_req_bits_fma,
  output  io_fpu_cp_req_bits_div,
  output  io_fpu_cp_req_bits_sqrt,
  output  io_fpu_cp_req_bits_round,
  output  io_fpu_cp_req_bits_wflags,
  output [2:0] io_fpu_cp_req_bits_rm,
  output [1:0] io_fpu_cp_req_bits_typ,
  output [64:0] io_fpu_cp_req_bits_in1,
  output [64:0] io_fpu_cp_req_bits_in2,
  output [64:0] io_fpu_cp_req_bits_in3,
  output  io_fpu_cp_resp_ready,
  input   io_fpu_cp_resp_valid,
  input  [64:0] io_fpu_cp_resp_bits_data,
  input  [4:0] io_fpu_cp_resp_bits_exc,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [6:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [6:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [10:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception
);
  reg  ex_ctrl_legal;
  reg [31:0] GEN_273;
  reg  ex_ctrl_fp;
  reg [31:0] GEN_274;
  reg  ex_ctrl_rocc;
  reg [31:0] GEN_275;
  reg  ex_ctrl_branch;
  reg [31:0] GEN_276;
  reg  ex_ctrl_jal;
  reg [31:0] GEN_277;
  reg  ex_ctrl_jalr;
  reg [31:0] GEN_278;
  reg  ex_ctrl_rxs2;
  reg [31:0] GEN_279;
  reg  ex_ctrl_rxs1;
  reg [31:0] GEN_280;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] GEN_281;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] GEN_282;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] GEN_283;
  reg  ex_ctrl_alu_dw;
  reg [31:0] GEN_284;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] GEN_285;
  reg  ex_ctrl_mem;
  reg [31:0] GEN_286;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] GEN_287;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] GEN_288;
  reg  ex_ctrl_rfs1;
  reg [31:0] GEN_289;
  reg  ex_ctrl_rfs2;
  reg [31:0] GEN_290;
  reg  ex_ctrl_rfs3;
  reg [31:0] GEN_291;
  reg  ex_ctrl_wfd;
  reg [31:0] GEN_292;
  reg  ex_ctrl_div;
  reg [31:0] GEN_293;
  reg  ex_ctrl_wxd;
  reg [31:0] GEN_294;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] GEN_295;
  reg  ex_ctrl_fence_i;
  reg [31:0] GEN_296;
  reg  ex_ctrl_fence;
  reg [31:0] GEN_297;
  reg  ex_ctrl_amo;
  reg [31:0] GEN_298;
  reg  mem_ctrl_legal;
  reg [31:0] GEN_299;
  reg  mem_ctrl_fp;
  reg [31:0] GEN_300;
  reg  mem_ctrl_rocc;
  reg [31:0] GEN_301;
  reg  mem_ctrl_branch;
  reg [31:0] GEN_302;
  reg  mem_ctrl_jal;
  reg [31:0] GEN_303;
  reg  mem_ctrl_jalr;
  reg [31:0] GEN_304;
  reg  mem_ctrl_rxs2;
  reg [31:0] GEN_305;
  reg  mem_ctrl_rxs1;
  reg [31:0] GEN_306;
  reg [1:0] mem_ctrl_sel_alu2;
  reg [31:0] GEN_307;
  reg [1:0] mem_ctrl_sel_alu1;
  reg [31:0] GEN_308;
  reg [2:0] mem_ctrl_sel_imm;
  reg [31:0] GEN_309;
  reg  mem_ctrl_alu_dw;
  reg [31:0] GEN_310;
  reg [3:0] mem_ctrl_alu_fn;
  reg [31:0] GEN_311;
  reg  mem_ctrl_mem;
  reg [31:0] GEN_312;
  reg [4:0] mem_ctrl_mem_cmd;
  reg [31:0] GEN_313;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] GEN_314;
  reg  mem_ctrl_rfs1;
  reg [31:0] GEN_315;
  reg  mem_ctrl_rfs2;
  reg [31:0] GEN_316;
  reg  mem_ctrl_rfs3;
  reg [31:0] GEN_317;
  reg  mem_ctrl_wfd;
  reg [31:0] GEN_318;
  reg  mem_ctrl_div;
  reg [31:0] GEN_319;
  reg  mem_ctrl_wxd;
  reg [31:0] GEN_320;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] GEN_321;
  reg  mem_ctrl_fence_i;
  reg [31:0] GEN_322;
  reg  mem_ctrl_fence;
  reg [31:0] GEN_323;
  reg  mem_ctrl_amo;
  reg [31:0] GEN_324;
  reg  wb_ctrl_legal;
  reg [31:0] GEN_325;
  reg  wb_ctrl_fp;
  reg [31:0] GEN_326;
  reg  wb_ctrl_rocc;
  reg [31:0] GEN_327;
  reg  wb_ctrl_branch;
  reg [31:0] GEN_328;
  reg  wb_ctrl_jal;
  reg [31:0] GEN_329;
  reg  wb_ctrl_jalr;
  reg [31:0] GEN_330;
  reg  wb_ctrl_rxs2;
  reg [31:0] GEN_331;
  reg  wb_ctrl_rxs1;
  reg [31:0] GEN_332;
  reg [1:0] wb_ctrl_sel_alu2;
  reg [31:0] GEN_333;
  reg [1:0] wb_ctrl_sel_alu1;
  reg [31:0] GEN_334;
  reg [2:0] wb_ctrl_sel_imm;
  reg [31:0] GEN_335;
  reg  wb_ctrl_alu_dw;
  reg [31:0] GEN_336;
  reg [3:0] wb_ctrl_alu_fn;
  reg [31:0] GEN_337;
  reg  wb_ctrl_mem;
  reg [31:0] GEN_338;
  reg [4:0] wb_ctrl_mem_cmd;
  reg [31:0] GEN_339;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] GEN_340;
  reg  wb_ctrl_rfs1;
  reg [31:0] GEN_341;
  reg  wb_ctrl_rfs2;
  reg [31:0] GEN_342;
  reg  wb_ctrl_rfs3;
  reg [31:0] GEN_343;
  reg  wb_ctrl_wfd;
  reg [31:0] GEN_344;
  reg  wb_ctrl_div;
  reg [31:0] GEN_345;
  reg  wb_ctrl_wxd;
  reg [31:0] GEN_346;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] GEN_347;
  reg  wb_ctrl_fence_i;
  reg [31:0] GEN_348;
  reg  wb_ctrl_fence;
  reg [31:0] GEN_349;
  reg  wb_ctrl_amo;
  reg [31:0] GEN_350;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] GEN_351;
  reg  ex_reg_valid;
  reg [31:0] GEN_352;
  reg  ex_reg_rvc;
  reg [31:0] GEN_353;
  reg  ex_reg_btb_hit;
  reg [31:0] GEN_354;
  reg  ex_reg_btb_resp_taken;
  reg [31:0] GEN_355;
  reg [1:0] ex_reg_btb_resp_mask;
  reg [31:0] GEN_356;
  reg  ex_reg_btb_resp_bridx;
  reg [31:0] GEN_357;
  reg [38:0] ex_reg_btb_resp_target;
  reg [63:0] GEN_358;
  reg [5:0] ex_reg_btb_resp_entry;
  reg [31:0] GEN_359;
  reg [6:0] ex_reg_btb_resp_bht_history;
  reg [31:0] GEN_360;
  reg [1:0] ex_reg_btb_resp_bht_value;
  reg [31:0] GEN_361;
  reg  ex_reg_xcpt;
  reg [31:0] GEN_362;
  reg  ex_reg_flush_pipe;
  reg [31:0] GEN_363;
  reg  ex_reg_load_use;
  reg [31:0] GEN_364;
  reg [63:0] ex_reg_cause;
  reg [63:0] GEN_365;
  reg  ex_reg_replay;
  reg [31:0] GEN_366;
  reg [39:0] ex_reg_pc;
  reg [63:0] GEN_367;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_368;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] GEN_369;
  reg  mem_reg_valid;
  reg [31:0] GEN_370;
  reg  mem_reg_rvc;
  reg [31:0] GEN_371;
  reg  mem_reg_btb_hit;
  reg [31:0] GEN_372;
  reg  mem_reg_btb_resp_taken;
  reg [31:0] GEN_373;
  reg [1:0] mem_reg_btb_resp_mask;
  reg [31:0] GEN_374;
  reg  mem_reg_btb_resp_bridx;
  reg [31:0] GEN_375;
  reg [38:0] mem_reg_btb_resp_target;
  reg [63:0] GEN_376;
  reg [5:0] mem_reg_btb_resp_entry;
  reg [31:0] GEN_377;
  reg [6:0] mem_reg_btb_resp_bht_history;
  reg [31:0] GEN_378;
  reg [1:0] mem_reg_btb_resp_bht_value;
  reg [31:0] GEN_379;
  reg  mem_reg_xcpt;
  reg [31:0] GEN_380;
  reg  mem_reg_replay;
  reg [31:0] GEN_381;
  reg  mem_reg_flush_pipe;
  reg [31:0] GEN_382;
  reg [63:0] mem_reg_cause;
  reg [63:0] GEN_383;
  reg  mem_reg_slow_bypass;
  reg [31:0] GEN_384;
  reg  mem_reg_load;
  reg [31:0] GEN_385;
  reg  mem_reg_store;
  reg [31:0] GEN_386;
  reg [39:0] mem_reg_pc;
  reg [63:0] GEN_387;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_388;
  reg [63:0] mem_reg_wdata;
  reg [63:0] GEN_389;
  reg [63:0] mem_reg_rs2;
  reg [63:0] GEN_390;
  wire  take_pc_mem;
  reg  wb_reg_valid;
  reg [31:0] GEN_391;
  reg  wb_reg_xcpt;
  reg [31:0] GEN_392;
  reg  wb_reg_replay;
  reg [31:0] GEN_393;
  reg [63:0] wb_reg_cause;
  reg [63:0] GEN_394;
  reg [39:0] wb_reg_pc;
  reg [63:0] GEN_395;
  reg [31:0] wb_reg_inst;
  reg [31:0] GEN_396;
  reg [63:0] wb_reg_wdata;
  reg [63:0] GEN_397;
  reg [63:0] wb_reg_rs2;
  reg [63:0] GEN_398;
  wire  take_pc_wb;
  wire  take_pc_mem_wb;
  wire  ibuf_clk;
  wire  ibuf_reset;
  wire  ibuf_io_imem_ready;
  wire  ibuf_io_imem_valid;
  wire  ibuf_io_imem_bits_btb_valid;
  wire  ibuf_io_imem_bits_btb_bits_taken;
  wire [1:0] ibuf_io_imem_bits_btb_bits_mask;
  wire  ibuf_io_imem_bits_btb_bits_bridx;
  wire [38:0] ibuf_io_imem_bits_btb_bits_target;
  wire [5:0] ibuf_io_imem_bits_btb_bits_entry;
  wire [6:0] ibuf_io_imem_bits_btb_bits_bht_history;
  wire [1:0] ibuf_io_imem_bits_btb_bits_bht_value;
  wire [39:0] ibuf_io_imem_bits_pc;
  wire [31:0] ibuf_io_imem_bits_data;
  wire [1:0] ibuf_io_imem_bits_mask;
  wire  ibuf_io_imem_bits_xcpt_if;
  wire  ibuf_io_imem_bits_replay;
  wire  ibuf_io_kill;
  wire [39:0] ibuf_io_pc;
  wire  ibuf_io_btb_resp_taken;
  wire [1:0] ibuf_io_btb_resp_mask;
  wire  ibuf_io_btb_resp_bridx;
  wire [38:0] ibuf_io_btb_resp_target;
  wire [5:0] ibuf_io_btb_resp_entry;
  wire [6:0] ibuf_io_btb_resp_bht_history;
  wire [1:0] ibuf_io_btb_resp_bht_value;
  wire  ibuf_io_inst_0_ready;
  wire  ibuf_io_inst_0_valid;
  wire  ibuf_io_inst_0_bits_pf0;
  wire  ibuf_io_inst_0_bits_pf1;
  wire  ibuf_io_inst_0_bits_replay;
  wire  ibuf_io_inst_0_bits_btb_hit;
  wire  ibuf_io_inst_0_bits_rvc;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3;
  wire  id_ctrl_legal;
  wire  id_ctrl_fp;
  wire  id_ctrl_rocc;
  wire  id_ctrl_branch;
  wire  id_ctrl_jal;
  wire  id_ctrl_jalr;
  wire  id_ctrl_rxs2;
  wire  id_ctrl_rxs1;
  wire [1:0] id_ctrl_sel_alu2;
  wire [1:0] id_ctrl_sel_alu1;
  wire [2:0] id_ctrl_sel_imm;
  wire  id_ctrl_alu_dw;
  wire [3:0] id_ctrl_alu_fn;
  wire  id_ctrl_mem;
  wire [4:0] id_ctrl_mem_cmd;
  wire [2:0] id_ctrl_mem_type;
  wire  id_ctrl_rfs1;
  wire  id_ctrl_rfs2;
  wire  id_ctrl_rfs3;
  wire  id_ctrl_wfd;
  wire  id_ctrl_div;
  wire  id_ctrl_wxd;
  wire [2:0] id_ctrl_csr;
  wire  id_ctrl_fence_i;
  wire  id_ctrl_fence;
  wire  id_ctrl_amo;
  wire [31:0] T_6645;
  wire  T_6647;
  wire [31:0] T_6649;
  wire  T_6651;
  wire [31:0] T_6653;
  wire  T_6655;
  wire [31:0] T_6657;
  wire  T_6659;
  wire [31:0] T_6661;
  wire  T_6663;
  wire [31:0] T_6665;
  wire  T_6667;
  wire [31:0] T_6669;
  wire  T_6671;
  wire [31:0] T_6673;
  wire  T_6675;
  wire [31:0] T_6677;
  wire  T_6679;
  wire [31:0] T_6681;
  wire  T_6683;
  wire [31:0] T_6685;
  wire  T_6687;
  wire [31:0] T_6689;
  wire  T_6691;
  wire [31:0] T_6693;
  wire  T_6695;
  wire [31:0] T_6697;
  wire  T_6699;
  wire [31:0] T_6701;
  wire  T_6703;
  wire  T_6707;
  wire [31:0] T_6709;
  wire  T_6711;
  wire  T_6715;
  wire [31:0] T_6717;
  wire  T_6719;
  wire [31:0] T_6721;
  wire  T_6723;
  wire  T_6727;
  wire [31:0] T_6729;
  wire  T_6731;
  wire [31:0] T_6733;
  wire  T_6735;
  wire [31:0] T_6737;
  wire  T_6739;
  wire [31:0] T_6741;
  wire  T_6743;
  wire [31:0] T_6745;
  wire  T_6747;
  wire  T_6749;
  wire [31:0] T_6751;
  wire  T_6753;
  wire [31:0] T_6755;
  wire  T_6757;
  wire [31:0] T_6759;
  wire  T_6761;
  wire [31:0] T_6763;
  wire  T_6765;
  wire  T_6769;
  wire [31:0] T_6771;
  wire  T_6773;
  wire  T_6775;
  wire [31:0] T_6777;
  wire  T_6779;
  wire [31:0] T_6781;
  wire  T_6783;
  wire [31:0] T_6785;
  wire  T_6787;
  wire [31:0] T_6789;
  wire  T_6791;
  wire [31:0] T_6793;
  wire  T_6795;
  wire [31:0] T_6797;
  wire  T_6799;
  wire [31:0] T_6801;
  wire  T_6803;
  wire  T_6806;
  wire  T_6807;
  wire  T_6808;
  wire  T_6809;
  wire  T_6810;
  wire  T_6811;
  wire  T_6812;
  wire  T_6813;
  wire  T_6814;
  wire  T_6815;
  wire  T_6816;
  wire  T_6817;
  wire  T_6818;
  wire  T_6819;
  wire  T_6820;
  wire  T_6821;
  wire  T_6822;
  wire  T_6823;
  wire  T_6824;
  wire  T_6825;
  wire  T_6826;
  wire  T_6827;
  wire  T_6828;
  wire  T_6829;
  wire  T_6830;
  wire  T_6831;
  wire  T_6832;
  wire  T_6833;
  wire  T_6834;
  wire  T_6835;
  wire  T_6836;
  wire  T_6837;
  wire  T_6838;
  wire  T_6839;
  wire  T_6840;
  wire  T_6841;
  wire  T_6842;
  wire  T_6843;
  wire  T_6844;
  wire  T_6845;
  wire [31:0] T_6847;
  wire  T_6849;
  wire [31:0] T_6851;
  wire  T_6853;
  wire  T_6856;
  wire [31:0] T_6859;
  wire  T_6861;
  wire [31:0] T_6865;
  wire  T_6867;
  wire [31:0] T_6871;
  wire  T_6873;
  wire [31:0] T_6877;
  wire  T_6879;
  wire [31:0] T_6881;
  wire  T_6883;
  wire [31:0] T_6885;
  wire  T_6887;
  wire  T_6890;
  wire  T_6891;
  wire [31:0] T_6893;
  wire  T_6895;
  wire [31:0] T_6897;
  wire  T_6899;
  wire [31:0] T_6901;
  wire  T_6903;
  wire [31:0] T_6905;
  wire  T_6907;
  wire [31:0] T_6909;
  wire  T_6911;
  wire  T_6914;
  wire  T_6915;
  wire  T_6916;
  wire  T_6917;
  wire [31:0] T_6919;
  wire  T_6921;
  wire [31:0] T_6923;
  wire  T_6925;
  wire [31:0] T_6927;
  wire  T_6929;
  wire [31:0] T_6931;
  wire  T_6933;
  wire [31:0] T_6935;
  wire  T_6937;
  wire  T_6940;
  wire  T_6941;
  wire  T_6942;
  wire  T_6943;
  wire  T_6947;
  wire [31:0] T_6949;
  wire  T_6951;
  wire [31:0] T_6953;
  wire  T_6955;
  wire  T_6958;
  wire  T_6959;
  wire  T_6960;
  wire [1:0] T_6961;
  wire [31:0] T_6963;
  wire  T_6965;
  wire [31:0] T_6967;
  wire  T_6969;
  wire [31:0] T_6971;
  wire  T_6973;
  wire  T_6976;
  wire  T_6977;
  wire  T_6978;
  wire  T_6979;
  wire  T_6983;
  wire  T_6986;
  wire [1:0] T_6987;
  wire  T_6991;
  wire  T_6995;
  wire  T_6998;
  wire [31:0] T_7000;
  wire  T_7002;
  wire  T_7005;
  wire [31:0] T_7007;
  wire  T_7009;
  wire [31:0] T_7011;
  wire  T_7013;
  wire  T_7017;
  wire  T_7020;
  wire  T_7021;
  wire [1:0] T_7022;
  wire [2:0] T_7023;
  wire [31:0] T_7025;
  wire  T_7027;
  wire [31:0] T_7029;
  wire  T_7031;
  wire  T_7034;
  wire [31:0] T_7036;
  wire  T_7038;
  wire [31:0] T_7040;
  wire  T_7042;
  wire [31:0] T_7044;
  wire  T_7046;
  wire  T_7049;
  wire  T_7050;
  wire [31:0] T_7052;
  wire  T_7054;
  wire [31:0] T_7056;
  wire  T_7058;
  wire  T_7062;
  wire [31:0] T_7064;
  wire  T_7066;
  wire [31:0] T_7068;
  wire  T_7070;
  wire [31:0] T_7072;
  wire  T_7074;
  wire  T_7077;
  wire  T_7078;
  wire  T_7079;
  wire  T_7080;
  wire  T_7081;
  wire [31:0] T_7083;
  wire  T_7085;
  wire [31:0] T_7087;
  wire  T_7089;
  wire [31:0] T_7091;
  wire  T_7093;
  wire [31:0] T_7095;
  wire  T_7097;
  wire  T_7100;
  wire  T_7101;
  wire  T_7102;
  wire  T_7106;
  wire [31:0] T_7108;
  wire  T_7110;
  wire  T_7113;
  wire  T_7114;
  wire  T_7115;
  wire [1:0] T_7116;
  wire [1:0] T_7117;
  wire [3:0] T_7118;
  wire [31:0] T_7120;
  wire  T_7122;
  wire [31:0] T_7124;
  wire  T_7126;
  wire [31:0] T_7128;
  wire  T_7130;
  wire  T_7133;
  wire  T_7134;
  wire  T_7135;
  wire  T_7136;
  wire  T_7137;
  wire  T_7138;
  wire  T_7139;
  wire [31:0] T_7141;
  wire  T_7143;
  wire [31:0] T_7145;
  wire  T_7147;
  wire [31:0] T_7149;
  wire  T_7151;
  wire [31:0] T_7153;
  wire  T_7155;
  wire  T_7158;
  wire  T_7159;
  wire  T_7160;
  wire [31:0] T_7162;
  wire  T_7164;
  wire [31:0] T_7166;
  wire  T_7168;
  wire  T_7171;
  wire [31:0] T_7173;
  wire  T_7175;
  wire [31:0] T_7177;
  wire  T_7179;
  wire [31:0] T_7181;
  wire  T_7183;
  wire  T_7186;
  wire  T_7187;
  wire  T_7188;
  wire [31:0] T_7190;
  wire  T_7192;
  wire [1:0] T_7196;
  wire [1:0] T_7197;
  wire [2:0] T_7198;
  wire [4:0] T_7199;
  wire [31:0] T_7201;
  wire  T_7203;
  wire [31:0] T_7207;
  wire  T_7209;
  wire [31:0] T_7213;
  wire  T_7215;
  wire [1:0] T_7218;
  wire [2:0] T_7219;
  wire [31:0] T_7221;
  wire  T_7223;
  wire [31:0] T_7225;
  wire  T_7227;
  wire [31:0] T_7229;
  wire  T_7231;
  wire  T_7234;
  wire  T_7235;
  wire [31:0] T_7237;
  wire  T_7239;
  wire [31:0] T_7241;
  wire  T_7243;
  wire [31:0] T_7245;
  wire  T_7247;
  wire  T_7250;
  wire  T_7251;
  wire  T_7252;
  wire [31:0] T_7256;
  wire  T_7258;
  wire  T_7262;
  wire  T_7265;
  wire  T_7266;
  wire  T_7267;
  wire [31:0] T_7269;
  wire  T_7271;
  wire  T_7277;
  wire  T_7281;
  wire [31:0] T_7283;
  wire  T_7285;
  wire  T_7289;
  wire [31:0] T_7291;
  wire  T_7293;
  wire [31:0] T_7295;
  wire  T_7297;
  wire [31:0] T_7299;
  wire  T_7301;
  wire  T_7304;
  wire  T_7305;
  wire  T_7306;
  wire  T_7307;
  wire  T_7308;
  wire  T_7309;
  wire [31:0] T_7311;
  wire  T_7313;
  wire [31:0] T_7317;
  wire  T_7319;
  wire [31:0] T_7323;
  wire  T_7325;
  wire [1:0] T_7328;
  wire [2:0] T_7329;
  wire [31:0] T_7331;
  wire  T_7333;
  wire  T_7339;
  wire [31:0] T_7343;
  wire  T_7345;
  wire  id_load_use;
  reg  id_reg_fence;
  reg [31:0] GEN_399;
  reg [63:0] T_7352 [0:30];
  reg [63:0] GEN_400;
  wire [63:0] T_7352_T_7361_data;
  wire [4:0] T_7352_T_7361_addr;
  wire  T_7352_T_7361_en;
  reg [63:0] GEN_401;
  wire [63:0] T_7352_T_7371_data;
  wire [4:0] T_7352_T_7371_addr;
  wire  T_7352_T_7371_en;
  reg [63:0] GEN_402;
  wire [63:0] T_7352_T_8104_data;
  wire [4:0] T_7352_T_8104_addr;
  wire  T_7352_T_8104_mask;
  wire  T_7352_T_8104_en;
  wire [63:0] id_rs_0;
  wire  T_7356;
  wire [4:0] T_7359;
  wire [4:0] T_7360;
  wire [63:0] T_7362;
  wire [63:0] id_rs_1;
  wire [4:0] T_7369;
  wire [4:0] T_7370;
  wire [63:0] T_7372;
  wire  ctrl_killd;
  wire  csr_clk;
  wire  csr_reset;
  wire  csr_io_prci_reset;
  wire  csr_io_prci_id;
  wire  csr_io_prci_interrupts_meip;
  wire  csr_io_prci_interrupts_seip;
  wire  csr_io_prci_interrupts_debug;
  wire  csr_io_prci_interrupts_mtip;
  wire  csr_io_prci_interrupts_msip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [63:0] csr_io_rw_rdata;
  wire [63:0] csr_io_rw_wdata;
  wire  csr_io_csr_stall;
  wire  csr_io_csr_xcpt;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [30:0] csr_io_status_zero3;
  wire  csr_io_status_sd_rv32;
  wire [1:0] csr_io_status_zero2;
  wire [4:0] csr_io_status_vm;
  wire [3:0] csr_io_status_zero1;
  wire  csr_io_status_mxr;
  wire  csr_io_status_pum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [6:0] csr_io_ptbr_asid;
  wire [37:0] csr_io_ptbr_ppn;
  wire [39:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire [63:0] csr_io_cause;
  wire [39:0] csr_io_pc;
  wire [39:0] csr_io_badaddr;
  wire  csr_io_fatc;
  wire [63:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_rocc_cmd_ready;
  wire  csr_io_rocc_cmd_valid;
  wire [6:0] csr_io_rocc_cmd_bits_inst_funct;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs1;
  wire  csr_io_rocc_cmd_bits_inst_xd;
  wire  csr_io_rocc_cmd_bits_inst_xs1;
  wire  csr_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rd;
  wire [6:0] csr_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] csr_io_rocc_cmd_bits_rs1;
  wire [63:0] csr_io_rocc_cmd_bits_rs2;
  wire  csr_io_rocc_cmd_bits_status_debug;
  wire [1:0] csr_io_rocc_cmd_bits_status_prv;
  wire  csr_io_rocc_cmd_bits_status_sd;
  wire [30:0] csr_io_rocc_cmd_bits_status_zero3;
  wire  csr_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] csr_io_rocc_cmd_bits_status_zero2;
  wire [4:0] csr_io_rocc_cmd_bits_status_vm;
  wire [3:0] csr_io_rocc_cmd_bits_status_zero1;
  wire  csr_io_rocc_cmd_bits_status_mxr;
  wire  csr_io_rocc_cmd_bits_status_pum;
  wire  csr_io_rocc_cmd_bits_status_mprv;
  wire [1:0] csr_io_rocc_cmd_bits_status_xs;
  wire [1:0] csr_io_rocc_cmd_bits_status_fs;
  wire [1:0] csr_io_rocc_cmd_bits_status_mpp;
  wire [1:0] csr_io_rocc_cmd_bits_status_hpp;
  wire  csr_io_rocc_cmd_bits_status_spp;
  wire  csr_io_rocc_cmd_bits_status_mpie;
  wire  csr_io_rocc_cmd_bits_status_hpie;
  wire  csr_io_rocc_cmd_bits_status_spie;
  wire  csr_io_rocc_cmd_bits_status_upie;
  wire  csr_io_rocc_cmd_bits_status_mie;
  wire  csr_io_rocc_cmd_bits_status_hie;
  wire  csr_io_rocc_cmd_bits_status_sie;
  wire  csr_io_rocc_cmd_bits_status_uie;
  wire  csr_io_rocc_resp_ready;
  wire  csr_io_rocc_resp_valid;
  wire [4:0] csr_io_rocc_resp_bits_rd;
  wire [63:0] csr_io_rocc_resp_bits_data;
  wire  csr_io_rocc_mem_req_ready;
  wire  csr_io_rocc_mem_req_valid;
  wire [39:0] csr_io_rocc_mem_req_bits_addr;
  wire [6:0] csr_io_rocc_mem_req_bits_tag;
  wire [4:0] csr_io_rocc_mem_req_bits_cmd;
  wire [2:0] csr_io_rocc_mem_req_bits_typ;
  wire  csr_io_rocc_mem_req_bits_phys;
  wire [63:0] csr_io_rocc_mem_req_bits_data;
  wire  csr_io_rocc_mem_s1_kill;
  wire [63:0] csr_io_rocc_mem_s1_data;
  wire  csr_io_rocc_mem_s2_nack;
  wire  csr_io_rocc_mem_resp_valid;
  wire [39:0] csr_io_rocc_mem_resp_bits_addr;
  wire [6:0] csr_io_rocc_mem_resp_bits_tag;
  wire [4:0] csr_io_rocc_mem_resp_bits_cmd;
  wire [2:0] csr_io_rocc_mem_resp_bits_typ;
  wire [63:0] csr_io_rocc_mem_resp_bits_data;
  wire  csr_io_rocc_mem_resp_bits_replay;
  wire  csr_io_rocc_mem_resp_bits_has_data;
  wire [63:0] csr_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] csr_io_rocc_mem_resp_bits_store_data;
  wire  csr_io_rocc_mem_replay_next;
  wire  csr_io_rocc_mem_xcpt_ma_ld;
  wire  csr_io_rocc_mem_xcpt_ma_st;
  wire  csr_io_rocc_mem_xcpt_pf_ld;
  wire  csr_io_rocc_mem_xcpt_pf_st;
  wire  csr_io_rocc_mem_invalidate_lr;
  wire  csr_io_rocc_mem_ordered;
  wire  csr_io_rocc_busy;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_rocc_autl_acquire_ready;
  wire  csr_io_rocc_autl_acquire_valid;
  wire [25:0] csr_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] csr_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_acquire_bits_addr_beat;
  wire  csr_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] csr_io_rocc_autl_acquire_bits_a_type;
  wire [10:0] csr_io_rocc_autl_acquire_bits_union;
  wire [63:0] csr_io_rocc_autl_acquire_bits_data;
  wire  csr_io_rocc_autl_grant_ready;
  wire  csr_io_rocc_autl_grant_valid;
  wire [2:0] csr_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] csr_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_grant_bits_manager_xact_id;
  wire  csr_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] csr_io_rocc_autl_grant_bits_g_type;
  wire [63:0] csr_io_rocc_autl_grant_bits_data;
  wire  csr_io_rocc_fpu_req_ready;
  wire  csr_io_rocc_fpu_req_valid;
  wire [4:0] csr_io_rocc_fpu_req_bits_cmd;
  wire  csr_io_rocc_fpu_req_bits_ldst;
  wire  csr_io_rocc_fpu_req_bits_wen;
  wire  csr_io_rocc_fpu_req_bits_ren1;
  wire  csr_io_rocc_fpu_req_bits_ren2;
  wire  csr_io_rocc_fpu_req_bits_ren3;
  wire  csr_io_rocc_fpu_req_bits_swap12;
  wire  csr_io_rocc_fpu_req_bits_swap23;
  wire  csr_io_rocc_fpu_req_bits_single;
  wire  csr_io_rocc_fpu_req_bits_fromint;
  wire  csr_io_rocc_fpu_req_bits_toint;
  wire  csr_io_rocc_fpu_req_bits_fastpipe;
  wire  csr_io_rocc_fpu_req_bits_fma;
  wire  csr_io_rocc_fpu_req_bits_div;
  wire  csr_io_rocc_fpu_req_bits_sqrt;
  wire  csr_io_rocc_fpu_req_bits_round;
  wire  csr_io_rocc_fpu_req_bits_wflags;
  wire [2:0] csr_io_rocc_fpu_req_bits_rm;
  wire [1:0] csr_io_rocc_fpu_req_bits_typ;
  wire [64:0] csr_io_rocc_fpu_req_bits_in1;
  wire [64:0] csr_io_rocc_fpu_req_bits_in2;
  wire [64:0] csr_io_rocc_fpu_req_bits_in3;
  wire  csr_io_rocc_fpu_resp_ready;
  wire  csr_io_rocc_fpu_resp_valid;
  wire [64:0] csr_io_rocc_fpu_resp_bits_data;
  wire [4:0] csr_io_rocc_fpu_resp_bits_exc;
  wire  csr_io_rocc_exception;
  wire  csr_io_interrupt;
  wire [63:0] csr_io_interrupt_cause;
  wire [3:0] csr_io_bp_0_control_ttype;
  wire  csr_io_bp_0_control_dmode;
  wire [5:0] csr_io_bp_0_control_maskmax;
  wire [39:0] csr_io_bp_0_control_reserved;
  wire  csr_io_bp_0_control_action;
  wire  csr_io_bp_0_control_chain;
  wire [1:0] csr_io_bp_0_control_zero;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_x;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_r;
  wire [38:0] csr_io_bp_0_address;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  T_7374;
  wire  T_7375;
  wire  T_7376;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire [11:0] id_csr_addr;
  wire  T_7380;
  wire  T_7381;
  wire [11:0] T_7511;
  wire  T_7513;
  wire [11:0] T_7515;
  wire  T_7517;
  wire  T_7520;
  wire  T_7523;
  wire  T_7524;
  wire  id_csr_flush;
  wire  T_7526;
  wire  T_7528;
  wire  T_7530;
  wire  T_7531;
  wire  T_7532;
  wire  T_7534;
  wire  T_7536;
  wire  T_7537;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  T_7538;
  wire  id_fence_next;
  wire  T_7540;
  wire  id_mem_busy;
  wire  T_7546;
  wire  T_7548;
  wire  T_7549;
  wire  T_7551;
  wire  T_7552;
  wire  T_7553;
  wire  T_7554;
  wire  T_7555;
  wire  T_7556;
  wire  T_7557;
  wire  bpu_clk;
  wire  bpu_reset;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_status_sd;
  wire [30:0] bpu_io_status_zero3;
  wire  bpu_io_status_sd_rv32;
  wire [1:0] bpu_io_status_zero2;
  wire [4:0] bpu_io_status_vm;
  wire [3:0] bpu_io_status_zero1;
  wire  bpu_io_status_mxr;
  wire  bpu_io_status_pum;
  wire  bpu_io_status_mprv;
  wire [1:0] bpu_io_status_xs;
  wire [1:0] bpu_io_status_fs;
  wire [1:0] bpu_io_status_mpp;
  wire [1:0] bpu_io_status_hpp;
  wire  bpu_io_status_spp;
  wire  bpu_io_status_mpie;
  wire  bpu_io_status_hpie;
  wire  bpu_io_status_spie;
  wire  bpu_io_status_upie;
  wire  bpu_io_status_mie;
  wire  bpu_io_status_hie;
  wire  bpu_io_status_sie;
  wire  bpu_io_status_uie;
  wire [3:0] bpu_io_bp_0_control_ttype;
  wire  bpu_io_bp_0_control_dmode;
  wire [5:0] bpu_io_bp_0_control_maskmax;
  wire [39:0] bpu_io_bp_0_control_reserved;
  wire  bpu_io_bp_0_control_action;
  wire  bpu_io_bp_0_control_chain;
  wire [1:0] bpu_io_bp_0_control_zero;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_x;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_r;
  wire [38:0] bpu_io_bp_0_address;
  wire [38:0] bpu_io_pc;
  wire [38:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  bpu_io_debug_if;
  wire  bpu_io_debug_ld;
  wire  bpu_io_debug_st;
  wire  id_xcpt_if;
  wire  T_7562;
  wire  T_7563;
  wire  T_7564;
  wire  id_xcpt;
  wire [1:0] T_7565;
  wire [1:0] T_7566;
  wire [3:0] T_7567;
  wire [63:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  T_7571;
  wire  T_7572;
  wire  T_7574;
  wire  T_7575;
  wire  T_7577;
  wire  T_7578;
  wire  id_bypass_src_0_1;
  wire  T_7579;
  wire  id_bypass_src_0_2;
  wire  id_bypass_src_0_3;
  wire  T_7581;
  wire  T_7582;
  wire  id_bypass_src_1_1;
  wire  T_7583;
  wire  id_bypass_src_1_2;
  wire  id_bypass_src_1_3;
  wire [63:0] bypass_mux_0;
  wire [63:0] bypass_mux_1;
  wire [63:0] bypass_mux_2;
  wire [63:0] bypass_mux_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] GEN_403;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] GEN_404;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] GEN_405;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] GEN_406;
  reg [61:0] ex_reg_rs_msb_0;
  reg [63:0] GEN_407;
  reg [61:0] ex_reg_rs_msb_1;
  reg [63:0] GEN_408;
  wire [63:0] T_7612;
  wire [63:0] GEN_0;
  wire [63:0] GEN_2;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] ex_rs_0;
  wire [63:0] T_7613;
  wire [63:0] GEN_1;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] ex_rs_1;
  wire  T_7614;
  wire  T_7616;
  wire  T_7617;
  wire  T_7618;
  wire  T_7619;
  wire [10:0] T_7620;
  wire [10:0] T_7621;
  wire [10:0] T_7622;
  wire  T_7623;
  wire  T_7624;
  wire  T_7625;
  wire [7:0] T_7626;
  wire [7:0] T_7627;
  wire [7:0] T_7628;
  wire  T_7631;
  wire  T_7633;
  wire  T_7634;
  wire  T_7635;
  wire  T_7636;
  wire  T_7637;
  wire  T_7638;
  wire  T_7639;
  wire  T_7640;
  wire  T_7641;
  wire [5:0] T_7646;
  wire [5:0] T_7647;
  wire  T_7650;
  wire  T_7652;
  wire [3:0] T_7653;
  wire [3:0] T_7655;
  wire [3:0] T_7656;
  wire [3:0] T_7657;
  wire [3:0] T_7658;
  wire [3:0] T_7659;
  wire  T_7662;
  wire  T_7665;
  wire  T_7668;
  wire  T_7670;
  wire  T_7672;
  wire [9:0] T_7673;
  wire [10:0] T_7674;
  wire  T_7675;
  wire [7:0] T_7676;
  wire [8:0] T_7677;
  wire [10:0] T_7678;
  wire  T_7679;
  wire [11:0] T_7680;
  wire [20:0] T_7681;
  wire [31:0] T_7682;
  wire [31:0] ex_imm;
  wire [63:0] T_7684;
  wire [39:0] T_7685;
  wire  T_7686;
  wire [39:0] T_7687;
  wire  T_7688;
  wire [63:0] ex_op1;
  wire [63:0] T_7690;
  wire [3:0] T_7693;
  wire  T_7694;
  wire [3:0] T_7695;
  wire  T_7696;
  wire [31:0] T_7697;
  wire  T_7698;
  wire [63:0] ex_op2;
  wire  alu_clk;
  wire  alu_reset;
  wire  alu_io_dw;
  wire [3:0] alu_io_fn;
  wire [63:0] alu_io_in2;
  wire [63:0] alu_io_in1;
  wire [63:0] alu_io_out;
  wire [63:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [63:0] T_7699;
  wire [63:0] T_7700;
  wire  div_clk;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire  div_io_req_bits_dw;
  wire [63:0] div_io_req_bits_in1;
  wire [63:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [63:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  T_7701;
  wire  T_7703;
  wire  T_7705;
  wire  T_7706;
  wire  T_7707;
  wire  T_7710;
  wire  T_7714;
  wire [63:0] GEN_8;
  wire  GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire [5:0] GEN_13;
  wire [6:0] GEN_14;
  wire [1:0] GEN_15;
  wire  T_7718;
  wire  T_7720;
  wire  T_7721;
  wire  T_7722;
  wire [1:0] GEN_16;
  wire  GEN_17;
  wire [3:0] GEN_18;
  wire  GEN_19;
  wire [1:0] GEN_20;
  wire [1:0] GEN_21;
  wire  GEN_22;
  wire  T_7724;
  wire  T_7725;
  wire  T_7726;
  wire  GEN_23;
  wire  GEN_24;
  wire  T_7729;
  wire  T_7730;
  wire  T_7731;
  wire [1:0] T_7736;
  wire [1:0] T_7737;
  wire [1:0] T_7738;
  wire  T_7740;
  wire  T_7741;
  wire [1:0] T_7742;
  wire [61:0] T_7743;
  wire [1:0] GEN_25;
  wire [61:0] GEN_26;
  wire  T_7744;
  wire  T_7745;
  wire  T_7746;
  wire [1:0] T_7751;
  wire [1:0] T_7752;
  wire [1:0] T_7753;
  wire  T_7755;
  wire  T_7756;
  wire [1:0] T_7757;
  wire [61:0] T_7758;
  wire [1:0] GEN_27;
  wire [61:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [1:0] GEN_37;
  wire [1:0] GEN_38;
  wire [2:0] GEN_39;
  wire  GEN_40;
  wire [3:0] GEN_41;
  wire  GEN_42;
  wire [4:0] GEN_43;
  wire [2:0] GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire [2:0] GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [61:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [61:0] GEN_63;
  wire  T_7761;
  wire  T_7762;
  wire [31:0] GEN_64;
  wire [39:0] GEN_65;
  wire  T_7763;
  wire  ex_pc_valid;
  wire  T_7765;
  wire  wb_dcache_miss;
  wire  T_7767;
  wire  T_7768;
  wire  T_7770;
  wire  T_7771;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  T_7772;
  wire  T_7773;
  wire  replay_ex;
  wire  T_7774;
  wire  T_7776;
  wire  ctrl_killx;
  wire  T_7777;
  wire [2:0] T_7783_0;
  wire [2:0] T_7783_1;
  wire [2:0] T_7783_2;
  wire [2:0] T_7783_3;
  wire  T_7785;
  wire  T_7786;
  wire  T_7787;
  wire  T_7788;
  wire  T_7791;
  wire  T_7792;
  wire  T_7793;
  wire  ex_slow_bypass;
  wire  T_7794;
  wire  T_7795;
  wire  ex_xcpt;
  wire [63:0] ex_cause;
  wire  mem_br_taken;
  wire [39:0] T_7797;
  wire  T_7798;
  wire  T_7801;
  wire  T_7802;
  wire [10:0] T_7807;
  wire [7:0] T_7811;
  wire [7:0] T_7812;
  wire [7:0] T_7813;
  wire  T_7819;
  wire  T_7820;
  wire  T_7822;
  wire  T_7823;
  wire [5:0] T_7831;
  wire [3:0] T_7838;
  wire [3:0] T_7841;
  wire [9:0] T_7858;
  wire [10:0] T_7859;
  wire  T_7860;
  wire [7:0] T_7861;
  wire [8:0] T_7862;
  wire [10:0] T_7863;
  wire  T_7864;
  wire [11:0] T_7865;
  wire [20:0] T_7866;
  wire [31:0] T_7867;
  wire [31:0] T_7868;
  wire [9:0] T_7928;
  wire [10:0] T_7929;
  wire  T_7930;
  wire [7:0] T_7931;
  wire [8:0] T_7932;
  wire [20:0] T_7936;
  wire [31:0] T_7937;
  wire [31:0] T_7938;
  wire [3:0] T_7941;
  wire [31:0] T_7942;
  wire [31:0] T_7943;
  wire [39:0] GEN_174;
  wire [40:0] T_7944;
  wire [39:0] T_7945;
  wire [39:0] mem_br_target;
  wire [25:0] T_7946;
  wire [1:0] T_7947;
  wire [1:0] T_7948;
  wire  T_7950;
  wire  T_7952;
  wire  T_7953;
  wire  T_7955;
  wire [25:0] T_7956;
  wire  T_7958;
  wire  T_7961;
  wire  T_7962;
  wire  T_7964;
  wire  T_7965;
  wire  T_7966;
  wire  T_7967;
  wire [38:0] T_7968;
  wire [39:0] T_7969;
  wire [39:0] T_7970;
  wire [39:0] T_7971;
  wire [39:0] T_7973;
  wire [39:0] T_7974;
  wire [39:0] mem_npc;
  wire  T_7975;
  wire  T_7976;
  wire  T_7978;
  wire  mem_wrong_npc;
  wire  T_7980;
  wire  T_7982;
  wire [63:0] T_7983;
  wire [63:0] T_7984;
  wire [63:0] mem_int_wdata;
  wire  T_7985;
  wire  mem_cfi;
  wire  T_7987;
  wire  mem_cfi_taken;
  wire  T_7988;
  wire  T_7989;
  wire  T_7991;
  wire  T_7994;
  wire  T_7997;
  wire  T_8000;
  wire [63:0] GEN_66;
  wire  T_8001;
  wire  T_8002;
  wire  T_8003;
  wire  T_8005;
  wire  T_8006;
  wire  T_8007;
  wire  T_8008;
  wire  T_8009;
  wire  T_8010;
  wire  T_8011;
  wire  T_8013;
  wire  T_8017;
  wire  T_8018;
  wire  GEN_67;
  wire [1:0] GEN_68;
  wire  GEN_69;
  wire [38:0] GEN_70;
  wire [5:0] GEN_71;
  wire [6:0] GEN_72;
  wire [1:0] GEN_73;
  wire  T_8019;
  wire  T_8020;
  wire [63:0] GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire [1:0] GEN_83;
  wire [1:0] GEN_84;
  wire [2:0] GEN_85;
  wire  GEN_86;
  wire [3:0] GEN_87;
  wire  GEN_88;
  wire [4:0] GEN_89;
  wire [2:0] GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire [1:0] GEN_106;
  wire  GEN_107;
  wire [38:0] GEN_108;
  wire [5:0] GEN_109;
  wire [6:0] GEN_110;
  wire [1:0] GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire [31:0] GEN_114;
  wire [39:0] GEN_115;
  wire [63:0] GEN_116;
  wire [63:0] GEN_117;
  wire  T_8021;
  wire  T_8022;
  wire  mem_breakpoint;
  wire  T_8023;
  wire  T_8024;
  wire  mem_debug_breakpoint;
  wire  T_8028;
  wire  T_8030;
  wire  T_8032;
  wire  T_8034;
  wire  T_8036;
  wire  T_8038;
  wire  T_8039;
  wire  T_8040;
  wire  mem_new_xcpt;
  wire [2:0] T_8041;
  wire [2:0] T_8042;
  wire [2:0] T_8043;
  wire [2:0] T_8045;
  wire [3:0] mem_new_cause;
  wire  T_8046;
  wire  T_8047;
  wire  mem_xcpt;
  wire [63:0] mem_cause;
  wire  dcache_kill_mem;
  wire  T_8049;
  wire  fpu_kill_mem;
  wire  T_8050;
  wire  replay_mem;
  wire  T_8051;
  wire  T_8052;
  wire  T_8054;
  wire  killm_common;
  wire  T_8055;
  reg  T_8056;
  reg [31:0] GEN_409;
  wire  T_8057;
  wire  T_8058;
  wire  ctrl_killm;
  wire  T_8060;
  wire  T_8062;
  wire  T_8063;
  wire  T_8066;
  wire [63:0] GEN_118;
  wire  T_8067;
  wire  T_8068;
  wire  T_8071;
  wire  T_8072;
  wire [63:0] T_8073;
  wire [63:0] GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire [1:0] GEN_128;
  wire [1:0] GEN_129;
  wire [2:0] GEN_130;
  wire  GEN_131;
  wire [3:0] GEN_132;
  wire  GEN_133;
  wire [4:0] GEN_134;
  wire [2:0] GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire [2:0] GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire [63:0] GEN_146;
  wire [63:0] GEN_147;
  wire [31:0] GEN_148;
  wire [39:0] GEN_149;
  wire  T_8074;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  T_8077;
  wire  replay_wb_rocc;
  wire  replay_wb;
  wire  wb_xcpt;
  wire  T_8078;
  wire  T_8079;
  wire  T_8080;
  wire  dmem_resp_xpu;
  wire [4:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  T_8084;
  wire  T_8086;
  wire [63:0] ll_wdata;
  wire [4:0] ll_waddr;
  wire  T_8087;
  wire  ll_wen;
  wire  T_8088;
  wire  GEN_150;
  wire [4:0] GEN_151;
  wire  GEN_152;
  wire  T_8092;
  wire  T_8093;
  wire  T_8095;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [4:0] rf_waddr;
  wire  T_8096;
  wire  T_8097;
  wire [63:0] T_8098;
  wire [63:0] T_8099;
  wire [63:0] rf_wdata;
  wire  T_8101;
  wire [4:0] T_8103;
  wire  T_8105;
  wire [63:0] GEN_153;
  wire  T_8106;
  wire [63:0] GEN_154;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire  GEN_164;
  wire [63:0] GEN_167;
  wire [63:0] GEN_168;
  wire [25:0] T_8107;
  wire [1:0] T_8108;
  wire [1:0] T_8109;
  wire  T_8111;
  wire  T_8113;
  wire  T_8114;
  wire  T_8116;
  wire [25:0] T_8117;
  wire  T_8119;
  wire  T_8122;
  wire  T_8123;
  wire  T_8125;
  wire  T_8126;
  wire  T_8127;
  wire  T_8128;
  wire [38:0] T_8129;
  wire [39:0] T_8130;
  wire [11:0] T_8131;
  wire [2:0] T_8132;
  wire  T_8134;
  wire  T_8135;
  wire  T_8137;
  wire  T_8138;
  wire  T_8140;
  wire  T_8141;
  reg [31:0] T_8143;
  reg [31:0] GEN_410;
  wire [30:0] T_8144;
  wire [31:0] GEN_175;
  wire [31:0] T_8145;
  wire [31:0] T_8148;
  wire [31:0] T_8150;
  wire [31:0] T_8151;
  wire [31:0] T_8152;
  wire [31:0] GEN_169;
  wire [31:0] T_8154;
  wire  T_8155;
  wire  T_8156;
  wire [31:0] T_8157;
  wire  T_8158;
  wire  T_8159;
  wire [31:0] T_8160;
  wire  T_8161;
  wire  T_8162;
  wire  T_8163;
  wire  id_sboard_hazard;
  wire  T_8164;
  wire [31:0] T_8166;
  wire [31:0] T_8168;
  wire [31:0] T_8169;
  wire  T_8170;
  wire [31:0] GEN_170;
  wire  T_8171;
  wire  T_8172;
  wire  T_8173;
  wire  T_8174;
  wire  T_8175;
  wire  ex_cannot_bypass;
  wire  T_8176;
  wire  T_8177;
  wire  T_8178;
  wire  T_8179;
  wire  T_8180;
  wire  T_8181;
  wire  T_8182;
  wire  T_8183;
  wire  data_hazard_ex;
  wire  T_8185;
  wire  T_8187;
  wire  T_8188;
  wire  T_8189;
  wire  T_8191;
  wire  T_8192;
  wire  T_8193;
  wire  T_8194;
  wire  fp_data_hazard_ex;
  wire  T_8195;
  wire  T_8196;
  wire  id_ex_hazard;
  wire  T_8198;
  wire  T_8199;
  wire  T_8200;
  wire  T_8201;
  wire  T_8202;
  wire  mem_cannot_bypass;
  wire  T_8203;
  wire  T_8204;
  wire  T_8205;
  wire  T_8206;
  wire  T_8207;
  wire  T_8208;
  wire  T_8209;
  wire  T_8210;
  wire  data_hazard_mem;
  wire  T_8212;
  wire  T_8214;
  wire  T_8215;
  wire  T_8216;
  wire  T_8218;
  wire  T_8219;
  wire  T_8220;
  wire  T_8221;
  wire  fp_data_hazard_mem;
  wire  T_8222;
  wire  T_8223;
  wire  id_mem_hazard;
  wire  T_8224;
  wire  T_8225;
  wire  T_8226;
  wire  T_8227;
  wire  T_8228;
  wire  T_8229;
  wire  T_8230;
  wire  T_8231;
  wire  T_8232;
  wire  T_8233;
  wire  data_hazard_wb;
  wire  T_8235;
  wire  T_8237;
  wire  T_8238;
  wire  T_8239;
  wire  T_8241;
  wire  T_8242;
  wire  T_8243;
  wire  T_8244;
  wire  fp_data_hazard_wb;
  wire  T_8245;
  wire  T_8246;
  wire  id_wb_hazard;
  reg [31:0] T_8248;
  reg [31:0] GEN_411;
  wire  T_8250;
  wire  T_8251;
  wire  T_8252;
  wire [31:0] T_8256;
  wire [31:0] T_8257;
  wire [31:0] GEN_171;
  wire  T_8259;
  wire [31:0] T_8261;
  wire [31:0] T_8263;
  wire [31:0] T_8264;
  wire [31:0] T_8265;
  wire  T_8266;
  wire [31:0] GEN_172;
  wire [31:0] T_8268;
  wire [31:0] T_8270;
  wire [31:0] T_8271;
  wire [31:0] T_8272;
  wire  T_8273;
  wire [31:0] GEN_173;
  wire  T_8275;
  wire  T_8276;
  wire [31:0] T_8277;
  wire  T_8278;
  wire  T_8279;
  wire [31:0] T_8280;
  wire  T_8281;
  wire  T_8282;
  wire [31:0] T_8283;
  wire  T_8284;
  wire  T_8285;
  wire [31:0] T_8286;
  wire  T_8287;
  wire  T_8288;
  wire  T_8289;
  wire  T_8290;
  wire  T_8291;
  wire  id_stall_fpu;
  reg  dcache_blocked;
  reg [31:0] GEN_412;
  wire  T_8295;
  wire  T_8296;
  reg  rocc_blocked;
  reg [31:0] GEN_413;
  wire  T_8299;
  wire  T_8302;
  wire  T_8303;
  wire  T_8304;
  wire  T_8305;
  wire  T_8306;
  wire  T_8307;
  wire  T_8308;
  wire  T_8309;
  wire  T_8310;
  wire  T_8311;
  wire  T_8312;
  wire  T_8313;
  wire  T_8314;
  wire  ctrl_stalld;
  wire  T_8316;
  wire  T_8317;
  wire  T_8318;
  wire  T_8319;
  wire  T_8320;
  wire  T_8323;
  wire [39:0] T_8324;
  wire [39:0] T_8325;
  wire  T_8326;
  wire  T_8328;
  wire  T_8329;
  wire  T_8331;
  wire  T_8332;
  wire  T_8333;
  wire  T_8336;
  wire  T_8338;
  wire  T_8339;
  wire  T_8340;
  wire  T_8341;
  wire  T_8342;
  wire  T_8344;
  wire  T_8345;
  wire  T_8346;
  wire [4:0] T_8347;
  wire [4:0] T_8350;
  wire  T_8351;
  wire  T_8352;
  wire [1:0] T_8355;
  wire [39:0] GEN_176;
  wire [40:0] T_8356;
  wire [39:0] T_8357;
  wire [38:0] T_8358;
  wire [38:0] T_8360;
  wire [38:0] T_8361;
  wire  T_8365;
  wire  T_8369;
  wire  T_8370;
  wire  T_8373;
  wire  T_8374;
  wire  T_8375;
  wire [5:0] ex_dcache_tag;
  wire [25:0] T_8377;
  wire [1:0] T_8378;
  wire [1:0] T_8379;
  wire  T_8381;
  wire  T_8383;
  wire  T_8384;
  wire  T_8386;
  wire [25:0] T_8387;
  wire  T_8389;
  wire  T_8392;
  wire  T_8393;
  wire  T_8395;
  wire  T_8396;
  wire  T_8397;
  wire  T_8398;
  wire [38:0] T_8399;
  wire [39:0] T_8400;
  wire [63:0] T_8401;
  wire  T_8402;
  wire  T_8404;
  wire  T_8405;
  wire [1:0] T_8406;
  wire [1:0] T_8407;
  wire [3:0] T_8408;
  wire  T_8410;
  wire  T_8411;
  wire  T_8413;
  wire  T_8416;
  wire  T_8417;
  wire  T_8420;
  wire [6:0] T_8439_funct;
  wire [4:0] T_8439_rs2;
  wire [4:0] T_8439_rs1;
  wire  T_8439_xd;
  wire  T_8439_xs1;
  wire  T_8439_xs2;
  wire [4:0] T_8439_rd;
  wire [6:0] T_8439_opcode;
  wire [31:0] T_8449;
  wire [6:0] T_8450;
  wire [4:0] T_8451;
  wire  T_8452;
  wire  T_8453;
  wire  T_8454;
  wire [4:0] T_8455;
  wire [4:0] T_8456;
  wire [6:0] T_8457;
  wire [31:0] T_8458;
  wire [4:0] T_8460;
  wire [4:0] T_8461;
  reg [63:0] T_8462;
  reg [63:0] GEN_414;
  reg [63:0] T_8463;
  reg [63:0] GEN_415;
  wire [4:0] T_8464;
  reg [63:0] T_8465;
  reg [63:0] GEN_416;
  reg [63:0] T_8466;
  reg [63:0] GEN_417;
  wire  T_8468;
  wire  GEN_155;
  reg [31:0] GEN_418;
  wire [63:0] GEN_156;
  reg [63:0] GEN_419;
  wire  GEN_157;
  reg [31:0] GEN_420;
  wire [4:0] GEN_158;
  reg [31:0] GEN_421;
  wire  GEN_159;
  reg [31:0] GEN_422;
  wire  GEN_162;
  reg [31:0] GEN_423;
  wire  GEN_163;
  reg [31:0] GEN_424;
  wire  GEN_165;
  reg [31:0] GEN_425;
  wire  GEN_166;
  reg [31:0] GEN_426;
  wire  GEN_177;
  reg [31:0] GEN_427;
  wire  GEN_178;
  reg [31:0] GEN_428;
  wire  GEN_179;
  reg [31:0] GEN_429;
  wire  GEN_180;
  reg [31:0] GEN_430;
  wire  GEN_181;
  reg [31:0] GEN_431;
  wire  GEN_182;
  reg [31:0] GEN_432;
  wire  GEN_183;
  reg [31:0] GEN_433;
  wire  GEN_184;
  reg [31:0] GEN_434;
  wire  GEN_185;
  reg [31:0] GEN_435;
  wire  GEN_186;
  reg [31:0] GEN_436;
  wire  GEN_187;
  reg [31:0] GEN_437;
  wire [2:0] GEN_188;
  reg [31:0] GEN_438;
  wire [1:0] GEN_189;
  reg [31:0] GEN_439;
  wire [64:0] GEN_190;
  reg [95:0] GEN_440;
  wire [64:0] GEN_191;
  reg [95:0] GEN_441;
  wire [64:0] GEN_192;
  reg [95:0] GEN_442;
  wire  GEN_193;
  reg [31:0] GEN_443;
  wire  GEN_194;
  reg [31:0] GEN_444;
  wire  GEN_195;
  reg [31:0] GEN_445;
  wire  GEN_196;
  reg [31:0] GEN_446;
  wire  GEN_197;
  reg [31:0] GEN_447;
  wire [39:0] GEN_198;
  reg [63:0] GEN_448;
  wire [6:0] GEN_199;
  reg [31:0] GEN_449;
  wire [4:0] GEN_200;
  reg [31:0] GEN_450;
  wire [2:0] GEN_201;
  reg [31:0] GEN_451;
  wire [63:0] GEN_202;
  reg [63:0] GEN_452;
  wire  GEN_203;
  reg [31:0] GEN_453;
  wire  GEN_204;
  reg [31:0] GEN_454;
  wire [63:0] GEN_205;
  reg [63:0] GEN_455;
  wire [63:0] GEN_206;
  reg [63:0] GEN_456;
  wire  GEN_207;
  reg [31:0] GEN_457;
  wire  GEN_208;
  reg [31:0] GEN_458;
  wire  GEN_209;
  reg [31:0] GEN_459;
  wire  GEN_210;
  reg [31:0] GEN_460;
  wire  GEN_211;
  reg [31:0] GEN_461;
  wire  GEN_212;
  reg [31:0] GEN_462;
  wire  GEN_213;
  reg [31:0] GEN_463;
  wire  GEN_214;
  reg [31:0] GEN_464;
  wire [2:0] GEN_215;
  reg [31:0] GEN_465;
  wire [1:0] GEN_216;
  reg [31:0] GEN_466;
  wire [2:0] GEN_217;
  reg [31:0] GEN_467;
  wire  GEN_218;
  reg [31:0] GEN_468;
  wire [3:0] GEN_219;
  reg [31:0] GEN_469;
  wire [63:0] GEN_220;
  reg [63:0] GEN_470;
  wire  GEN_221;
  reg [31:0] GEN_471;
  wire  GEN_222;
  reg [31:0] GEN_472;
  wire [64:0] GEN_223;
  reg [95:0] GEN_473;
  wire [4:0] GEN_224;
  reg [31:0] GEN_474;
  wire  GEN_225;
  reg [31:0] GEN_475;
  wire  GEN_226;
  reg [31:0] GEN_476;
  wire [4:0] GEN_227;
  reg [31:0] GEN_477;
  wire [63:0] GEN_228;
  reg [63:0] GEN_478;
  wire  GEN_229;
  reg [31:0] GEN_479;
  wire [39:0] GEN_230;
  reg [63:0] GEN_480;
  wire [6:0] GEN_231;
  reg [31:0] GEN_481;
  wire [4:0] GEN_232;
  reg [31:0] GEN_482;
  wire [2:0] GEN_233;
  reg [31:0] GEN_483;
  wire  GEN_234;
  reg [31:0] GEN_484;
  wire [63:0] GEN_235;
  reg [63:0] GEN_485;
  wire  GEN_236;
  reg [31:0] GEN_486;
  wire [63:0] GEN_237;
  reg [63:0] GEN_487;
  wire  GEN_238;
  reg [31:0] GEN_488;
  wire  GEN_239;
  reg [31:0] GEN_489;
  wire  GEN_240;
  reg [31:0] GEN_490;
  wire [25:0] GEN_241;
  reg [31:0] GEN_491;
  wire [1:0] GEN_242;
  reg [31:0] GEN_492;
  wire [2:0] GEN_243;
  reg [31:0] GEN_493;
  wire  GEN_244;
  reg [31:0] GEN_494;
  wire [2:0] GEN_245;
  reg [31:0] GEN_495;
  wire [10:0] GEN_246;
  reg [31:0] GEN_496;
  wire [63:0] GEN_247;
  reg [63:0] GEN_497;
  wire  GEN_248;
  reg [31:0] GEN_498;
  wire  GEN_249;
  reg [31:0] GEN_499;
  wire [4:0] GEN_250;
  reg [31:0] GEN_500;
  wire  GEN_251;
  reg [31:0] GEN_501;
  wire  GEN_252;
  reg [31:0] GEN_502;
  wire  GEN_253;
  reg [31:0] GEN_503;
  wire  GEN_254;
  reg [31:0] GEN_504;
  wire  GEN_255;
  reg [31:0] GEN_505;
  wire  GEN_256;
  reg [31:0] GEN_506;
  wire  GEN_257;
  reg [31:0] GEN_507;
  wire  GEN_258;
  reg [31:0] GEN_508;
  wire  GEN_259;
  reg [31:0] GEN_509;
  wire  GEN_260;
  reg [31:0] GEN_510;
  wire  GEN_261;
  reg [31:0] GEN_511;
  wire  GEN_262;
  reg [31:0] GEN_512;
  wire  GEN_263;
  reg [31:0] GEN_513;
  wire  GEN_264;
  reg [31:0] GEN_514;
  wire  GEN_265;
  reg [31:0] GEN_515;
  wire  GEN_266;
  reg [31:0] GEN_516;
  wire [2:0] GEN_267;
  reg [31:0] GEN_517;
  wire [1:0] GEN_268;
  reg [31:0] GEN_518;
  wire [64:0] GEN_269;
  reg [95:0] GEN_519;
  wire [64:0] GEN_270;
  reg [95:0] GEN_520;
  wire [64:0] GEN_271;
  reg [95:0] GEN_521;
  wire  GEN_272;
  reg [31:0] GEN_522;
  IBuf ibuf (
    .clk(ibuf_clk),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_valid(ibuf_io_imem_bits_btb_valid),
    .io_imem_bits_btb_bits_taken(ibuf_io_imem_bits_btb_bits_taken),
    .io_imem_bits_btb_bits_mask(ibuf_io_imem_bits_btb_bits_mask),
    .io_imem_bits_btb_bits_bridx(ibuf_io_imem_bits_btb_bits_bridx),
    .io_imem_bits_btb_bits_target(ibuf_io_imem_bits_btb_bits_target),
    .io_imem_bits_btb_bits_entry(ibuf_io_imem_bits_btb_bits_entry),
    .io_imem_bits_btb_bits_bht_history(ibuf_io_imem_bits_btb_bits_bht_history),
    .io_imem_bits_btb_bits_bht_value(ibuf_io_imem_bits_btb_bits_bht_value),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_mask(ibuf_io_imem_bits_mask),
    .io_imem_bits_xcpt_if(ibuf_io_imem_bits_xcpt_if),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_btb_resp_taken(ibuf_io_btb_resp_taken),
    .io_btb_resp_mask(ibuf_io_btb_resp_mask),
    .io_btb_resp_bridx(ibuf_io_btb_resp_bridx),
    .io_btb_resp_target(ibuf_io_btb_resp_target),
    .io_btb_resp_entry(ibuf_io_btb_resp_entry),
    .io_btb_resp_bht_history(ibuf_io_btb_resp_bht_history),
    .io_btb_resp_bht_value(ibuf_io_btb_resp_bht_value),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_pf0(ibuf_io_inst_0_bits_pf0),
    .io_inst_0_bits_pf1(ibuf_io_inst_0_bits_pf1),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_btb_hit(ibuf_io_inst_0_bits_btb_hit),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3)
  );
  CSRFile csr (
    .clk(csr_clk),
    .reset(csr_reset),
    .io_prci_reset(csr_io_prci_reset),
    .io_prci_id(csr_io_prci_id),
    .io_prci_interrupts_meip(csr_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(csr_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(csr_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(csr_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(csr_io_prci_interrupts_msip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_csr_stall(csr_io_csr_stall),
    .io_csr_xcpt(csr_io_csr_xcpt),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero3(csr_io_status_zero3),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_vm(csr_io_status_vm),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_pum(csr_io_status_pum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_asid(csr_io_ptbr_asid),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fatc(csr_io_fatc),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_rocc_cmd_ready(csr_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(csr_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(csr_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(csr_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(csr_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(csr_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(csr_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(csr_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(csr_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(csr_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(csr_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(csr_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(csr_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(csr_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(csr_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(csr_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(csr_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(csr_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(csr_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(csr_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(csr_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(csr_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(csr_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(csr_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(csr_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(csr_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(csr_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(csr_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(csr_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(csr_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(csr_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(csr_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(csr_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(csr_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(csr_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(csr_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(csr_io_rocc_resp_ready),
    .io_rocc_resp_valid(csr_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(csr_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(csr_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(csr_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(csr_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(csr_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(csr_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(csr_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(csr_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(csr_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(csr_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(csr_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(csr_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(csr_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(csr_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(csr_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(csr_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(csr_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(csr_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(csr_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(csr_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(csr_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(csr_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(csr_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(csr_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(csr_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(csr_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(csr_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(csr_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(csr_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(csr_io_rocc_mem_ordered),
    .io_rocc_busy(csr_io_rocc_busy),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(csr_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(csr_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(csr_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(csr_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(csr_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(csr_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(csr_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(csr_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(csr_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(csr_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(csr_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(csr_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(csr_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(csr_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(csr_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(csr_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(csr_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(csr_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(csr_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(csr_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(csr_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(csr_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(csr_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(csr_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(csr_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(csr_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(csr_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(csr_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(csr_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(csr_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(csr_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(csr_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(csr_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(csr_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(csr_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(csr_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(csr_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(csr_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(csr_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(csr_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(csr_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(csr_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(csr_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(csr_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(csr_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(csr_io_rocc_exception),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_ttype(csr_io_bp_0_control_ttype),
    .io_bp_0_control_dmode(csr_io_bp_0_control_dmode),
    .io_bp_0_control_maskmax(csr_io_bp_0_control_maskmax),
    .io_bp_0_control_reserved(csr_io_bp_0_control_reserved),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_chain(csr_io_bp_0_control_chain),
    .io_bp_0_control_zero(csr_io_bp_0_control_zero),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address)
  );
  BreakpointUnit bpu (
    .clk(bpu_clk),
    .reset(bpu_reset),
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_status_sd(bpu_io_status_sd),
    .io_status_zero3(bpu_io_status_zero3),
    .io_status_sd_rv32(bpu_io_status_sd_rv32),
    .io_status_zero2(bpu_io_status_zero2),
    .io_status_vm(bpu_io_status_vm),
    .io_status_zero1(bpu_io_status_zero1),
    .io_status_mxr(bpu_io_status_mxr),
    .io_status_pum(bpu_io_status_pum),
    .io_status_mprv(bpu_io_status_mprv),
    .io_status_xs(bpu_io_status_xs),
    .io_status_fs(bpu_io_status_fs),
    .io_status_mpp(bpu_io_status_mpp),
    .io_status_hpp(bpu_io_status_hpp),
    .io_status_spp(bpu_io_status_spp),
    .io_status_mpie(bpu_io_status_mpie),
    .io_status_hpie(bpu_io_status_hpie),
    .io_status_spie(bpu_io_status_spie),
    .io_status_upie(bpu_io_status_upie),
    .io_status_mie(bpu_io_status_mie),
    .io_status_hie(bpu_io_status_hie),
    .io_status_sie(bpu_io_status_sie),
    .io_status_uie(bpu_io_status_uie),
    .io_bp_0_control_ttype(bpu_io_bp_0_control_ttype),
    .io_bp_0_control_dmode(bpu_io_bp_0_control_dmode),
    .io_bp_0_control_maskmax(bpu_io_bp_0_control_maskmax),
    .io_bp_0_control_reserved(bpu_io_bp_0_control_reserved),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_chain(bpu_io_bp_0_control_chain),
    .io_bp_0_control_zero(bpu_io_bp_0_control_zero),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st)
  );
  ALU alu (
    .clk(alu_clk),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clk(div_clk),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_imem_req_bits_pc = T_8325;
  assign io_imem_req_bits_speculative = T_8062;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign io_imem_btb_update_valid = T_8342;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_pc = T_8361;
  assign io_imem_btb_update_bits_target = io_imem_req_bits_pc[38:0];
  assign io_imem_btb_update_bits_taken = GEN_155;
  assign io_imem_btb_update_bits_isValid = T_8345;
  assign io_imem_btb_update_bits_isJump = T_8346;
  assign io_imem_btb_update_bits_isReturn = T_8352;
  assign io_imem_btb_update_bits_br_pc = T_8357[38:0];
  assign io_imem_bht_update_valid = T_8365;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_ras_update_valid = T_8336;
  assign io_imem_ras_update_bits_isCall = T_8370;
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_returnAddr = mem_int_wdata[38:0];
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_flush_icache = T_8329;
  assign io_imem_flush_tlb = csr_io_fatc;
  assign io_dmem_req_valid = T_8375;
  assign io_dmem_req_bits_addr = T_8400;
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_data = GEN_156;
  assign io_dmem_s1_kill = T_8402;
  assign io_dmem_s1_data = T_8401;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr_asid = csr_io_ptbr_asid;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_status_zero3 = csr_io_status_zero3;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_pum = csr_io_status_pum;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_mpp = csr_io_status_mpp;
  assign io_ptw_status_hpp = csr_io_status_hpp;
  assign io_ptw_status_spp = csr_io_status_spp;
  assign io_ptw_status_mpie = csr_io_status_mpie;
  assign io_ptw_status_hpie = csr_io_status_hpie;
  assign io_ptw_status_spie = csr_io_status_spie;
  assign io_ptw_status_upie = csr_io_status_upie;
  assign io_ptw_status_mie = csr_io_status_mie;
  assign io_ptw_status_hie = csr_io_status_hie;
  assign io_ptw_status_sie = csr_io_status_sie;
  assign io_ptw_status_uie = csr_io_status_uie;
  assign io_fpu_inst = ibuf_io_inst_0_bits_inst_bits;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = T_8374;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_valid = T_8373;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_killm = killm_common;
  assign io_fpu_cp_req_valid = GEN_157;
  assign io_fpu_cp_req_bits_cmd = GEN_158;
  assign io_fpu_cp_req_bits_ldst = GEN_159;
  assign io_fpu_cp_req_bits_wen = GEN_162;
  assign io_fpu_cp_req_bits_ren1 = GEN_163;
  assign io_fpu_cp_req_bits_ren2 = GEN_165;
  assign io_fpu_cp_req_bits_ren3 = GEN_166;
  assign io_fpu_cp_req_bits_swap12 = GEN_177;
  assign io_fpu_cp_req_bits_swap23 = GEN_178;
  assign io_fpu_cp_req_bits_single = GEN_179;
  assign io_fpu_cp_req_bits_fromint = GEN_180;
  assign io_fpu_cp_req_bits_toint = GEN_181;
  assign io_fpu_cp_req_bits_fastpipe = GEN_182;
  assign io_fpu_cp_req_bits_fma = GEN_183;
  assign io_fpu_cp_req_bits_div = GEN_184;
  assign io_fpu_cp_req_bits_sqrt = GEN_185;
  assign io_fpu_cp_req_bits_round = GEN_186;
  assign io_fpu_cp_req_bits_wflags = GEN_187;
  assign io_fpu_cp_req_bits_rm = GEN_188;
  assign io_fpu_cp_req_bits_typ = GEN_189;
  assign io_fpu_cp_req_bits_in1 = GEN_190;
  assign io_fpu_cp_req_bits_in2 = GEN_191;
  assign io_fpu_cp_req_bits_in3 = GEN_192;
  assign io_fpu_cp_resp_ready = GEN_193;
  assign io_rocc_cmd_valid = T_8417;
  assign io_rocc_cmd_bits_inst_funct = T_8439_funct;
  assign io_rocc_cmd_bits_inst_rs2 = T_8439_rs2;
  assign io_rocc_cmd_bits_inst_rs1 = T_8439_rs1;
  assign io_rocc_cmd_bits_inst_xd = T_8439_xd;
  assign io_rocc_cmd_bits_inst_xs1 = T_8439_xs1;
  assign io_rocc_cmd_bits_inst_xs2 = T_8439_xs2;
  assign io_rocc_cmd_bits_inst_rd = T_8439_rd;
  assign io_rocc_cmd_bits_inst_opcode = T_8439_opcode;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign io_rocc_cmd_bits_status_debug = csr_io_status_debug;
  assign io_rocc_cmd_bits_status_prv = csr_io_status_prv;
  assign io_rocc_cmd_bits_status_sd = csr_io_status_sd;
  assign io_rocc_cmd_bits_status_zero3 = csr_io_status_zero3;
  assign io_rocc_cmd_bits_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_rocc_cmd_bits_status_zero2 = csr_io_status_zero2;
  assign io_rocc_cmd_bits_status_vm = csr_io_status_vm;
  assign io_rocc_cmd_bits_status_zero1 = csr_io_status_zero1;
  assign io_rocc_cmd_bits_status_mxr = csr_io_status_mxr;
  assign io_rocc_cmd_bits_status_pum = csr_io_status_pum;
  assign io_rocc_cmd_bits_status_mprv = csr_io_status_mprv;
  assign io_rocc_cmd_bits_status_xs = csr_io_status_xs;
  assign io_rocc_cmd_bits_status_fs = csr_io_status_fs;
  assign io_rocc_cmd_bits_status_mpp = csr_io_status_mpp;
  assign io_rocc_cmd_bits_status_hpp = csr_io_status_hpp;
  assign io_rocc_cmd_bits_status_spp = csr_io_status_spp;
  assign io_rocc_cmd_bits_status_mpie = csr_io_status_mpie;
  assign io_rocc_cmd_bits_status_hpie = csr_io_status_hpie;
  assign io_rocc_cmd_bits_status_spie = csr_io_status_spie;
  assign io_rocc_cmd_bits_status_upie = csr_io_status_upie;
  assign io_rocc_cmd_bits_status_mie = csr_io_status_mie;
  assign io_rocc_cmd_bits_status_hie = csr_io_status_hie;
  assign io_rocc_cmd_bits_status_sie = csr_io_status_sie;
  assign io_rocc_cmd_bits_status_uie = csr_io_status_uie;
  assign io_rocc_resp_ready = GEN_194;
  assign io_rocc_mem_req_ready = GEN_195;
  assign io_rocc_mem_s2_nack = GEN_196;
  assign io_rocc_mem_resp_valid = GEN_197;
  assign io_rocc_mem_resp_bits_addr = GEN_198;
  assign io_rocc_mem_resp_bits_tag = GEN_199;
  assign io_rocc_mem_resp_bits_cmd = GEN_200;
  assign io_rocc_mem_resp_bits_typ = GEN_201;
  assign io_rocc_mem_resp_bits_data = GEN_202;
  assign io_rocc_mem_resp_bits_replay = GEN_203;
  assign io_rocc_mem_resp_bits_has_data = GEN_204;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_205;
  assign io_rocc_mem_resp_bits_store_data = GEN_206;
  assign io_rocc_mem_replay_next = GEN_207;
  assign io_rocc_mem_xcpt_ma_ld = GEN_208;
  assign io_rocc_mem_xcpt_ma_st = GEN_209;
  assign io_rocc_mem_xcpt_pf_ld = GEN_210;
  assign io_rocc_mem_xcpt_pf_st = GEN_211;
  assign io_rocc_mem_ordered = GEN_212;
  assign io_rocc_autl_acquire_ready = GEN_213;
  assign io_rocc_autl_grant_valid = GEN_214;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_215;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_216;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_217;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_218;
  assign io_rocc_autl_grant_bits_g_type = GEN_219;
  assign io_rocc_autl_grant_bits_data = GEN_220;
  assign io_rocc_fpu_req_ready = GEN_221;
  assign io_rocc_fpu_resp_valid = GEN_222;
  assign io_rocc_fpu_resp_bits_data = GEN_223;
  assign io_rocc_fpu_resp_bits_exc = GEN_224;
  assign io_rocc_exception = T_8420;
  assign take_pc_mem = T_7989;
  assign take_pc_wb = T_8079;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign ibuf_clk = clk;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_imem_bits_btb_valid = io_imem_resp_bits_btb_valid;
  assign ibuf_io_imem_bits_btb_bits_taken = io_imem_resp_bits_btb_bits_taken;
  assign ibuf_io_imem_bits_btb_bits_mask = io_imem_resp_bits_btb_bits_mask;
  assign ibuf_io_imem_bits_btb_bits_bridx = io_imem_resp_bits_btb_bits_bridx;
  assign ibuf_io_imem_bits_btb_bits_target = io_imem_resp_bits_btb_bits_target;
  assign ibuf_io_imem_bits_btb_bits_entry = io_imem_resp_bits_btb_bits_entry;
  assign ibuf_io_imem_bits_btb_bits_bht_history = io_imem_resp_bits_btb_bits_bht_history;
  assign ibuf_io_imem_bits_btb_bits_bht_value = io_imem_resp_bits_btb_bits_bht_value;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_mask = io_imem_resp_bits_mask;
  assign ibuf_io_imem_bits_xcpt_if = io_imem_resp_bits_xcpt_if;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_kill = take_pc_mem_wb;
  assign ibuf_io_inst_0_ready = T_8332;
  assign id_ctrl_legal = T_6845;
  assign id_ctrl_fp = T_6856;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_branch = T_6861;
  assign id_ctrl_jal = T_6867;
  assign id_ctrl_jalr = T_6873;
  assign id_ctrl_rxs2 = T_6891;
  assign id_ctrl_rxs1 = T_6917;
  assign id_ctrl_sel_alu2 = T_6961;
  assign id_ctrl_sel_alu1 = T_6987;
  assign id_ctrl_sel_imm = T_7023;
  assign id_ctrl_alu_dw = T_7034;
  assign id_ctrl_alu_fn = T_7118;
  assign id_ctrl_mem = T_7139;
  assign id_ctrl_mem_cmd = T_7199;
  assign id_ctrl_mem_type = T_7219;
  assign id_ctrl_rfs1 = T_7235;
  assign id_ctrl_rfs2 = T_7252;
  assign id_ctrl_rfs3 = T_7231;
  assign id_ctrl_wfd = T_7267;
  assign id_ctrl_div = T_7271;
  assign id_ctrl_wxd = T_7309;
  assign id_ctrl_csr = T_7329;
  assign id_ctrl_fence_i = T_7333;
  assign id_ctrl_fence = T_7339;
  assign id_ctrl_amo = T_7345;
  assign T_6645 = ibuf_io_inst_0_bits_inst_bits & 32'h207f;
  assign T_6647 = T_6645 == 32'h3;
  assign T_6649 = ibuf_io_inst_0_bits_inst_bits & 32'h106f;
  assign T_6651 = T_6649 == 32'h3;
  assign T_6653 = ibuf_io_inst_0_bits_inst_bits & 32'h607f;
  assign T_6655 = T_6653 == 32'hf;
  assign T_6657 = ibuf_io_inst_0_bits_inst_bits & 32'h7077;
  assign T_6659 = T_6657 == 32'h13;
  assign T_6661 = ibuf_io_inst_0_bits_inst_bits & 32'h5f;
  assign T_6663 = T_6661 == 32'h17;
  assign T_6665 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00007f;
  assign T_6667 = T_6665 == 32'h33;
  assign T_6669 = ibuf_io_inst_0_bits_inst_bits & 32'hbe007077;
  assign T_6671 = T_6669 == 32'h33;
  assign T_6673 = ibuf_io_inst_0_bits_inst_bits & 32'h4000073;
  assign T_6675 = T_6673 == 32'h43;
  assign T_6677 = ibuf_io_inst_0_bits_inst_bits & 32'he400007f;
  assign T_6679 = T_6677 == 32'h53;
  assign T_6681 = ibuf_io_inst_0_bits_inst_bits & 32'h707b;
  assign T_6683 = T_6681 == 32'h63;
  assign T_6685 = ibuf_io_inst_0_bits_inst_bits & 32'h7f;
  assign T_6687 = T_6685 == 32'h6f;
  assign T_6689 = ibuf_io_inst_0_bits_inst_bits & 32'hffefffff;
  assign T_6691 = T_6689 == 32'h73;
  assign T_6693 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00305f;
  assign T_6695 = T_6693 == 32'h1013;
  assign T_6697 = ibuf_io_inst_0_bits_inst_bits & 32'hfe00305f;
  assign T_6699 = T_6697 == 32'h101b;
  assign T_6701 = ibuf_io_inst_0_bits_inst_bits & 32'h605b;
  assign T_6703 = T_6701 == 32'h2003;
  assign T_6707 = T_6645 == 32'h2013;
  assign T_6709 = ibuf_io_inst_0_bits_inst_bits & 32'h1800607f;
  assign T_6711 = T_6709 == 32'h202f;
  assign T_6715 = T_6645 == 32'h2073;
  assign T_6717 = ibuf_io_inst_0_bits_inst_bits & 32'hbc00707f;
  assign T_6719 = T_6717 == 32'h5013;
  assign T_6721 = ibuf_io_inst_0_bits_inst_bits & 32'hbe00705f;
  assign T_6723 = T_6721 == 32'h501b;
  assign T_6727 = T_6669 == 32'h5033;
  assign T_6729 = ibuf_io_inst_0_bits_inst_bits & 32'hfe004077;
  assign T_6731 = T_6729 == 32'h2004033;
  assign T_6733 = ibuf_io_inst_0_bits_inst_bits & 32'he800607f;
  assign T_6735 = T_6733 == 32'h800202f;
  assign T_6737 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0607f;
  assign T_6739 = T_6737 == 32'h1000202f;
  assign T_6741 = ibuf_io_inst_0_bits_inst_bits & 32'hdfffffff;
  assign T_6743 = T_6741 == 32'h10200073;
  assign T_6745 = ibuf_io_inst_0_bits_inst_bits & 32'hfff07fff;
  assign T_6747 = T_6745 == 32'h10400073;
  assign T_6749 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073;
  assign T_6751 = ibuf_io_inst_0_bits_inst_bits & 32'hf400607f;
  assign T_6753 = T_6751 == 32'h20000053;
  assign T_6755 = ibuf_io_inst_0_bits_inst_bits & 32'h7c00607f;
  assign T_6757 = T_6755 == 32'h20000053;
  assign T_6759 = ibuf_io_inst_0_bits_inst_bits & 32'h7c00507f;
  assign T_6761 = T_6759 == 32'h20000053;
  assign T_6763 = ibuf_io_inst_0_bits_inst_bits & 32'h7ff0007f;
  assign T_6765 = T_6763 == 32'h40100053;
  assign T_6769 = T_6763 == 32'h42000053;
  assign T_6771 = ibuf_io_inst_0_bits_inst_bits & 32'hfdf0007f;
  assign T_6773 = T_6771 == 32'h58000053;
  assign T_6775 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073;
  assign T_6777 = ibuf_io_inst_0_bits_inst_bits & 32'hedc0007f;
  assign T_6779 = T_6777 == 32'hc0000053;
  assign T_6781 = ibuf_io_inst_0_bits_inst_bits & 32'hfdf0607f;
  assign T_6783 = T_6781 == 32'he0000053;
  assign T_6785 = ibuf_io_inst_0_bits_inst_bits & 32'hedf0707f;
  assign T_6787 = T_6785 == 32'he0000053;
  assign T_6789 = ibuf_io_inst_0_bits_inst_bits & 32'h603f;
  assign T_6791 = T_6789 == 32'h23;
  assign T_6793 = ibuf_io_inst_0_bits_inst_bits & 32'h306f;
  assign T_6795 = T_6793 == 32'h1063;
  assign T_6797 = ibuf_io_inst_0_bits_inst_bits & 32'h407f;
  assign T_6799 = T_6797 == 32'h4063;
  assign T_6801 = ibuf_io_inst_0_bits_inst_bits & 32'hfc007077;
  assign T_6803 = T_6801 == 32'h33;
  assign T_6806 = T_6647 | T_6651;
  assign T_6807 = T_6806 | T_6655;
  assign T_6808 = T_6807 | T_6659;
  assign T_6809 = T_6808 | T_6663;
  assign T_6810 = T_6809 | T_6667;
  assign T_6811 = T_6810 | T_6671;
  assign T_6812 = T_6811 | T_6675;
  assign T_6813 = T_6812 | T_6679;
  assign T_6814 = T_6813 | T_6683;
  assign T_6815 = T_6814 | T_6687;
  assign T_6816 = T_6815 | T_6691;
  assign T_6817 = T_6816 | T_6695;
  assign T_6818 = T_6817 | T_6699;
  assign T_6819 = T_6818 | T_6703;
  assign T_6820 = T_6819 | T_6707;
  assign T_6821 = T_6820 | T_6711;
  assign T_6822 = T_6821 | T_6715;
  assign T_6823 = T_6822 | T_6719;
  assign T_6824 = T_6823 | T_6723;
  assign T_6825 = T_6824 | T_6727;
  assign T_6826 = T_6825 | T_6731;
  assign T_6827 = T_6826 | T_6735;
  assign T_6828 = T_6827 | T_6739;
  assign T_6829 = T_6828 | T_6743;
  assign T_6830 = T_6829 | T_6747;
  assign T_6831 = T_6830 | T_6749;
  assign T_6832 = T_6831 | T_6753;
  assign T_6833 = T_6832 | T_6757;
  assign T_6834 = T_6833 | T_6761;
  assign T_6835 = T_6834 | T_6765;
  assign T_6836 = T_6835 | T_6769;
  assign T_6837 = T_6836 | T_6773;
  assign T_6838 = T_6837 | T_6775;
  assign T_6839 = T_6838 | T_6779;
  assign T_6840 = T_6839 | T_6783;
  assign T_6841 = T_6840 | T_6787;
  assign T_6842 = T_6841 | T_6791;
  assign T_6843 = T_6842 | T_6795;
  assign T_6844 = T_6843 | T_6799;
  assign T_6845 = T_6844 | T_6803;
  assign T_6847 = ibuf_io_inst_0_bits_inst_bits & 32'h5c;
  assign T_6849 = T_6847 == 32'h4;
  assign T_6851 = ibuf_io_inst_0_bits_inst_bits & 32'h60;
  assign T_6853 = T_6851 == 32'h40;
  assign T_6856 = T_6849 | T_6853;
  assign T_6859 = ibuf_io_inst_0_bits_inst_bits & 32'h74;
  assign T_6861 = T_6859 == 32'h60;
  assign T_6865 = ibuf_io_inst_0_bits_inst_bits & 32'h68;
  assign T_6867 = T_6865 == 32'h68;
  assign T_6871 = ibuf_io_inst_0_bits_inst_bits & 32'h203c;
  assign T_6873 = T_6871 == 32'h24;
  assign T_6877 = ibuf_io_inst_0_bits_inst_bits & 32'h64;
  assign T_6879 = T_6877 == 32'h20;
  assign T_6881 = ibuf_io_inst_0_bits_inst_bits & 32'h34;
  assign T_6883 = T_6881 == 32'h20;
  assign T_6885 = ibuf_io_inst_0_bits_inst_bits & 32'h2048;
  assign T_6887 = T_6885 == 32'h2008;
  assign T_6890 = T_6879 | T_6883;
  assign T_6891 = T_6890 | T_6887;
  assign T_6893 = ibuf_io_inst_0_bits_inst_bits & 32'h44;
  assign T_6895 = T_6893 == 32'h0;
  assign T_6897 = ibuf_io_inst_0_bits_inst_bits & 32'h4024;
  assign T_6899 = T_6897 == 32'h20;
  assign T_6901 = ibuf_io_inst_0_bits_inst_bits & 32'h38;
  assign T_6903 = T_6901 == 32'h20;
  assign T_6905 = ibuf_io_inst_0_bits_inst_bits & 32'h2050;
  assign T_6907 = T_6905 == 32'h2000;
  assign T_6909 = ibuf_io_inst_0_bits_inst_bits & 32'h90000034;
  assign T_6911 = T_6909 == 32'h90000010;
  assign T_6914 = T_6895 | T_6899;
  assign T_6915 = T_6914 | T_6903;
  assign T_6916 = T_6915 | T_6907;
  assign T_6917 = T_6916 | T_6911;
  assign T_6919 = ibuf_io_inst_0_bits_inst_bits & 32'h58;
  assign T_6921 = T_6919 == 32'h0;
  assign T_6923 = ibuf_io_inst_0_bits_inst_bits & 32'h20;
  assign T_6925 = T_6923 == 32'h0;
  assign T_6927 = ibuf_io_inst_0_bits_inst_bits & 32'hc;
  assign T_6929 = T_6927 == 32'h4;
  assign T_6931 = ibuf_io_inst_0_bits_inst_bits & 32'h48;
  assign T_6933 = T_6931 == 32'h48;
  assign T_6935 = ibuf_io_inst_0_bits_inst_bits & 32'h4050;
  assign T_6937 = T_6935 == 32'h4050;
  assign T_6940 = T_6921 | T_6925;
  assign T_6941 = T_6940 | T_6929;
  assign T_6942 = T_6941 | T_6933;
  assign T_6943 = T_6942 | T_6937;
  assign T_6947 = T_6931 == 32'h0;
  assign T_6949 = ibuf_io_inst_0_bits_inst_bits & 32'h18;
  assign T_6951 = T_6949 == 32'h0;
  assign T_6953 = ibuf_io_inst_0_bits_inst_bits & 32'h4008;
  assign T_6955 = T_6953 == 32'h4000;
  assign T_6958 = T_6947 | T_6895;
  assign T_6959 = T_6958 | T_6951;
  assign T_6960 = T_6959 | T_6955;
  assign T_6961 = {T_6960,T_6943};
  assign T_6963 = ibuf_io_inst_0_bits_inst_bits & 32'h4004;
  assign T_6965 = T_6963 == 32'h0;
  assign T_6967 = ibuf_io_inst_0_bits_inst_bits & 32'h50;
  assign T_6969 = T_6967 == 32'h0;
  assign T_6971 = ibuf_io_inst_0_bits_inst_bits & 32'h24;
  assign T_6973 = T_6971 == 32'h0;
  assign T_6976 = T_6965 | T_6969;
  assign T_6977 = T_6976 | T_6895;
  assign T_6978 = T_6977 | T_6973;
  assign T_6979 = T_6978 | T_6951;
  assign T_6983 = T_6881 == 32'h14;
  assign T_6986 = T_6983 | T_6933;
  assign T_6987 = {T_6986,T_6979};
  assign T_6991 = T_6949 == 32'h8;
  assign T_6995 = T_6893 == 32'h40;
  assign T_6998 = T_6991 | T_6995;
  assign T_7000 = ibuf_io_inst_0_bits_inst_bits & 32'h14;
  assign T_7002 = T_7000 == 32'h14;
  assign T_7005 = T_6991 | T_7002;
  assign T_7007 = ibuf_io_inst_0_bits_inst_bits & 32'h30;
  assign T_7009 = T_7007 == 32'h0;
  assign T_7011 = ibuf_io_inst_0_bits_inst_bits & 32'h201c;
  assign T_7013 = T_7011 == 32'h4;
  assign T_7017 = T_7000 == 32'h10;
  assign T_7020 = T_7009 | T_7013;
  assign T_7021 = T_7020 | T_7017;
  assign T_7022 = {T_7021,T_7005};
  assign T_7023 = {T_7022,T_6998};
  assign T_7025 = ibuf_io_inst_0_bits_inst_bits & 32'h10;
  assign T_7027 = T_7025 == 32'h0;
  assign T_7029 = ibuf_io_inst_0_bits_inst_bits & 32'h8;
  assign T_7031 = T_7029 == 32'h0;
  assign T_7034 = T_7027 | T_7031;
  assign T_7036 = ibuf_io_inst_0_bits_inst_bits & 32'h3054;
  assign T_7038 = T_7036 == 32'h1010;
  assign T_7040 = ibuf_io_inst_0_bits_inst_bits & 32'h1058;
  assign T_7042 = T_7040 == 32'h1040;
  assign T_7044 = ibuf_io_inst_0_bits_inst_bits & 32'h7044;
  assign T_7046 = T_7044 == 32'h7000;
  assign T_7049 = T_7038 | T_7042;
  assign T_7050 = T_7049 | T_7046;
  assign T_7052 = ibuf_io_inst_0_bits_inst_bits & 32'h4054;
  assign T_7054 = T_7052 == 32'h40;
  assign T_7056 = ibuf_io_inst_0_bits_inst_bits & 32'h2058;
  assign T_7058 = T_7056 == 32'h2040;
  assign T_7062 = T_7036 == 32'h3010;
  assign T_7064 = ibuf_io_inst_0_bits_inst_bits & 32'h6054;
  assign T_7066 = T_7064 == 32'h6010;
  assign T_7068 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034;
  assign T_7070 = T_7068 == 32'h40000030;
  assign T_7072 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054;
  assign T_7074 = T_7072 == 32'h40001010;
  assign T_7077 = T_7054 | T_7058;
  assign T_7078 = T_7077 | T_7062;
  assign T_7079 = T_7078 | T_7066;
  assign T_7080 = T_7079 | T_7070;
  assign T_7081 = T_7080 | T_7074;
  assign T_7083 = ibuf_io_inst_0_bits_inst_bits & 32'h2054;
  assign T_7085 = T_7083 == 32'h2010;
  assign T_7087 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054;
  assign T_7089 = T_7087 == 32'h4010;
  assign T_7091 = ibuf_io_inst_0_bits_inst_bits & 32'h5054;
  assign T_7093 = T_7091 == 32'h4010;
  assign T_7095 = ibuf_io_inst_0_bits_inst_bits & 32'h4058;
  assign T_7097 = T_7095 == 32'h4040;
  assign T_7100 = T_7085 | T_7089;
  assign T_7101 = T_7100 | T_7093;
  assign T_7102 = T_7101 | T_7097;
  assign T_7106 = T_7064 == 32'h2010;
  assign T_7108 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054;
  assign T_7110 = T_7108 == 32'h40001010;
  assign T_7113 = T_7106 | T_7097;
  assign T_7114 = T_7113 | T_7070;
  assign T_7115 = T_7114 | T_7110;
  assign T_7116 = {T_7081,T_7050};
  assign T_7117 = {T_7115,T_7102};
  assign T_7118 = {T_7117,T_7116};
  assign T_7120 = ibuf_io_inst_0_bits_inst_bits & 32'h405f;
  assign T_7122 = T_7120 == 32'h3;
  assign T_7124 = ibuf_io_inst_0_bits_inst_bits & 32'h107f;
  assign T_7126 = T_7124 == 32'h3;
  assign T_7128 = ibuf_io_inst_0_bits_inst_bits & 32'h707f;
  assign T_7130 = T_7128 == 32'h100f;
  assign T_7133 = T_7122 | T_6647;
  assign T_7134 = T_7133 | T_7126;
  assign T_7135 = T_7134 | T_7130;
  assign T_7136 = T_7135 | T_6703;
  assign T_7137 = T_7136 | T_6711;
  assign T_7138 = T_7137 | T_6735;
  assign T_7139 = T_7138 | T_6739;
  assign T_7141 = ibuf_io_inst_0_bits_inst_bits & 32'h2008;
  assign T_7143 = T_7141 == 32'h8;
  assign T_7145 = ibuf_io_inst_0_bits_inst_bits & 32'h28;
  assign T_7147 = T_7145 == 32'h20;
  assign T_7149 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020;
  assign T_7151 = T_7149 == 32'h18000020;
  assign T_7153 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020;
  assign T_7155 = T_7153 == 32'h20000020;
  assign T_7158 = T_7143 | T_7147;
  assign T_7159 = T_7158 | T_7151;
  assign T_7160 = T_7159 | T_7155;
  assign T_7162 = ibuf_io_inst_0_bits_inst_bits & 32'h10002008;
  assign T_7164 = T_7162 == 32'h10002008;
  assign T_7166 = ibuf_io_inst_0_bits_inst_bits & 32'h40002008;
  assign T_7168 = T_7166 == 32'h40002008;
  assign T_7171 = T_7164 | T_7168;
  assign T_7173 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008;
  assign T_7175 = T_7173 == 32'h8000008;
  assign T_7177 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008;
  assign T_7179 = T_7177 == 32'h10000008;
  assign T_7181 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008;
  assign T_7183 = T_7181 == 32'h80000008;
  assign T_7186 = T_7143 | T_7175;
  assign T_7187 = T_7186 | T_7179;
  assign T_7188 = T_7187 | T_7183;
  assign T_7190 = ibuf_io_inst_0_bits_inst_bits & 32'h18002008;
  assign T_7192 = T_7190 == 32'h2008;
  assign T_7196 = {T_7171,T_7160};
  assign T_7197 = {1'h0,T_7192};
  assign T_7198 = {T_7197,T_7188};
  assign T_7199 = {T_7198,T_7196};
  assign T_7201 = ibuf_io_inst_0_bits_inst_bits & 32'h1000;
  assign T_7203 = T_7201 == 32'h1000;
  assign T_7207 = ibuf_io_inst_0_bits_inst_bits & 32'h2000;
  assign T_7209 = T_7207 == 32'h2000;
  assign T_7213 = ibuf_io_inst_0_bits_inst_bits & 32'h4000;
  assign T_7215 = T_7213 == 32'h4000;
  assign T_7218 = {T_7215,T_7209};
  assign T_7219 = {T_7218,T_7203};
  assign T_7221 = ibuf_io_inst_0_bits_inst_bits & 32'h80000060;
  assign T_7223 = T_7221 == 32'h40;
  assign T_7225 = ibuf_io_inst_0_bits_inst_bits & 32'h10000060;
  assign T_7227 = T_7225 == 32'h40;
  assign T_7229 = ibuf_io_inst_0_bits_inst_bits & 32'h70;
  assign T_7231 = T_7229 == 32'h40;
  assign T_7234 = T_7223 | T_7227;
  assign T_7235 = T_7234 | T_7231;
  assign T_7237 = ibuf_io_inst_0_bits_inst_bits & 32'h7c;
  assign T_7239 = T_7237 == 32'h24;
  assign T_7241 = ibuf_io_inst_0_bits_inst_bits & 32'h40000060;
  assign T_7243 = T_7241 == 32'h40;
  assign T_7245 = ibuf_io_inst_0_bits_inst_bits & 32'h90000060;
  assign T_7247 = T_7245 == 32'h10000040;
  assign T_7250 = T_7239 | T_7243;
  assign T_7251 = T_7250 | T_7231;
  assign T_7252 = T_7251 | T_7247;
  assign T_7256 = ibuf_io_inst_0_bits_inst_bits & 32'h3c;
  assign T_7258 = T_7256 == 32'h4;
  assign T_7262 = T_7225 == 32'h10000040;
  assign T_7265 = T_7258 | T_7223;
  assign T_7266 = T_7265 | T_7231;
  assign T_7267 = T_7266 | T_7262;
  assign T_7269 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074;
  assign T_7271 = T_7269 == 32'h2000030;
  assign T_7277 = T_6877 == 32'h0;
  assign T_7281 = T_6967 == 32'h10;
  assign T_7283 = ibuf_io_inst_0_bits_inst_bits & 32'h2024;
  assign T_7285 = T_7283 == 32'h24;
  assign T_7289 = T_7145 == 32'h28;
  assign T_7291 = ibuf_io_inst_0_bits_inst_bits & 32'h1030;
  assign T_7293 = T_7291 == 32'h1030;
  assign T_7295 = ibuf_io_inst_0_bits_inst_bits & 32'h2030;
  assign T_7297 = T_7295 == 32'h2030;
  assign T_7299 = ibuf_io_inst_0_bits_inst_bits & 32'h90000010;
  assign T_7301 = T_7299 == 32'h80000010;
  assign T_7304 = T_7277 | T_7281;
  assign T_7305 = T_7304 | T_7285;
  assign T_7306 = T_7305 | T_7289;
  assign T_7307 = T_7306 | T_7293;
  assign T_7308 = T_7307 | T_7297;
  assign T_7309 = T_7308 | T_7301;
  assign T_7311 = ibuf_io_inst_0_bits_inst_bits & 32'h1070;
  assign T_7313 = T_7311 == 32'h1070;
  assign T_7317 = ibuf_io_inst_0_bits_inst_bits & 32'h2070;
  assign T_7319 = T_7317 == 32'h2070;
  assign T_7323 = ibuf_io_inst_0_bits_inst_bits & 32'h3070;
  assign T_7325 = T_7323 == 32'h70;
  assign T_7328 = {T_7325,T_7319};
  assign T_7329 = {T_7328,T_7313};
  assign T_7331 = ibuf_io_inst_0_bits_inst_bits & 32'h3058;
  assign T_7333 = T_7331 == 32'h1008;
  assign T_7339 = T_7331 == 32'h8;
  assign T_7343 = ibuf_io_inst_0_bits_inst_bits & 32'h6048;
  assign T_7345 = T_7343 == 32'h2008;
  assign id_load_use = T_8225;
  assign T_7352_T_7361_addr = T_7360;
  assign T_7352_T_7361_en = 1'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_7352_T_7361_data = T_7352[T_7352_T_7361_addr];
  `else
  assign T_7352_T_7361_data = T_7352_T_7361_addr >= 5'h1f ? GEN_401[63:0] : T_7352[T_7352_T_7361_addr];
  `endif
  assign T_7352_T_7371_addr = T_7370;
  assign T_7352_T_7371_en = 1'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign T_7352_T_7371_data = T_7352[T_7352_T_7371_addr];
  `else
  assign T_7352_T_7371_data = T_7352_T_7371_addr >= 5'h1f ? GEN_402[63:0] : T_7352[T_7352_T_7371_addr];
  `endif
  assign T_7352_T_8104_data = rf_wdata;
  assign T_7352_T_8104_addr = T_8103;
  assign T_7352_T_8104_mask = GEN_164;
  assign T_7352_T_8104_en = GEN_164;
  assign id_rs_0 = GEN_167;
  assign T_7356 = ibuf_io_inst_0_bits_inst_rs1 == 5'h0;
  assign T_7359 = ibuf_io_inst_0_bits_inst_rs1;
  assign T_7360 = ~ T_7359;
  assign T_7362 = T_7352_T_7361_data;
  assign id_rs_1 = GEN_168;
  assign T_7369 = ibuf_io_inst_0_bits_inst_rs2;
  assign T_7370 = ~ T_7369;
  assign T_7372 = T_7352_T_7371_data;
  assign ctrl_killd = T_8320;
  assign csr_clk = clk;
  assign csr_reset = reset;
  assign csr_io_prci_reset = io_prci_reset;
  assign csr_io_prci_id = io_prci_id;
  assign csr_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign csr_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign csr_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign csr_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign csr_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign csr_io_rw_addr = T_8131;
  assign csr_io_rw_cmd = T_8132;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_exception = wb_reg_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_cause = wb_reg_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = T_8130;
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_rocc_cmd_ready = GEN_225;
  assign csr_io_rocc_resp_valid = GEN_226;
  assign csr_io_rocc_resp_bits_rd = GEN_227;
  assign csr_io_rocc_resp_bits_data = GEN_228;
  assign csr_io_rocc_mem_req_valid = GEN_229;
  assign csr_io_rocc_mem_req_bits_addr = GEN_230;
  assign csr_io_rocc_mem_req_bits_tag = GEN_231;
  assign csr_io_rocc_mem_req_bits_cmd = GEN_232;
  assign csr_io_rocc_mem_req_bits_typ = GEN_233;
  assign csr_io_rocc_mem_req_bits_phys = GEN_234;
  assign csr_io_rocc_mem_req_bits_data = GEN_235;
  assign csr_io_rocc_mem_s1_kill = GEN_236;
  assign csr_io_rocc_mem_s1_data = GEN_237;
  assign csr_io_rocc_mem_invalidate_lr = GEN_238;
  assign csr_io_rocc_busy = GEN_239;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign csr_io_rocc_autl_acquire_valid = GEN_240;
  assign csr_io_rocc_autl_acquire_bits_addr_block = GEN_241;
  assign csr_io_rocc_autl_acquire_bits_client_xact_id = GEN_242;
  assign csr_io_rocc_autl_acquire_bits_addr_beat = GEN_243;
  assign csr_io_rocc_autl_acquire_bits_is_builtin_type = GEN_244;
  assign csr_io_rocc_autl_acquire_bits_a_type = GEN_245;
  assign csr_io_rocc_autl_acquire_bits_union = GEN_246;
  assign csr_io_rocc_autl_acquire_bits_data = GEN_247;
  assign csr_io_rocc_autl_grant_ready = GEN_248;
  assign csr_io_rocc_fpu_req_valid = GEN_249;
  assign csr_io_rocc_fpu_req_bits_cmd = GEN_250;
  assign csr_io_rocc_fpu_req_bits_ldst = GEN_251;
  assign csr_io_rocc_fpu_req_bits_wen = GEN_252;
  assign csr_io_rocc_fpu_req_bits_ren1 = GEN_253;
  assign csr_io_rocc_fpu_req_bits_ren2 = GEN_254;
  assign csr_io_rocc_fpu_req_bits_ren3 = GEN_255;
  assign csr_io_rocc_fpu_req_bits_swap12 = GEN_256;
  assign csr_io_rocc_fpu_req_bits_swap23 = GEN_257;
  assign csr_io_rocc_fpu_req_bits_single = GEN_258;
  assign csr_io_rocc_fpu_req_bits_fromint = GEN_259;
  assign csr_io_rocc_fpu_req_bits_toint = GEN_260;
  assign csr_io_rocc_fpu_req_bits_fastpipe = GEN_261;
  assign csr_io_rocc_fpu_req_bits_fma = GEN_262;
  assign csr_io_rocc_fpu_req_bits_div = GEN_263;
  assign csr_io_rocc_fpu_req_bits_sqrt = GEN_264;
  assign csr_io_rocc_fpu_req_bits_round = GEN_265;
  assign csr_io_rocc_fpu_req_bits_wflags = GEN_266;
  assign csr_io_rocc_fpu_req_bits_rm = GEN_267;
  assign csr_io_rocc_fpu_req_bits_typ = GEN_268;
  assign csr_io_rocc_fpu_req_bits_in1 = GEN_269;
  assign csr_io_rocc_fpu_req_bits_in2 = GEN_270;
  assign csr_io_rocc_fpu_req_bits_in3 = GEN_271;
  assign csr_io_rocc_fpu_resp_ready = GEN_272;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign T_7374 = id_ctrl_csr == 3'h2;
  assign T_7375 = id_ctrl_csr == 3'h3;
  assign T_7376 = T_7374 | T_7375;
  assign id_csr_ren = T_7376 & T_7356;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_csr_addr = ibuf_io_inst_0_bits_inst_bits[31:20];
  assign T_7380 = id_csr_ren == 1'h0;
  assign T_7381 = id_csr_en & T_7380;
  assign T_7511 = id_csr_addr & 12'h46;
  assign T_7513 = T_7511 == 12'h40;
  assign T_7515 = id_csr_addr & 12'h244;
  assign T_7517 = T_7515 == 12'h240;
  assign T_7520 = T_7513 | T_7517;
  assign T_7523 = T_7520 == 1'h0;
  assign T_7524 = T_7381 & T_7523;
  assign id_csr_flush = id_system_insn | T_7524;
  assign T_7526 = id_ctrl_legal == 1'h0;
  assign T_7528 = csr_io_status_fs != 2'h0;
  assign T_7530 = T_7528 == 1'h0;
  assign T_7531 = id_ctrl_fp & T_7530;
  assign T_7532 = T_7526 | T_7531;
  assign T_7534 = csr_io_status_xs != 2'h0;
  assign T_7536 = T_7534 == 1'h0;
  assign T_7537 = id_ctrl_rocc & T_7536;
  assign id_illegal_insn = T_7532 | T_7537;
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26];
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25];
  assign T_7538 = id_ctrl_amo & id_amo_rl;
  assign id_fence_next = id_ctrl_fence | T_7538;
  assign T_7540 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = T_7540 | io_dmem_req_valid;
  assign T_7546 = wb_reg_valid & wb_ctrl_rocc;
  assign T_7548 = id_reg_fence & id_mem_busy;
  assign T_7549 = id_fence_next | T_7548;
  assign T_7551 = id_ctrl_amo & id_amo_aq;
  assign T_7552 = T_7551 | id_ctrl_fence_i;
  assign T_7553 = id_ctrl_mem | id_ctrl_rocc;
  assign T_7554 = id_reg_fence & T_7553;
  assign T_7555 = T_7552 | T_7554;
  assign T_7556 = T_7555 | id_csr_en;
  assign T_7557 = id_mem_busy & T_7556;
  assign bpu_clk = clk;
  assign bpu_reset = reset;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_status_sd = csr_io_status_sd;
  assign bpu_io_status_zero3 = csr_io_status_zero3;
  assign bpu_io_status_sd_rv32 = csr_io_status_sd_rv32;
  assign bpu_io_status_zero2 = csr_io_status_zero2;
  assign bpu_io_status_vm = csr_io_status_vm;
  assign bpu_io_status_zero1 = csr_io_status_zero1;
  assign bpu_io_status_mxr = csr_io_status_mxr;
  assign bpu_io_status_pum = csr_io_status_pum;
  assign bpu_io_status_mprv = csr_io_status_mprv;
  assign bpu_io_status_xs = csr_io_status_xs;
  assign bpu_io_status_fs = csr_io_status_fs;
  assign bpu_io_status_mpp = csr_io_status_mpp;
  assign bpu_io_status_hpp = csr_io_status_hpp;
  assign bpu_io_status_spp = csr_io_status_spp;
  assign bpu_io_status_mpie = csr_io_status_mpie;
  assign bpu_io_status_hpie = csr_io_status_hpie;
  assign bpu_io_status_spie = csr_io_status_spie;
  assign bpu_io_status_upie = csr_io_status_upie;
  assign bpu_io_status_mie = csr_io_status_mie;
  assign bpu_io_status_hie = csr_io_status_hie;
  assign bpu_io_status_sie = csr_io_status_sie;
  assign bpu_io_status_uie = csr_io_status_uie;
  assign bpu_io_bp_0_control_ttype = csr_io_bp_0_control_ttype;
  assign bpu_io_bp_0_control_dmode = csr_io_bp_0_control_dmode;
  assign bpu_io_bp_0_control_maskmax = csr_io_bp_0_control_maskmax;
  assign bpu_io_bp_0_control_reserved = csr_io_bp_0_control_reserved;
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action;
  assign bpu_io_bp_0_control_chain = csr_io_bp_0_control_chain;
  assign bpu_io_bp_0_control_zero = csr_io_bp_0_control_zero;
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = ibuf_io_pc[38:0];
  assign bpu_io_ea = mem_reg_wdata[38:0];
  assign id_xcpt_if = ibuf_io_inst_0_bits_pf0 | ibuf_io_inst_0_bits_pf1;
  assign T_7562 = csr_io_interrupt | bpu_io_debug_if;
  assign T_7563 = T_7562 | bpu_io_xcpt_if;
  assign T_7564 = T_7563 | id_xcpt_if;
  assign id_xcpt = T_7564 | id_illegal_insn;
  assign T_7565 = id_xcpt_if ? 2'h1 : 2'h2;
  assign T_7566 = bpu_io_xcpt_if ? 2'h3 : T_7565;
  assign T_7567 = bpu_io_debug_if ? 4'hd : {{2'd0}, T_7566};
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{60'd0}, T_7567};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign T_7571 = ex_reg_valid & ex_ctrl_wxd;
  assign T_7572 = mem_reg_valid & mem_ctrl_wxd;
  assign T_7574 = mem_ctrl_mem == 1'h0;
  assign T_7575 = T_7572 & T_7574;
  assign T_7577 = 5'h0 == ibuf_io_inst_0_bits_inst_rs1;
  assign T_7578 = ex_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_1 = T_7571 & T_7578;
  assign T_7579 = mem_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_2 = T_7575 & T_7579;
  assign id_bypass_src_0_3 = T_7572 & T_7579;
  assign T_7581 = 5'h0 == ibuf_io_inst_0_bits_inst_rs2;
  assign T_7582 = ex_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_1 = T_7571 & T_7582;
  assign T_7583 = mem_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_2 = T_7575 & T_7583;
  assign id_bypass_src_1_3 = T_7572 & T_7583;
  assign bypass_mux_0 = 64'h0;
  assign bypass_mux_1 = mem_reg_wdata;
  assign bypass_mux_2 = wb_reg_wdata;
  assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
  assign T_7612 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign GEN_0 = GEN_4;
  assign GEN_2 = 2'h1 == ex_reg_rs_lsb_0 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_3 = 2'h2 == ex_reg_rs_lsb_0 ? bypass_mux_2 : GEN_2;
  assign GEN_4 = 2'h3 == ex_reg_rs_lsb_0 ? bypass_mux_3 : GEN_3;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? GEN_0 : T_7612;
  assign T_7613 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign GEN_1 = GEN_7;
  assign GEN_5 = 2'h1 == ex_reg_rs_lsb_1 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_6 = 2'h2 == ex_reg_rs_lsb_1 ? bypass_mux_2 : GEN_5;
  assign GEN_7 = 2'h3 == ex_reg_rs_lsb_1 ? bypass_mux_3 : GEN_6;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? GEN_1 : T_7613;
  assign T_7614 = ex_ctrl_sel_imm == 3'h5;
  assign T_7616 = ex_reg_inst[31];
  assign T_7617 = $signed(T_7616);
  assign T_7618 = T_7614 ? $signed(1'sh0) : $signed(T_7617);
  assign T_7619 = ex_ctrl_sel_imm == 3'h2;
  assign T_7620 = ex_reg_inst[30:20];
  assign T_7621 = $signed(T_7620);
  assign T_7622 = T_7619 ? $signed(T_7621) : $signed({11{T_7618}});
  assign T_7623 = ex_ctrl_sel_imm != 3'h2;
  assign T_7624 = ex_ctrl_sel_imm != 3'h3;
  assign T_7625 = T_7623 & T_7624;
  assign T_7626 = ex_reg_inst[19:12];
  assign T_7627 = $signed(T_7626);
  assign T_7628 = T_7625 ? $signed({8{T_7618}}) : $signed(T_7627);
  assign T_7631 = T_7619 | T_7614;
  assign T_7633 = ex_ctrl_sel_imm == 3'h3;
  assign T_7634 = ex_reg_inst[20];
  assign T_7635 = $signed(T_7634);
  assign T_7636 = ex_ctrl_sel_imm == 3'h1;
  assign T_7637 = ex_reg_inst[7];
  assign T_7638 = $signed(T_7637);
  assign T_7639 = T_7636 ? $signed(T_7638) : $signed(T_7618);
  assign T_7640 = T_7633 ? $signed(T_7635) : $signed(T_7639);
  assign T_7641 = T_7631 ? $signed(1'sh0) : $signed(T_7640);
  assign T_7646 = ex_reg_inst[30:25];
  assign T_7647 = T_7631 ? 6'h0 : T_7646;
  assign T_7650 = ex_ctrl_sel_imm == 3'h0;
  assign T_7652 = T_7650 | T_7636;
  assign T_7653 = ex_reg_inst[11:8];
  assign T_7655 = ex_reg_inst[19:16];
  assign T_7656 = ex_reg_inst[24:21];
  assign T_7657 = T_7614 ? T_7655 : T_7656;
  assign T_7658 = T_7652 ? T_7653 : T_7657;
  assign T_7659 = T_7619 ? 4'h0 : T_7658;
  assign T_7662 = ex_ctrl_sel_imm == 3'h4;
  assign T_7665 = ex_reg_inst[15];
  assign T_7668 = T_7614 ? T_7665 : 1'h0;
  assign T_7670 = T_7662 ? T_7634 : T_7668;
  assign T_7672 = T_7650 ? T_7637 : T_7670;
  assign T_7673 = {T_7647,T_7659};
  assign T_7674 = {T_7673,T_7672};
  assign T_7675 = $unsigned(T_7641);
  assign T_7676 = $unsigned(T_7628);
  assign T_7677 = {T_7676,T_7675};
  assign T_7678 = $unsigned(T_7622);
  assign T_7679 = $unsigned(T_7618);
  assign T_7680 = {T_7679,T_7678};
  assign T_7681 = {T_7680,T_7677};
  assign T_7682 = {T_7681,T_7674};
  assign ex_imm = $signed(T_7682);
  assign T_7684 = $signed(ex_rs_0);
  assign T_7685 = $signed(ex_reg_pc);
  assign T_7686 = 2'h2 == ex_ctrl_sel_alu1;
  assign T_7687 = T_7686 ? $signed(T_7685) : $signed(40'sh0);
  assign T_7688 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = T_7688 ? $signed(T_7684) : $signed({{24{T_7687[39]}},T_7687});
  assign T_7690 = $signed(ex_rs_1);
  assign T_7693 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign T_7694 = 2'h1 == ex_ctrl_sel_alu2;
  assign T_7695 = T_7694 ? $signed(T_7693) : $signed(4'sh0);
  assign T_7696 = 2'h3 == ex_ctrl_sel_alu2;
  assign T_7697 = T_7696 ? $signed(ex_imm) : $signed({{28{T_7695[3]}},T_7695});
  assign T_7698 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = T_7698 ? $signed(T_7690) : $signed({{32{T_7697[31]}},T_7697});
  assign alu_clk = clk;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = T_7699;
  assign alu_io_in1 = T_7700;
  assign T_7699 = $unsigned(ex_op2);
  assign T_7700 = $unsigned(ex_op1);
  assign div_clk = clk;
  assign div_reset = reset;
  assign div_io_req_valid = T_7701;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_dw = ex_ctrl_alu_dw;
  assign div_io_req_bits_in1 = ex_rs_0;
  assign div_io_req_bits_in2 = ex_rs_1;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = T_8057;
  assign div_io_resp_ready = GEN_150;
  assign T_7701 = ex_reg_valid & ex_ctrl_div;
  assign T_7703 = ctrl_killd == 1'h0;
  assign T_7705 = take_pc_mem_wb == 1'h0;
  assign T_7706 = T_7705 & ibuf_io_inst_0_valid;
  assign T_7707 = T_7706 & ibuf_io_inst_0_bits_replay;
  assign T_7710 = T_7703 & id_xcpt;
  assign T_7714 = T_7706 & csr_io_interrupt;
  assign GEN_8 = id_xcpt ? id_cause : ex_reg_cause;
  assign GEN_9 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_taken : ex_reg_btb_resp_taken;
  assign GEN_10 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_mask : ex_reg_btb_resp_mask;
  assign GEN_11 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bridx : ex_reg_btb_resp_bridx;
  assign GEN_12 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_target : ex_reg_btb_resp_target;
  assign GEN_13 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_entry : ex_reg_btb_resp_entry;
  assign GEN_14 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bht_history : ex_reg_btb_resp_bht_history;
  assign GEN_15 = ibuf_io_inst_0_bits_btb_hit ? ibuf_io_btb_resp_bht_value : ex_reg_btb_resp_bht_value;
  assign T_7718 = bpu_io_xcpt_if == 1'h0;
  assign T_7720 = ibuf_io_inst_0_bits_pf0 == 1'h0;
  assign T_7721 = T_7718 & T_7720;
  assign T_7722 = T_7721 & ibuf_io_inst_0_bits_pf1;
  assign GEN_16 = T_7722 ? 2'h1 : 2'h0;
  assign GEN_17 = T_7722 ? 1'h1 : ibuf_io_inst_0_bits_rvc;
  assign GEN_18 = id_xcpt ? 4'h0 : id_ctrl_alu_fn;
  assign GEN_19 = id_xcpt ? 1'h1 : id_ctrl_alu_dw;
  assign GEN_20 = id_xcpt ? 2'h2 : id_ctrl_sel_alu1;
  assign GEN_21 = id_xcpt ? GEN_16 : id_ctrl_sel_alu2;
  assign GEN_22 = id_xcpt ? GEN_17 : ibuf_io_inst_0_bits_rvc;
  assign T_7724 = id_ctrl_fence_i | id_csr_flush;
  assign T_7725 = T_7724 | csr_io_singleStep;
  assign T_7726 = id_ctrl_jalr & csr_io_status_debug;
  assign GEN_23 = T_7726 ? 1'h1 : T_7725;
  assign GEN_24 = T_7726 ? 1'h1 : id_ctrl_fence_i;
  assign T_7729 = T_7577 | id_bypass_src_0_1;
  assign T_7730 = T_7729 | id_bypass_src_0_2;
  assign T_7731 = T_7730 | id_bypass_src_0_3;
  assign T_7736 = id_bypass_src_0_2 ? 2'h2 : 2'h3;
  assign T_7737 = id_bypass_src_0_1 ? 2'h1 : T_7736;
  assign T_7738 = T_7577 ? 2'h0 : T_7737;
  assign T_7740 = T_7731 == 1'h0;
  assign T_7741 = id_ctrl_rxs1 & T_7740;
  assign T_7742 = id_rs_0[1:0];
  assign T_7743 = id_rs_0[63:2];
  assign GEN_25 = T_7741 ? T_7742 : T_7738;
  assign GEN_26 = T_7741 ? T_7743 : ex_reg_rs_msb_0;
  assign T_7744 = T_7581 | id_bypass_src_1_1;
  assign T_7745 = T_7744 | id_bypass_src_1_2;
  assign T_7746 = T_7745 | id_bypass_src_1_3;
  assign T_7751 = id_bypass_src_1_2 ? 2'h2 : 2'h3;
  assign T_7752 = id_bypass_src_1_1 ? 2'h1 : T_7751;
  assign T_7753 = T_7581 ? 2'h0 : T_7752;
  assign T_7755 = T_7746 == 1'h0;
  assign T_7756 = id_ctrl_rxs2 & T_7755;
  assign T_7757 = id_rs_1[1:0];
  assign T_7758 = id_rs_1[63:2];
  assign GEN_27 = T_7756 ? T_7757 : T_7753;
  assign GEN_28 = T_7756 ? T_7758 : ex_reg_rs_msb_1;
  assign GEN_29 = T_7703 ? id_ctrl_legal : ex_ctrl_legal;
  assign GEN_30 = T_7703 ? id_ctrl_fp : ex_ctrl_fp;
  assign GEN_31 = T_7703 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign GEN_32 = T_7703 ? id_ctrl_branch : ex_ctrl_branch;
  assign GEN_33 = T_7703 ? id_ctrl_jal : ex_ctrl_jal;
  assign GEN_34 = T_7703 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign GEN_35 = T_7703 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign GEN_36 = T_7703 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign GEN_37 = T_7703 ? GEN_21 : ex_ctrl_sel_alu2;
  assign GEN_38 = T_7703 ? GEN_20 : ex_ctrl_sel_alu1;
  assign GEN_39 = T_7703 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign GEN_40 = T_7703 ? GEN_19 : ex_ctrl_alu_dw;
  assign GEN_41 = T_7703 ? GEN_18 : ex_ctrl_alu_fn;
  assign GEN_42 = T_7703 ? id_ctrl_mem : ex_ctrl_mem;
  assign GEN_43 = T_7703 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign GEN_44 = T_7703 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign GEN_45 = T_7703 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign GEN_46 = T_7703 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign GEN_47 = T_7703 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign GEN_48 = T_7703 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign GEN_49 = T_7703 ? id_ctrl_div : ex_ctrl_div;
  assign GEN_50 = T_7703 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign GEN_51 = T_7703 ? id_csr : ex_ctrl_csr;
  assign GEN_52 = T_7703 ? GEN_24 : ex_ctrl_fence_i;
  assign GEN_53 = T_7703 ? id_ctrl_fence : ex_ctrl_fence;
  assign GEN_54 = T_7703 ? id_ctrl_amo : ex_ctrl_amo;
  assign GEN_55 = T_7703 ? GEN_22 : ex_reg_rvc;
  assign GEN_56 = T_7703 ? GEN_23 : ex_reg_flush_pipe;
  assign GEN_57 = T_7703 ? id_load_use : ex_reg_load_use;
  assign GEN_58 = T_7703 ? T_7731 : ex_reg_rs_bypass_0;
  assign GEN_59 = T_7703 ? GEN_25 : ex_reg_rs_lsb_0;
  assign GEN_60 = T_7703 ? GEN_26 : ex_reg_rs_msb_0;
  assign GEN_61 = T_7703 ? T_7746 : ex_reg_rs_bypass_1;
  assign GEN_62 = T_7703 ? GEN_27 : ex_reg_rs_lsb_1;
  assign GEN_63 = T_7703 ? GEN_28 : ex_reg_rs_msb_1;
  assign T_7761 = T_7703 | csr_io_interrupt;
  assign T_7762 = T_7761 | ibuf_io_inst_0_bits_replay;
  assign GEN_64 = T_7762 ? ibuf_io_inst_0_bits_inst_bits : ex_reg_inst;
  assign GEN_65 = T_7762 ? ibuf_io_pc : ex_reg_pc;
  assign T_7763 = ex_reg_valid | ex_reg_replay;
  assign ex_pc_valid = T_7763 | ex_reg_xcpt_interrupt;
  assign T_7765 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & T_7765;
  assign T_7767 = io_dmem_req_ready == 1'h0;
  assign T_7768 = ex_ctrl_mem & T_7767;
  assign T_7770 = div_io_req_ready == 1'h0;
  assign T_7771 = ex_ctrl_div & T_7770;
  assign replay_ex_structural = T_7768 | T_7771;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T_7772 = replay_ex_structural | replay_ex_load_use;
  assign T_7773 = ex_reg_valid & T_7772;
  assign replay_ex = ex_reg_replay | T_7773;
  assign T_7774 = take_pc_mem_wb | replay_ex;
  assign T_7776 = ex_reg_valid == 1'h0;
  assign ctrl_killx = T_7774 | T_7776;
  assign T_7777 = ex_ctrl_mem_cmd == 5'h7;
  assign T_7783_0 = 3'h0;
  assign T_7783_1 = 3'h4;
  assign T_7783_2 = 3'h1;
  assign T_7783_3 = 3'h5;
  assign T_7785 = T_7783_0 == ex_ctrl_mem_type;
  assign T_7786 = T_7783_1 == ex_ctrl_mem_type;
  assign T_7787 = T_7783_2 == ex_ctrl_mem_type;
  assign T_7788 = T_7783_3 == ex_ctrl_mem_type;
  assign T_7791 = T_7785 | T_7786;
  assign T_7792 = T_7791 | T_7787;
  assign T_7793 = T_7792 | T_7788;
  assign ex_slow_bypass = T_7777 | T_7793;
  assign T_7794 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T_7795 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign ex_xcpt = T_7794 | T_7795;
  assign ex_cause = T_7794 ? ex_reg_cause : 64'h2;
  assign mem_br_taken = mem_reg_wdata[0];
  assign T_7797 = $signed(mem_reg_pc);
  assign T_7798 = mem_ctrl_branch & mem_br_taken;
  assign T_7801 = mem_reg_inst[31];
  assign T_7802 = $signed(T_7801);
  assign T_7807 = {11{T_7802}};
  assign T_7811 = mem_reg_inst[19:12];
  assign T_7812 = $signed(T_7811);
  assign T_7813 = {8{T_7802}};
  assign T_7819 = mem_reg_inst[20];
  assign T_7820 = $signed(T_7819);
  assign T_7822 = mem_reg_inst[7];
  assign T_7823 = $signed(T_7822);
  assign T_7831 = mem_reg_inst[30:25];
  assign T_7838 = mem_reg_inst[11:8];
  assign T_7841 = mem_reg_inst[24:21];
  assign T_7858 = {T_7831,T_7838};
  assign T_7859 = {T_7858,1'h0};
  assign T_7860 = $unsigned(T_7823);
  assign T_7861 = $unsigned(T_7813);
  assign T_7862 = {T_7861,T_7860};
  assign T_7863 = $unsigned(T_7807);
  assign T_7864 = $unsigned(T_7802);
  assign T_7865 = {T_7864,T_7863};
  assign T_7866 = {T_7865,T_7862};
  assign T_7867 = {T_7866,T_7859};
  assign T_7868 = $signed(T_7867);
  assign T_7928 = {T_7831,T_7841};
  assign T_7929 = {T_7928,1'h0};
  assign T_7930 = $unsigned(T_7820);
  assign T_7931 = $unsigned(T_7812);
  assign T_7932 = {T_7931,T_7930};
  assign T_7936 = {T_7865,T_7932};
  assign T_7937 = {T_7936,T_7929};
  assign T_7938 = $signed(T_7937);
  assign T_7941 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign T_7942 = mem_ctrl_jal ? $signed(T_7938) : $signed({{28{T_7941[3]}},T_7941});
  assign T_7943 = T_7798 ? $signed(T_7868) : $signed(T_7942);
  assign GEN_174 = {{8{T_7943[31]}},T_7943};
  assign T_7944 = $signed(T_7797) + $signed(GEN_174);
  assign T_7945 = T_7944[39:0];
  assign mem_br_target = $signed(T_7945);
  assign T_7946 = mem_reg_wdata[63:38];
  assign T_7947 = mem_reg_wdata[39:38];
  assign T_7948 = $signed(T_7947);
  assign T_7950 = T_7946 == 26'h0;
  assign T_7952 = T_7946 == 26'h1;
  assign T_7953 = T_7950 | T_7952;
  assign T_7955 = $signed(T_7948) != $signed(2'sh0);
  assign T_7956 = $signed(T_7946);
  assign T_7958 = $signed(T_7956) == $signed(26'sh3ffffff);
  assign T_7961 = $signed(T_7956) == $signed(26'sh3fffffe);
  assign T_7962 = T_7958 | T_7961;
  assign T_7964 = $signed(T_7948) == $signed(2'sh3);
  assign T_7965 = T_7948[0];
  assign T_7966 = T_7962 ? T_7964 : T_7965;
  assign T_7967 = T_7953 ? T_7955 : T_7966;
  assign T_7968 = mem_reg_wdata[38:0];
  assign T_7969 = {T_7967,T_7968};
  assign T_7970 = $signed(T_7969);
  assign T_7971 = mem_ctrl_jalr ? $signed(T_7970) : $signed(mem_br_target);
  assign T_7973 = $signed(T_7971) & $signed(40'shfffffffffe);
  assign T_7974 = $signed(T_7973);
  assign mem_npc = $unsigned(T_7974);
  assign T_7975 = mem_npc != ex_reg_pc;
  assign T_7976 = mem_npc != ibuf_io_pc;
  assign T_7978 = ibuf_io_inst_0_valid ? T_7976 : 1'h1;
  assign mem_wrong_npc = ex_pc_valid ? T_7975 : T_7978;
  assign T_7980 = mem_reg_xcpt == 1'h0;
  assign T_7982 = T_7980 & mem_ctrl_jalr;
  assign T_7983 = $signed(mem_reg_wdata);
  assign T_7984 = T_7982 ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(T_7983);
  assign mem_int_wdata = $unsigned(T_7984);
  assign T_7985 = mem_ctrl_branch | mem_ctrl_jalr;
  assign mem_cfi = T_7985 | mem_ctrl_jal;
  assign T_7987 = T_7798 | mem_ctrl_jalr;
  assign mem_cfi_taken = T_7987 | mem_ctrl_jal;
  assign T_7988 = mem_wrong_npc | mem_reg_flush_pipe;
  assign T_7989 = mem_reg_valid & T_7988;
  assign T_7991 = ctrl_killx == 1'h0;
  assign T_7994 = T_7705 & replay_ex;
  assign T_7997 = T_7991 & ex_xcpt;
  assign T_8000 = T_7705 & ex_reg_xcpt_interrupt;
  assign GEN_66 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign T_8001 = ex_ctrl_mem_cmd == 5'h0;
  assign T_8002 = ex_ctrl_mem_cmd == 5'h6;
  assign T_8003 = T_8001 | T_8002;
  assign T_8005 = T_8003 | T_7777;
  assign T_8006 = ex_ctrl_mem_cmd[3];
  assign T_8007 = ex_ctrl_mem_cmd == 5'h4;
  assign T_8008 = T_8006 | T_8007;
  assign T_8009 = T_8005 | T_8008;
  assign T_8010 = ex_ctrl_mem & T_8009;
  assign T_8011 = ex_ctrl_mem_cmd == 5'h1;
  assign T_8013 = T_8011 | T_7777;
  assign T_8017 = T_8013 | T_8008;
  assign T_8018 = ex_ctrl_mem & T_8017;
  assign GEN_67 = ex_reg_btb_hit ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign GEN_68 = ex_reg_btb_hit ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign GEN_69 = ex_reg_btb_hit ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign GEN_70 = ex_reg_btb_hit ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign GEN_71 = ex_reg_btb_hit ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign GEN_72 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign GEN_73 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T_8019 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T_8020 = ex_ctrl_rxs2 & T_8019;
  assign GEN_74 = T_8020 ? ex_rs_1 : mem_reg_rs2;
  assign GEN_75 = ex_pc_valid ? ex_ctrl_legal : mem_ctrl_legal;
  assign GEN_76 = ex_pc_valid ? ex_ctrl_fp : mem_ctrl_fp;
  assign GEN_77 = ex_pc_valid ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign GEN_78 = ex_pc_valid ? ex_ctrl_branch : mem_ctrl_branch;
  assign GEN_79 = ex_pc_valid ? ex_ctrl_jal : mem_ctrl_jal;
  assign GEN_80 = ex_pc_valid ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign GEN_81 = ex_pc_valid ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign GEN_82 = ex_pc_valid ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign GEN_83 = ex_pc_valid ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign GEN_84 = ex_pc_valid ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign GEN_85 = ex_pc_valid ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign GEN_86 = ex_pc_valid ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign GEN_87 = ex_pc_valid ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign GEN_88 = ex_pc_valid ? ex_ctrl_mem : mem_ctrl_mem;
  assign GEN_89 = ex_pc_valid ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign GEN_90 = ex_pc_valid ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign GEN_91 = ex_pc_valid ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign GEN_92 = ex_pc_valid ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign GEN_93 = ex_pc_valid ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign GEN_94 = ex_pc_valid ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign GEN_95 = ex_pc_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_96 = ex_pc_valid ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign GEN_97 = ex_pc_valid ? ex_ctrl_csr : mem_ctrl_csr;
  assign GEN_98 = ex_pc_valid ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign GEN_99 = ex_pc_valid ? ex_ctrl_fence : mem_ctrl_fence;
  assign GEN_100 = ex_pc_valid ? ex_ctrl_amo : mem_ctrl_amo;
  assign GEN_101 = ex_pc_valid ? ex_reg_rvc : mem_reg_rvc;
  assign GEN_102 = ex_pc_valid ? T_8010 : mem_reg_load;
  assign GEN_103 = ex_pc_valid ? T_8018 : mem_reg_store;
  assign GEN_104 = ex_pc_valid ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign GEN_105 = ex_pc_valid ? GEN_67 : mem_reg_btb_resp_taken;
  assign GEN_106 = ex_pc_valid ? GEN_68 : mem_reg_btb_resp_mask;
  assign GEN_107 = ex_pc_valid ? GEN_69 : mem_reg_btb_resp_bridx;
  assign GEN_108 = ex_pc_valid ? GEN_70 : mem_reg_btb_resp_target;
  assign GEN_109 = ex_pc_valid ? GEN_71 : mem_reg_btb_resp_entry;
  assign GEN_110 = ex_pc_valid ? GEN_72 : mem_reg_btb_resp_bht_history;
  assign GEN_111 = ex_pc_valid ? GEN_73 : mem_reg_btb_resp_bht_value;
  assign GEN_112 = ex_pc_valid ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign GEN_113 = ex_pc_valid ? ex_slow_bypass : mem_reg_slow_bypass;
  assign GEN_114 = ex_pc_valid ? ex_reg_inst : mem_reg_inst;
  assign GEN_115 = ex_pc_valid ? ex_reg_pc : mem_reg_pc;
  assign GEN_116 = ex_pc_valid ? alu_io_out : mem_reg_wdata;
  assign GEN_117 = ex_pc_valid ? GEN_74 : mem_reg_rs2;
  assign T_8021 = mem_reg_load & bpu_io_xcpt_ld;
  assign T_8022 = mem_reg_store & bpu_io_xcpt_st;
  assign mem_breakpoint = T_8021 | T_8022;
  assign T_8023 = mem_reg_load & bpu_io_debug_ld;
  assign T_8024 = mem_reg_store & bpu_io_debug_st;
  assign mem_debug_breakpoint = T_8023 | T_8024;
  assign T_8028 = mem_ctrl_mem & io_dmem_xcpt_ma_st;
  assign T_8030 = mem_ctrl_mem & io_dmem_xcpt_ma_ld;
  assign T_8032 = mem_ctrl_mem & io_dmem_xcpt_pf_st;
  assign T_8034 = mem_ctrl_mem & io_dmem_xcpt_pf_ld;
  assign T_8036 = mem_debug_breakpoint | mem_breakpoint;
  assign T_8038 = T_8036 | T_8028;
  assign T_8039 = T_8038 | T_8030;
  assign T_8040 = T_8039 | T_8032;
  assign mem_new_xcpt = T_8040 | T_8034;
  assign T_8041 = T_8032 ? 3'h7 : 3'h5;
  assign T_8042 = T_8030 ? 3'h4 : T_8041;
  assign T_8043 = T_8028 ? 3'h6 : T_8042;
  assign T_8045 = mem_breakpoint ? 3'h3 : T_8043;
  assign mem_new_cause = mem_debug_breakpoint ? 4'hd : {{1'd0}, T_8045};
  assign T_8046 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T_8047 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = T_8046 | T_8047;
  assign mem_cause = T_8046 ? mem_reg_cause : {{60'd0}, mem_new_cause};
  assign dcache_kill_mem = T_7572 & io_dmem_replay_next;
  assign T_8049 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = T_8049 & io_fpu_nack_mem;
  assign T_8050 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = T_8050 | fpu_kill_mem;
  assign T_8051 = dcache_kill_mem | take_pc_wb;
  assign T_8052 = T_8051 | mem_reg_xcpt;
  assign T_8054 = mem_reg_valid == 1'h0;
  assign killm_common = T_8052 | T_8054;
  assign T_8055 = div_io_req_ready & div_io_req_valid;
  assign T_8057 = killm_common & T_8056;
  assign T_8058 = killm_common | mem_xcpt;
  assign ctrl_killm = T_8058 | fpu_kill_mem;
  assign T_8060 = ctrl_killm == 1'h0;
  assign T_8062 = take_pc_wb == 1'h0;
  assign T_8063 = replay_mem & T_8062;
  assign T_8066 = mem_xcpt & T_8062;
  assign GEN_118 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign T_8067 = mem_reg_valid | mem_reg_replay;
  assign T_8068 = T_8067 | mem_reg_xcpt_interrupt;
  assign T_8071 = T_7980 & mem_ctrl_fp;
  assign T_8072 = T_8071 & mem_ctrl_wxd;
  assign T_8073 = T_8072 ? io_fpu_toint_data : mem_int_wdata;
  assign GEN_119 = mem_ctrl_rocc ? mem_reg_rs2 : wb_reg_rs2;
  assign GEN_120 = T_8068 ? mem_ctrl_legal : wb_ctrl_legal;
  assign GEN_121 = T_8068 ? mem_ctrl_fp : wb_ctrl_fp;
  assign GEN_122 = T_8068 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign GEN_123 = T_8068 ? mem_ctrl_branch : wb_ctrl_branch;
  assign GEN_124 = T_8068 ? mem_ctrl_jal : wb_ctrl_jal;
  assign GEN_125 = T_8068 ? mem_ctrl_jalr : wb_ctrl_jalr;
  assign GEN_126 = T_8068 ? mem_ctrl_rxs2 : wb_ctrl_rxs2;
  assign GEN_127 = T_8068 ? mem_ctrl_rxs1 : wb_ctrl_rxs1;
  assign GEN_128 = T_8068 ? mem_ctrl_sel_alu2 : wb_ctrl_sel_alu2;
  assign GEN_129 = T_8068 ? mem_ctrl_sel_alu1 : wb_ctrl_sel_alu1;
  assign GEN_130 = T_8068 ? mem_ctrl_sel_imm : wb_ctrl_sel_imm;
  assign GEN_131 = T_8068 ? mem_ctrl_alu_dw : wb_ctrl_alu_dw;
  assign GEN_132 = T_8068 ? mem_ctrl_alu_fn : wb_ctrl_alu_fn;
  assign GEN_133 = T_8068 ? mem_ctrl_mem : wb_ctrl_mem;
  assign GEN_134 = T_8068 ? mem_ctrl_mem_cmd : wb_ctrl_mem_cmd;
  assign GEN_135 = T_8068 ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign GEN_136 = T_8068 ? mem_ctrl_rfs1 : wb_ctrl_rfs1;
  assign GEN_137 = T_8068 ? mem_ctrl_rfs2 : wb_ctrl_rfs2;
  assign GEN_138 = T_8068 ? mem_ctrl_rfs3 : wb_ctrl_rfs3;
  assign GEN_139 = T_8068 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign GEN_140 = T_8068 ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_141 = T_8068 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign GEN_142 = T_8068 ? mem_ctrl_csr : wb_ctrl_csr;
  assign GEN_143 = T_8068 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign GEN_144 = T_8068 ? mem_ctrl_fence : wb_ctrl_fence;
  assign GEN_145 = T_8068 ? mem_ctrl_amo : wb_ctrl_amo;
  assign GEN_146 = T_8068 ? T_8073 : wb_reg_wdata;
  assign GEN_147 = T_8068 ? GEN_119 : wb_reg_rs2;
  assign GEN_148 = T_8068 ? mem_reg_inst : wb_reg_inst;
  assign GEN_149 = T_8068 ? mem_reg_pc : wb_reg_pc;
  assign T_8074 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = T_8074 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign T_8077 = io_rocc_cmd_ready == 1'h0;
  assign replay_wb_rocc = T_7546 & T_8077;
  assign replay_wb = replay_wb_common | replay_wb_rocc;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T_8078 = replay_wb | wb_xcpt;
  assign T_8079 = T_8078 | csr_io_eret;
  assign T_8080 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = T_8080 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign T_8084 = wb_reg_valid & wb_ctrl_wxd;
  assign T_8086 = T_8084 == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign ll_waddr = GEN_151;
  assign T_8087 = div_io_resp_ready & div_io_resp_valid;
  assign ll_wen = GEN_152;
  assign T_8088 = dmem_resp_replay & dmem_resp_xpu;
  assign GEN_150 = T_8088 ? 1'h0 : T_8086;
  assign GEN_151 = T_8088 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign GEN_152 = T_8088 ? 1'h1 : T_8087;
  assign T_8092 = replay_wb == 1'h0;
  assign T_8093 = wb_reg_valid & T_8092;
  assign T_8095 = wb_xcpt == 1'h0;
  assign wb_valid = T_8093 & T_8095;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | ll_wen;
  assign rf_waddr = ll_wen ? ll_waddr : wb_waddr;
  assign T_8096 = dmem_resp_valid & dmem_resp_xpu;
  assign T_8097 = wb_ctrl_csr != 3'h0;
  assign T_8098 = T_8097 ? csr_io_rw_rdata : wb_reg_wdata;
  assign T_8099 = ll_wen ? ll_wdata : T_8098;
  assign rf_wdata = T_8096 ? io_dmem_resp_bits_data : T_8099;
  assign T_8101 = rf_waddr != 5'h0;
  assign T_8103 = ~ rf_waddr;
  assign T_8105 = rf_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign GEN_153 = T_8105 ? rf_wdata : T_7362;
  assign T_8106 = rf_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign GEN_154 = T_8106 ? rf_wdata : T_7372;
  assign GEN_160 = T_8101 ? GEN_153 : T_7362;
  assign GEN_161 = T_8101 ? GEN_154 : T_7372;
  assign GEN_164 = rf_wen ? T_8101 : 1'h0;
  assign GEN_167 = rf_wen ? GEN_160 : T_7362;
  assign GEN_168 = rf_wen ? GEN_161 : T_7372;
  assign T_8107 = wb_reg_wdata[63:38];
  assign T_8108 = wb_reg_wdata[39:38];
  assign T_8109 = $signed(T_8108);
  assign T_8111 = T_8107 == 26'h0;
  assign T_8113 = T_8107 == 26'h1;
  assign T_8114 = T_8111 | T_8113;
  assign T_8116 = $signed(T_8109) != $signed(2'sh0);
  assign T_8117 = $signed(T_8107);
  assign T_8119 = $signed(T_8117) == $signed(26'sh3ffffff);
  assign T_8122 = $signed(T_8117) == $signed(26'sh3fffffe);
  assign T_8123 = T_8119 | T_8122;
  assign T_8125 = $signed(T_8109) == $signed(2'sh3);
  assign T_8126 = T_8109[0];
  assign T_8127 = T_8123 ? T_8125 : T_8126;
  assign T_8128 = T_8114 ? T_8116 : T_8127;
  assign T_8129 = wb_reg_wdata[38:0];
  assign T_8130 = {T_8128,T_8129};
  assign T_8131 = wb_reg_inst[31:20];
  assign T_8132 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T_8134 = ibuf_io_inst_0_bits_inst_rs1 != 5'h0;
  assign T_8135 = id_ctrl_rxs1 & T_8134;
  assign T_8137 = ibuf_io_inst_0_bits_inst_rs2 != 5'h0;
  assign T_8138 = id_ctrl_rxs2 & T_8137;
  assign T_8140 = ibuf_io_inst_0_bits_inst_rd != 5'h0;
  assign T_8141 = id_ctrl_wxd & T_8140;
  assign T_8144 = T_8143[31:1];
  assign GEN_175 = {{1'd0}, T_8144};
  assign T_8145 = GEN_175 << 1;
  assign T_8148 = 32'h1 << ll_waddr;
  assign T_8150 = ll_wen ? T_8148 : 32'h0;
  assign T_8151 = ~ T_8150;
  assign T_8152 = T_8145 & T_8151;
  assign GEN_169 = ll_wen ? T_8152 : T_8143;
  assign T_8154 = T_8145 >> ibuf_io_inst_0_bits_inst_rs1;
  assign T_8155 = T_8154[0];
  assign T_8156 = T_8135 & T_8155;
  assign T_8157 = T_8145 >> ibuf_io_inst_0_bits_inst_rs2;
  assign T_8158 = T_8157[0];
  assign T_8159 = T_8138 & T_8158;
  assign T_8160 = T_8145 >> ibuf_io_inst_0_bits_inst_rd;
  assign T_8161 = T_8160[0];
  assign T_8162 = T_8141 & T_8161;
  assign T_8163 = T_8156 | T_8159;
  assign id_sboard_hazard = T_8163 | T_8162;
  assign T_8164 = wb_set_sboard & wb_wen;
  assign T_8166 = 32'h1 << wb_waddr;
  assign T_8168 = T_8164 ? T_8166 : 32'h0;
  assign T_8169 = T_8152 | T_8168;
  assign T_8170 = ll_wen | T_8164;
  assign GEN_170 = T_8170 ? T_8169 : GEN_169;
  assign T_8171 = ex_ctrl_csr != 3'h0;
  assign T_8172 = T_8171 | ex_ctrl_jalr;
  assign T_8173 = T_8172 | ex_ctrl_mem;
  assign T_8174 = T_8173 | ex_ctrl_div;
  assign T_8175 = T_8174 | ex_ctrl_fp;
  assign ex_cannot_bypass = T_8175 | ex_ctrl_rocc;
  assign T_8176 = ibuf_io_inst_0_bits_inst_rs1 == ex_waddr;
  assign T_8177 = T_8135 & T_8176;
  assign T_8178 = ibuf_io_inst_0_bits_inst_rs2 == ex_waddr;
  assign T_8179 = T_8138 & T_8178;
  assign T_8180 = ibuf_io_inst_0_bits_inst_rd == ex_waddr;
  assign T_8181 = T_8141 & T_8180;
  assign T_8182 = T_8177 | T_8179;
  assign T_8183 = T_8182 | T_8181;
  assign data_hazard_ex = ex_ctrl_wxd & T_8183;
  assign T_8185 = io_fpu_dec_ren1 & T_8176;
  assign T_8187 = io_fpu_dec_ren2 & T_8178;
  assign T_8188 = ibuf_io_inst_0_bits_inst_rs3 == ex_waddr;
  assign T_8189 = io_fpu_dec_ren3 & T_8188;
  assign T_8191 = io_fpu_dec_wen & T_8180;
  assign T_8192 = T_8185 | T_8187;
  assign T_8193 = T_8192 | T_8189;
  assign T_8194 = T_8193 | T_8191;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T_8194;
  assign T_8195 = data_hazard_ex & ex_cannot_bypass;
  assign T_8196 = T_8195 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & T_8196;
  assign T_8198 = mem_ctrl_csr != 3'h0;
  assign T_8199 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign T_8200 = T_8198 | T_8199;
  assign T_8201 = T_8200 | mem_ctrl_div;
  assign T_8202 = T_8201 | mem_ctrl_fp;
  assign mem_cannot_bypass = T_8202 | mem_ctrl_rocc;
  assign T_8203 = ibuf_io_inst_0_bits_inst_rs1 == mem_waddr;
  assign T_8204 = T_8135 & T_8203;
  assign T_8205 = ibuf_io_inst_0_bits_inst_rs2 == mem_waddr;
  assign T_8206 = T_8138 & T_8205;
  assign T_8207 = ibuf_io_inst_0_bits_inst_rd == mem_waddr;
  assign T_8208 = T_8141 & T_8207;
  assign T_8209 = T_8204 | T_8206;
  assign T_8210 = T_8209 | T_8208;
  assign data_hazard_mem = mem_ctrl_wxd & T_8210;
  assign T_8212 = io_fpu_dec_ren1 & T_8203;
  assign T_8214 = io_fpu_dec_ren2 & T_8205;
  assign T_8215 = ibuf_io_inst_0_bits_inst_rs3 == mem_waddr;
  assign T_8216 = io_fpu_dec_ren3 & T_8215;
  assign T_8218 = io_fpu_dec_wen & T_8207;
  assign T_8219 = T_8212 | T_8214;
  assign T_8220 = T_8219 | T_8216;
  assign T_8221 = T_8220 | T_8218;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T_8221;
  assign T_8222 = data_hazard_mem & mem_cannot_bypass;
  assign T_8223 = T_8222 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & T_8223;
  assign T_8224 = mem_reg_valid & data_hazard_mem;
  assign T_8225 = T_8224 & mem_ctrl_mem;
  assign T_8226 = ibuf_io_inst_0_bits_inst_rs1 == wb_waddr;
  assign T_8227 = T_8135 & T_8226;
  assign T_8228 = ibuf_io_inst_0_bits_inst_rs2 == wb_waddr;
  assign T_8229 = T_8138 & T_8228;
  assign T_8230 = ibuf_io_inst_0_bits_inst_rd == wb_waddr;
  assign T_8231 = T_8141 & T_8230;
  assign T_8232 = T_8227 | T_8229;
  assign T_8233 = T_8232 | T_8231;
  assign data_hazard_wb = wb_ctrl_wxd & T_8233;
  assign T_8235 = io_fpu_dec_ren1 & T_8226;
  assign T_8237 = io_fpu_dec_ren2 & T_8228;
  assign T_8238 = ibuf_io_inst_0_bits_inst_rs3 == wb_waddr;
  assign T_8239 = io_fpu_dec_ren3 & T_8238;
  assign T_8241 = io_fpu_dec_wen & T_8230;
  assign T_8242 = T_8235 | T_8237;
  assign T_8243 = T_8242 | T_8239;
  assign T_8244 = T_8243 | T_8241;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T_8244;
  assign T_8245 = data_hazard_wb & wb_set_sboard;
  assign T_8246 = T_8245 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & T_8246;
  assign T_8250 = wb_dcache_miss & wb_ctrl_wfd;
  assign T_8251 = T_8250 | io_fpu_sboard_set;
  assign T_8252 = T_8251 & wb_valid;
  assign T_8256 = T_8252 ? T_8166 : 32'h0;
  assign T_8257 = T_8248 | T_8256;
  assign GEN_171 = T_8252 ? T_8257 : T_8248;
  assign T_8259 = dmem_resp_replay & T_8080;
  assign T_8261 = 32'h1 << dmem_resp_waddr;
  assign T_8263 = T_8259 ? T_8261 : 32'h0;
  assign T_8264 = ~ T_8263;
  assign T_8265 = T_8257 & T_8264;
  assign T_8266 = T_8252 | T_8259;
  assign GEN_172 = T_8266 ? T_8265 : GEN_171;
  assign T_8268 = 32'h1 << io_fpu_sboard_clra;
  assign T_8270 = io_fpu_sboard_clr ? T_8268 : 32'h0;
  assign T_8271 = ~ T_8270;
  assign T_8272 = T_8265 & T_8271;
  assign T_8273 = T_8266 | io_fpu_sboard_clr;
  assign GEN_173 = T_8273 ? T_8272 : GEN_172;
  assign T_8275 = io_fpu_fcsr_rdy == 1'h0;
  assign T_8276 = id_csr_en & T_8275;
  assign T_8277 = T_8248 >> ibuf_io_inst_0_bits_inst_rs1;
  assign T_8278 = T_8277[0];
  assign T_8279 = io_fpu_dec_ren1 & T_8278;
  assign T_8280 = T_8248 >> ibuf_io_inst_0_bits_inst_rs2;
  assign T_8281 = T_8280[0];
  assign T_8282 = io_fpu_dec_ren2 & T_8281;
  assign T_8283 = T_8248 >> ibuf_io_inst_0_bits_inst_rs3;
  assign T_8284 = T_8283[0];
  assign T_8285 = io_fpu_dec_ren3 & T_8284;
  assign T_8286 = T_8248 >> ibuf_io_inst_0_bits_inst_rd;
  assign T_8287 = T_8286[0];
  assign T_8288 = io_fpu_dec_wen & T_8287;
  assign T_8289 = T_8279 | T_8282;
  assign T_8290 = T_8289 | T_8285;
  assign T_8291 = T_8290 | T_8288;
  assign id_stall_fpu = T_8276 | T_8291;
  assign T_8295 = io_dmem_req_valid | dcache_blocked;
  assign T_8296 = T_7767 & T_8295;
  assign T_8299 = wb_reg_xcpt == 1'h0;
  assign T_8302 = T_8299 & T_8077;
  assign T_8303 = io_rocc_cmd_valid | rocc_blocked;
  assign T_8304 = T_8302 & T_8303;
  assign T_8305 = id_ex_hazard | id_mem_hazard;
  assign T_8306 = T_8305 | id_wb_hazard;
  assign T_8307 = T_8306 | id_sboard_hazard;
  assign T_8308 = id_ctrl_fp & id_stall_fpu;
  assign T_8309 = T_8307 | T_8308;
  assign T_8310 = id_ctrl_mem & dcache_blocked;
  assign T_8311 = T_8309 | T_8310;
  assign T_8312 = id_ctrl_rocc & rocc_blocked;
  assign T_8313 = T_8311 | T_8312;
  assign T_8314 = T_8313 | T_7557;
  assign ctrl_stalld = T_8314 | csr_io_csr_stall;
  assign T_8316 = ibuf_io_inst_0_valid == 1'h0;
  assign T_8317 = T_8316 | ibuf_io_inst_0_bits_replay;
  assign T_8318 = T_8317 | take_pc_mem_wb;
  assign T_8319 = T_8318 | ctrl_stalld;
  assign T_8320 = T_8319 | csr_io_interrupt;
  assign T_8323 = wb_xcpt | csr_io_eret;
  assign T_8324 = replay_wb ? wb_reg_pc : mem_npc;
  assign T_8325 = T_8323 ? csr_io_evec : T_8324;
  assign T_8326 = wb_reg_valid & wb_ctrl_fence_i;
  assign T_8328 = io_dmem_s2_nack == 1'h0;
  assign T_8329 = T_8326 & T_8328;
  assign T_8331 = ctrl_stalld == 1'h0;
  assign T_8332 = T_8331 | csr_io_interrupt;
  assign T_8333 = mem_reg_replay & mem_reg_btb_hit;
  assign T_8336 = mem_reg_valid & T_8062;
  assign T_8338 = mem_cfi == 1'h0;
  assign T_8339 = mem_cfi_taken | T_8338;
  assign T_8340 = T_8336 & T_8339;
  assign T_8341 = T_8340 & mem_wrong_npc;
  assign T_8342 = T_8333 | T_8341;
  assign T_8344 = mem_reg_replay == 1'h0;
  assign T_8345 = T_8344 & mem_cfi;
  assign T_8346 = mem_ctrl_jal | mem_ctrl_jalr;
  assign T_8347 = mem_reg_inst[19:15];
  assign T_8350 = T_8347 & 5'h19;
  assign T_8351 = 5'h1 == T_8350;
  assign T_8352 = mem_ctrl_jalr & T_8351;
  assign T_8355 = mem_reg_rvc ? 2'h0 : 2'h2;
  assign GEN_176 = {{38'd0}, T_8355};
  assign T_8356 = mem_reg_pc + GEN_176;
  assign T_8357 = T_8356[39:0];
  assign T_8358 = ~ io_imem_btb_update_bits_br_pc;
  assign T_8360 = T_8358 | 39'h3;
  assign T_8361 = ~ T_8360;
  assign T_8365 = T_8336 & mem_ctrl_branch;
  assign T_8369 = mem_waddr[0];
  assign T_8370 = io_imem_btb_update_bits_isJump & T_8369;
  assign T_8373 = T_7703 & id_ctrl_fp;
  assign T_8374 = dmem_resp_valid & T_8080;
  assign T_8375 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign T_8377 = ex_rs_0[63:38];
  assign T_8378 = alu_io_adder_out[39:38];
  assign T_8379 = $signed(T_8378);
  assign T_8381 = T_8377 == 26'h0;
  assign T_8383 = T_8377 == 26'h1;
  assign T_8384 = T_8381 | T_8383;
  assign T_8386 = $signed(T_8379) != $signed(2'sh0);
  assign T_8387 = $signed(T_8377);
  assign T_8389 = $signed(T_8387) == $signed(26'sh3ffffff);
  assign T_8392 = $signed(T_8387) == $signed(26'sh3fffffe);
  assign T_8393 = T_8389 | T_8392;
  assign T_8395 = $signed(T_8379) == $signed(2'sh3);
  assign T_8396 = T_8379[0];
  assign T_8397 = T_8393 ? T_8395 : T_8396;
  assign T_8398 = T_8384 ? T_8386 : T_8397;
  assign T_8399 = alu_io_adder_out[38:0];
  assign T_8400 = {T_8398,T_8399};
  assign T_8401 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign T_8402 = killm_common | mem_breakpoint;
  assign T_8404 = io_dmem_s1_kill == 1'h0;
  assign T_8405 = mem_xcpt & T_8404;
  assign T_8406 = {io_dmem_xcpt_pf_ld,io_dmem_xcpt_pf_st};
  assign T_8407 = {io_dmem_xcpt_ma_ld,io_dmem_xcpt_ma_st};
  assign T_8408 = {T_8407,T_8406};
  assign T_8410 = T_8408 != 4'h0;
  assign T_8411 = T_8410 | reset;
  assign T_8413 = T_8411 == 1'h0;
  assign T_8416 = replay_wb_common == 1'h0;
  assign T_8417 = T_7546 & T_8416;
  assign T_8420 = wb_xcpt & T_7534;
  assign T_8439_funct = T_8457;
  assign T_8439_rs2 = T_8456;
  assign T_8439_rs1 = T_8455;
  assign T_8439_xd = T_8454;
  assign T_8439_xs1 = T_8453;
  assign T_8439_xs2 = T_8452;
  assign T_8439_rd = T_8451;
  assign T_8439_opcode = T_8450;
  assign T_8449 = wb_reg_inst;
  assign T_8450 = T_8449[6:0];
  assign T_8451 = T_8449[11:7];
  assign T_8452 = T_8449[12];
  assign T_8453 = T_8449[13];
  assign T_8454 = T_8449[14];
  assign T_8455 = T_8449[19:15];
  assign T_8456 = T_8449[24:20];
  assign T_8457 = T_8449[31:25];
  assign T_8458 = csr_io_time[31:0];
  assign T_8460 = rf_wen ? rf_waddr : 5'h0;
  assign T_8461 = wb_reg_inst[19:15];
  assign T_8464 = wb_reg_inst[24:20];
  assign T_8468 = reset == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_155 = GEN_418[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_156 = GEN_419[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_157 = GEN_420[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_158 = GEN_421[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_159 = GEN_422[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_162 = GEN_423[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_163 = GEN_424[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_165 = GEN_425[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_166 = GEN_426[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_177 = GEN_427[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_178 = GEN_428[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_179 = GEN_429[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_180 = GEN_430[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_181 = GEN_431[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_182 = GEN_432[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_183 = GEN_433[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_184 = GEN_434[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_185 = GEN_435[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_186 = GEN_436[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_187 = GEN_437[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_188 = GEN_438[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_189 = GEN_439[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_190 = GEN_440[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_191 = GEN_441[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_192 = GEN_442[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_193 = GEN_443[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_194 = GEN_444[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_195 = GEN_445[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_196 = GEN_446[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_197 = GEN_447[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_198 = GEN_448[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_199 = GEN_449[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_200 = GEN_450[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_201 = GEN_451[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_202 = GEN_452[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_203 = GEN_453[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_204 = GEN_454[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_205 = GEN_455[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_206 = GEN_456[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_207 = GEN_457[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_208 = GEN_458[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_209 = GEN_459[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_210 = GEN_460[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_211 = GEN_461[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_212 = GEN_462[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_213 = GEN_463[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_214 = GEN_464[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_215 = GEN_465[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_216 = GEN_466[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_217 = GEN_467[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_218 = GEN_468[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_219 = GEN_469[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_220 = GEN_470[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_221 = GEN_471[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_222 = GEN_472[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_223 = GEN_473[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_224 = GEN_474[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_225 = GEN_475[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_226 = GEN_476[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_227 = GEN_477[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_228 = GEN_478[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_229 = GEN_479[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_230 = GEN_480[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_231 = GEN_481[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_232 = GEN_482[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_233 = GEN_483[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_234 = GEN_484[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_235 = GEN_485[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_236 = GEN_486[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_237 = GEN_487[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_238 = GEN_488[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_239 = GEN_489[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_240 = GEN_490[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_241 = GEN_491[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_242 = GEN_492[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_243 = GEN_493[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_244 = GEN_494[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_245 = GEN_495[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_246 = GEN_496[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_247 = GEN_497[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_248 = GEN_498[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_249 = GEN_499[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_250 = GEN_500[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_251 = GEN_501[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_252 = GEN_502[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_253 = GEN_503[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_254 = GEN_504[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_255 = GEN_505[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_256 = GEN_506[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_257 = GEN_507[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_258 = GEN_508[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_259 = GEN_509[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_260 = GEN_510[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_261 = GEN_511[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_262 = GEN_512[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_263 = GEN_513[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_264 = GEN_514[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_265 = GEN_515[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_266 = GEN_516[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_267 = GEN_517[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_268 = GEN_518[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_269 = GEN_519[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_270 = GEN_520[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_271 = GEN_521[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_272 = GEN_522[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_273 = {1{$random}};
  ex_ctrl_legal = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_274 = {1{$random}};
  ex_ctrl_fp = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_275 = {1{$random}};
  ex_ctrl_rocc = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_276 = {1{$random}};
  ex_ctrl_branch = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_277 = {1{$random}};
  ex_ctrl_jal = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_278 = {1{$random}};
  ex_ctrl_jalr = GEN_278[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_279 = {1{$random}};
  ex_ctrl_rxs2 = GEN_279[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_280 = {1{$random}};
  ex_ctrl_rxs1 = GEN_280[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_281 = {1{$random}};
  ex_ctrl_sel_alu2 = GEN_281[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_282 = {1{$random}};
  ex_ctrl_sel_alu1 = GEN_282[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_283 = {1{$random}};
  ex_ctrl_sel_imm = GEN_283[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_284 = {1{$random}};
  ex_ctrl_alu_dw = GEN_284[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_285 = {1{$random}};
  ex_ctrl_alu_fn = GEN_285[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_286 = {1{$random}};
  ex_ctrl_mem = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_287 = {1{$random}};
  ex_ctrl_mem_cmd = GEN_287[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_288 = {1{$random}};
  ex_ctrl_mem_type = GEN_288[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_289 = {1{$random}};
  ex_ctrl_rfs1 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_290 = {1{$random}};
  ex_ctrl_rfs2 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_291 = {1{$random}};
  ex_ctrl_rfs3 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_292 = {1{$random}};
  ex_ctrl_wfd = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_293 = {1{$random}};
  ex_ctrl_div = GEN_293[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_294 = {1{$random}};
  ex_ctrl_wxd = GEN_294[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_295 = {1{$random}};
  ex_ctrl_csr = GEN_295[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_296 = {1{$random}};
  ex_ctrl_fence_i = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_297 = {1{$random}};
  ex_ctrl_fence = GEN_297[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_298 = {1{$random}};
  ex_ctrl_amo = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_299 = {1{$random}};
  mem_ctrl_legal = GEN_299[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_300 = {1{$random}};
  mem_ctrl_fp = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_301 = {1{$random}};
  mem_ctrl_rocc = GEN_301[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_302 = {1{$random}};
  mem_ctrl_branch = GEN_302[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_303 = {1{$random}};
  mem_ctrl_jal = GEN_303[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_304 = {1{$random}};
  mem_ctrl_jalr = GEN_304[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_305 = {1{$random}};
  mem_ctrl_rxs2 = GEN_305[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_306 = {1{$random}};
  mem_ctrl_rxs1 = GEN_306[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_307 = {1{$random}};
  mem_ctrl_sel_alu2 = GEN_307[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_308 = {1{$random}};
  mem_ctrl_sel_alu1 = GEN_308[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_309 = {1{$random}};
  mem_ctrl_sel_imm = GEN_309[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_310 = {1{$random}};
  mem_ctrl_alu_dw = GEN_310[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_311 = {1{$random}};
  mem_ctrl_alu_fn = GEN_311[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_312 = {1{$random}};
  mem_ctrl_mem = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_313 = {1{$random}};
  mem_ctrl_mem_cmd = GEN_313[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_314 = {1{$random}};
  mem_ctrl_mem_type = GEN_314[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_315 = {1{$random}};
  mem_ctrl_rfs1 = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_316 = {1{$random}};
  mem_ctrl_rfs2 = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_317 = {1{$random}};
  mem_ctrl_rfs3 = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_318 = {1{$random}};
  mem_ctrl_wfd = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_319 = {1{$random}};
  mem_ctrl_div = GEN_319[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_320 = {1{$random}};
  mem_ctrl_wxd = GEN_320[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_321 = {1{$random}};
  mem_ctrl_csr = GEN_321[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_322 = {1{$random}};
  mem_ctrl_fence_i = GEN_322[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_323 = {1{$random}};
  mem_ctrl_fence = GEN_323[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_324 = {1{$random}};
  mem_ctrl_amo = GEN_324[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_325 = {1{$random}};
  wb_ctrl_legal = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_326 = {1{$random}};
  wb_ctrl_fp = GEN_326[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_327 = {1{$random}};
  wb_ctrl_rocc = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_328 = {1{$random}};
  wb_ctrl_branch = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_329 = {1{$random}};
  wb_ctrl_jal = GEN_329[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_330 = {1{$random}};
  wb_ctrl_jalr = GEN_330[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_331 = {1{$random}};
  wb_ctrl_rxs2 = GEN_331[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_332 = {1{$random}};
  wb_ctrl_rxs1 = GEN_332[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_333 = {1{$random}};
  wb_ctrl_sel_alu2 = GEN_333[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_334 = {1{$random}};
  wb_ctrl_sel_alu1 = GEN_334[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_335 = {1{$random}};
  wb_ctrl_sel_imm = GEN_335[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_336 = {1{$random}};
  wb_ctrl_alu_dw = GEN_336[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_337 = {1{$random}};
  wb_ctrl_alu_fn = GEN_337[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_338 = {1{$random}};
  wb_ctrl_mem = GEN_338[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_339 = {1{$random}};
  wb_ctrl_mem_cmd = GEN_339[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_340 = {1{$random}};
  wb_ctrl_mem_type = GEN_340[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_341 = {1{$random}};
  wb_ctrl_rfs1 = GEN_341[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_342 = {1{$random}};
  wb_ctrl_rfs2 = GEN_342[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_343 = {1{$random}};
  wb_ctrl_rfs3 = GEN_343[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_344 = {1{$random}};
  wb_ctrl_wfd = GEN_344[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_345 = {1{$random}};
  wb_ctrl_div = GEN_345[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_346 = {1{$random}};
  wb_ctrl_wxd = GEN_346[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_347 = {1{$random}};
  wb_ctrl_csr = GEN_347[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_348 = {1{$random}};
  wb_ctrl_fence_i = GEN_348[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_349 = {1{$random}};
  wb_ctrl_fence = GEN_349[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_350 = {1{$random}};
  wb_ctrl_amo = GEN_350[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_351 = {1{$random}};
  ex_reg_xcpt_interrupt = GEN_351[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_352 = {1{$random}};
  ex_reg_valid = GEN_352[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_353 = {1{$random}};
  ex_reg_rvc = GEN_353[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_354 = {1{$random}};
  ex_reg_btb_hit = GEN_354[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_355 = {1{$random}};
  ex_reg_btb_resp_taken = GEN_355[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_356 = {1{$random}};
  ex_reg_btb_resp_mask = GEN_356[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_357 = {1{$random}};
  ex_reg_btb_resp_bridx = GEN_357[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_358 = {2{$random}};
  ex_reg_btb_resp_target = GEN_358[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_359 = {1{$random}};
  ex_reg_btb_resp_entry = GEN_359[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_360 = {1{$random}};
  ex_reg_btb_resp_bht_history = GEN_360[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_361 = {1{$random}};
  ex_reg_btb_resp_bht_value = GEN_361[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_362 = {1{$random}};
  ex_reg_xcpt = GEN_362[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_363 = {1{$random}};
  ex_reg_flush_pipe = GEN_363[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_364 = {1{$random}};
  ex_reg_load_use = GEN_364[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_365 = {2{$random}};
  ex_reg_cause = GEN_365[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_366 = {1{$random}};
  ex_reg_replay = GEN_366[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_367 = {2{$random}};
  ex_reg_pc = GEN_367[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_368 = {1{$random}};
  ex_reg_inst = GEN_368[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_369 = {1{$random}};
  mem_reg_xcpt_interrupt = GEN_369[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_370 = {1{$random}};
  mem_reg_valid = GEN_370[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_371 = {1{$random}};
  mem_reg_rvc = GEN_371[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_372 = {1{$random}};
  mem_reg_btb_hit = GEN_372[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_373 = {1{$random}};
  mem_reg_btb_resp_taken = GEN_373[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_374 = {1{$random}};
  mem_reg_btb_resp_mask = GEN_374[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_375 = {1{$random}};
  mem_reg_btb_resp_bridx = GEN_375[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_376 = {2{$random}};
  mem_reg_btb_resp_target = GEN_376[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_377 = {1{$random}};
  mem_reg_btb_resp_entry = GEN_377[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_378 = {1{$random}};
  mem_reg_btb_resp_bht_history = GEN_378[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_379 = {1{$random}};
  mem_reg_btb_resp_bht_value = GEN_379[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_380 = {1{$random}};
  mem_reg_xcpt = GEN_380[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_381 = {1{$random}};
  mem_reg_replay = GEN_381[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_382 = {1{$random}};
  mem_reg_flush_pipe = GEN_382[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_383 = {2{$random}};
  mem_reg_cause = GEN_383[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_384 = {1{$random}};
  mem_reg_slow_bypass = GEN_384[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_385 = {1{$random}};
  mem_reg_load = GEN_385[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_386 = {1{$random}};
  mem_reg_store = GEN_386[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_387 = {2{$random}};
  mem_reg_pc = GEN_387[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_388 = {1{$random}};
  mem_reg_inst = GEN_388[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_389 = {2{$random}};
  mem_reg_wdata = GEN_389[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_390 = {2{$random}};
  mem_reg_rs2 = GEN_390[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_391 = {1{$random}};
  wb_reg_valid = GEN_391[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_392 = {1{$random}};
  wb_reg_xcpt = GEN_392[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_393 = {1{$random}};
  wb_reg_replay = GEN_393[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_394 = {2{$random}};
  wb_reg_cause = GEN_394[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_395 = {2{$random}};
  wb_reg_pc = GEN_395[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_396 = {1{$random}};
  wb_reg_inst = GEN_396[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_397 = {2{$random}};
  wb_reg_wdata = GEN_397[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_398 = {2{$random}};
  wb_reg_rs2 = GEN_398[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_399 = {1{$random}};
  id_reg_fence = GEN_399[0:0];
  `endif
  GEN_400 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    T_7352[initvar] = GEN_400[63:0];
  `endif
  GEN_401 = {2{$random}};
  GEN_402 = {2{$random}};
  `ifdef RANDOMIZE_REG_INIT
  GEN_403 = {1{$random}};
  ex_reg_rs_bypass_0 = GEN_403[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_404 = {1{$random}};
  ex_reg_rs_bypass_1 = GEN_404[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_405 = {1{$random}};
  ex_reg_rs_lsb_0 = GEN_405[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_406 = {1{$random}};
  ex_reg_rs_lsb_1 = GEN_406[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_407 = {2{$random}};
  ex_reg_rs_msb_0 = GEN_407[61:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_408 = {2{$random}};
  ex_reg_rs_msb_1 = GEN_408[61:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_409 = {1{$random}};
  T_8056 = GEN_409[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_410 = {1{$random}};
  T_8143 = GEN_410[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_411 = {1{$random}};
  T_8248 = GEN_411[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_412 = {1{$random}};
  dcache_blocked = GEN_412[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_413 = {1{$random}};
  rocc_blocked = GEN_413[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_414 = {2{$random}};
  T_8462 = GEN_414[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_415 = {2{$random}};
  T_8463 = GEN_415[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_416 = {2{$random}};
  T_8465 = GEN_416[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_417 = {2{$random}};
  T_8466 = GEN_417[63:0];
  `endif
  GEN_418 = {1{$random}};
  GEN_419 = {2{$random}};
  GEN_420 = {1{$random}};
  GEN_421 = {1{$random}};
  GEN_422 = {1{$random}};
  GEN_423 = {1{$random}};
  GEN_424 = {1{$random}};
  GEN_425 = {1{$random}};
  GEN_426 = {1{$random}};
  GEN_427 = {1{$random}};
  GEN_428 = {1{$random}};
  GEN_429 = {1{$random}};
  GEN_430 = {1{$random}};
  GEN_431 = {1{$random}};
  GEN_432 = {1{$random}};
  GEN_433 = {1{$random}};
  GEN_434 = {1{$random}};
  GEN_435 = {1{$random}};
  GEN_436 = {1{$random}};
  GEN_437 = {1{$random}};
  GEN_438 = {1{$random}};
  GEN_439 = {1{$random}};
  GEN_440 = {3{$random}};
  GEN_441 = {3{$random}};
  GEN_442 = {3{$random}};
  GEN_443 = {1{$random}};
  GEN_444 = {1{$random}};
  GEN_445 = {1{$random}};
  GEN_446 = {1{$random}};
  GEN_447 = {1{$random}};
  GEN_448 = {2{$random}};
  GEN_449 = {1{$random}};
  GEN_450 = {1{$random}};
  GEN_451 = {1{$random}};
  GEN_452 = {2{$random}};
  GEN_453 = {1{$random}};
  GEN_454 = {1{$random}};
  GEN_455 = {2{$random}};
  GEN_456 = {2{$random}};
  GEN_457 = {1{$random}};
  GEN_458 = {1{$random}};
  GEN_459 = {1{$random}};
  GEN_460 = {1{$random}};
  GEN_461 = {1{$random}};
  GEN_462 = {1{$random}};
  GEN_463 = {1{$random}};
  GEN_464 = {1{$random}};
  GEN_465 = {1{$random}};
  GEN_466 = {1{$random}};
  GEN_467 = {1{$random}};
  GEN_468 = {1{$random}};
  GEN_469 = {1{$random}};
  GEN_470 = {2{$random}};
  GEN_471 = {1{$random}};
  GEN_472 = {1{$random}};
  GEN_473 = {3{$random}};
  GEN_474 = {1{$random}};
  GEN_475 = {1{$random}};
  GEN_476 = {1{$random}};
  GEN_477 = {1{$random}};
  GEN_478 = {2{$random}};
  GEN_479 = {1{$random}};
  GEN_480 = {2{$random}};
  GEN_481 = {1{$random}};
  GEN_482 = {1{$random}};
  GEN_483 = {1{$random}};
  GEN_484 = {1{$random}};
  GEN_485 = {2{$random}};
  GEN_486 = {1{$random}};
  GEN_487 = {2{$random}};
  GEN_488 = {1{$random}};
  GEN_489 = {1{$random}};
  GEN_490 = {1{$random}};
  GEN_491 = {1{$random}};
  GEN_492 = {1{$random}};
  GEN_493 = {1{$random}};
  GEN_494 = {1{$random}};
  GEN_495 = {1{$random}};
  GEN_496 = {1{$random}};
  GEN_497 = {2{$random}};
  GEN_498 = {1{$random}};
  GEN_499 = {1{$random}};
  GEN_500 = {1{$random}};
  GEN_501 = {1{$random}};
  GEN_502 = {1{$random}};
  GEN_503 = {1{$random}};
  GEN_504 = {1{$random}};
  GEN_505 = {1{$random}};
  GEN_506 = {1{$random}};
  GEN_507 = {1{$random}};
  GEN_508 = {1{$random}};
  GEN_509 = {1{$random}};
  GEN_510 = {1{$random}};
  GEN_511 = {1{$random}};
  GEN_512 = {1{$random}};
  GEN_513 = {1{$random}};
  GEN_514 = {1{$random}};
  GEN_515 = {1{$random}};
  GEN_516 = {1{$random}};
  GEN_517 = {1{$random}};
  GEN_518 = {1{$random}};
  GEN_519 = {3{$random}};
  GEN_520 = {3{$random}};
  GEN_521 = {3{$random}};
  GEN_522 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_legal <= id_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_fp <= id_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rocc <= id_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_branch <= id_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_jal <= id_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_jalr <= id_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rxs2 <= id_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rxs1 <= id_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_xcpt) begin
          if(T_7722) begin
            ex_ctrl_sel_alu2 <= 2'h1;
          end else begin
            ex_ctrl_sel_alu2 <= 2'h0;
          end
        end else begin
          ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_xcpt) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_sel_imm <= id_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_xcpt) begin
          ex_ctrl_alu_dw <= 1'h1;
        end else begin
          ex_ctrl_alu_dw <= id_ctrl_alu_dw;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_xcpt) begin
          ex_ctrl_alu_fn <= 4'h0;
        end else begin
          ex_ctrl_alu_fn <= id_ctrl_alu_fn;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_mem <= id_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_mem_type <= id_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rfs1 <= id_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rfs2 <= id_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_rfs3 <= id_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_wfd <= id_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_div <= id_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_wxd <= id_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_csr_ren) begin
          ex_ctrl_csr <= 3'h5;
        end else begin
          ex_ctrl_csr <= id_ctrl_csr;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7726) begin
          ex_ctrl_fence_i <= 1'h1;
        end else begin
          ex_ctrl_fence_i <= id_ctrl_fence_i;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_fence <= id_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_ctrl_amo <= id_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_legal <= ex_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rocc <= ex_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu2 <= ex_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu1 <= ex_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_imm <= ex_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_dw <= ex_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_fn <= ex_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_type <= ex_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs3 <= ex_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence_i <= ex_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence <= ex_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_amo <= ex_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_legal <= mem_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_fp <= mem_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rocc <= mem_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_branch <= mem_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_jal <= mem_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_jalr <= mem_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rxs2 <= mem_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rxs1 <= mem_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_sel_alu2 <= mem_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_sel_alu1 <= mem_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_sel_imm <= mem_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_alu_dw <= mem_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_alu_fn <= mem_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_mem <= mem_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_mem_cmd <= mem_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_mem_type <= mem_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rfs1 <= mem_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rfs2 <= mem_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_rfs3 <= mem_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_wfd <= mem_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_div <= mem_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_wxd <= mem_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_csr <= mem_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_fence_i <= mem_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_fence <= mem_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_ctrl_amo <= mem_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt_interrupt <= T_7714;
    end
    if(1'h0) begin
    end else begin
      ex_reg_valid <= T_7703;
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(id_xcpt) begin
          if(T_7722) begin
            ex_reg_rvc <= 1'h1;
          end else begin
            ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
          end
        end else begin
          ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_hit <= ibuf_io_inst_0_bits_btb_hit;
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_taken <= ibuf_io_btb_resp_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_mask <= ibuf_io_btb_resp_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bridx <= ibuf_io_btb_resp_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_target <= ibuf_io_btb_resp_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_entry <= ibuf_io_btb_resp_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bht_history <= ibuf_io_btb_resp_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(ibuf_io_inst_0_bits_btb_hit) begin
        ex_reg_btb_resp_bht_value <= ibuf_io_btb_resp_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt <= T_7710;
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7726) begin
          ex_reg_flush_pipe <= 1'h1;
        end else begin
          ex_reg_flush_pipe <= T_7725;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_reg_load_use <= id_load_use;
      end
    end
    if(1'h0) begin
    end else begin
      if(id_xcpt) begin
        if(csr_io_interrupt) begin
          ex_reg_cause <= csr_io_interrupt_cause;
        end else begin
          ex_reg_cause <= {{60'd0}, T_7567};
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_replay <= T_7707;
    end
    if(1'h0) begin
    end else begin
      if(T_7762) begin
        ex_reg_pc <= ibuf_io_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7762) begin
        ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt_interrupt <= T_8000;
    end
    if(1'h0) begin
    end else begin
      mem_reg_valid <= T_7991;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_rvc <= ex_reg_rvc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_btb_hit <= ex_reg_btb_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt <= T_7997;
    end
    if(1'h0) begin
    end else begin
      mem_reg_replay <= T_7994;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_flush_pipe <= ex_reg_flush_pipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_xcpt) begin
        if(T_7794) begin
          mem_reg_cause <= ex_reg_cause;
        end else begin
          mem_reg_cause <= 64'h2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_load <= T_8010;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_store <= T_8018;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_wdata <= alu_io_out;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(T_8020) begin
          if(ex_reg_rs_bypass_1) begin
            mem_reg_rs2 <= GEN_1;
          end else begin
            mem_reg_rs2 <= T_7613;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      wb_reg_valid <= T_8060;
    end
    if(1'h0) begin
    end else begin
      wb_reg_xcpt <= T_8066;
    end
    if(1'h0) begin
    end else begin
      wb_reg_replay <= T_8063;
    end
    if(1'h0) begin
    end else begin
      if(mem_xcpt) begin
        if(T_8046) begin
          wb_reg_cause <= mem_reg_cause;
        end else begin
          wb_reg_cause <= {{60'd0}, mem_new_cause};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_reg_pc <= mem_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        wb_reg_inst <= mem_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        if(T_8072) begin
          wb_reg_wdata <= io_fpu_toint_data;
        end else begin
          wb_reg_wdata <= mem_int_wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_8068) begin
        if(mem_ctrl_rocc) begin
          wb_reg_rs2 <= mem_reg_rs2;
        end
      end
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T_7549;
    end
    if(T_7352_T_8104_en & T_7352_T_8104_mask) begin
      T_7352[T_7352_T_8104_addr] <= T_7352_T_8104_data;
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_reg_rs_bypass_0 <= T_7731;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        ex_reg_rs_bypass_1 <= T_7746;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7741) begin
          ex_reg_rs_lsb_0 <= T_7742;
        end else begin
          if(T_7577) begin
            ex_reg_rs_lsb_0 <= 2'h0;
          end else begin
            if(id_bypass_src_0_1) begin
              ex_reg_rs_lsb_0 <= 2'h1;
            end else begin
              if(id_bypass_src_0_2) begin
                ex_reg_rs_lsb_0 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_0 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7756) begin
          ex_reg_rs_lsb_1 <= T_7757;
        end else begin
          if(T_7581) begin
            ex_reg_rs_lsb_1 <= 2'h0;
          end else begin
            if(id_bypass_src_1_1) begin
              ex_reg_rs_lsb_1 <= 2'h1;
            end else begin
              if(id_bypass_src_1_2) begin
                ex_reg_rs_lsb_1 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_1 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7741) begin
          ex_reg_rs_msb_0 <= T_7743;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7703) begin
        if(T_7756) begin
          ex_reg_rs_msb_1 <= T_7758;
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_8056 <= T_8055;
    end
    if(reset) begin
      T_8143 <= 32'h0;
    end else begin
      if(T_8170) begin
        T_8143 <= T_8169;
      end else begin
        if(ll_wen) begin
          T_8143 <= T_8152;
        end
      end
    end
    if(reset) begin
      T_8248 <= 32'h0;
    end else begin
      if(T_8273) begin
        T_8248 <= T_8272;
      end else begin
        if(T_8266) begin
          T_8248 <= T_8265;
        end else begin
          if(T_8252) begin
            T_8248 <= T_8257;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      dcache_blocked <= T_8296;
    end
    if(1'h0) begin
    end else begin
      rocc_blocked <= T_8304;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_0) begin
        T_8462 <= GEN_0;
      end else begin
        T_8462 <= T_7612;
      end
    end
    if(1'h0) begin
    end else begin
      T_8463 <= T_8462;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_1) begin
        T_8465 <= GEN_1;
      end else begin
        T_8465 <= T_7613;
      end
    end
    if(1'h0) begin
    end else begin
      T_8466 <= T_8465;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8405 & T_8413) begin
          $fwrite(32'h80000002,"Assertion failed\n    at rocket.scala:632 assert(io.dmem.xcpt.asUInt.orR) // make sure s1_kill is exhaustive\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_8405 & T_8413) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8468) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_prci_id,T_8458,wb_valid,wb_reg_pc,T_8460,rf_wdata,rf_wen,T_8461,T_8463,T_8464,T_8466,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FlowThroughSerializer(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module ICache(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [19:0] io_s1_ppn,
  input   io_s1_kill,
  input   io_s2_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [15:0] io_resp_bits_data,
  output [63:0] io_resp_bits_datablock,
  input   io_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  reg [1:0] state;
  reg [31:0] GEN_5;
  reg  invalidated;
  reg [31:0] GEN_6;
  wire  stall;
  wire  rdy;
  reg [31:0] refill_addr;
  reg [31:0] GEN_7;
  wire  s1_any_tag_hit;
  reg  s1_valid;
  reg [31:0] GEN_8;
  reg [38:0] s1_vaddr;
  reg [63:0] GEN_9;
  wire [11:0] T_827;
  wire [31:0] s1_paddr;
  wire [19:0] s1_tag;
  wire  T_828;
  wire  s0_valid;
  wire [38:0] s0_vaddr;
  wire  T_830;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire [38:0] GEN_0;
  wire  T_839;
  wire  T_840;
  wire  out_valid;
  wire [5:0] s1_idx;
  wire  s1_hit;
  wire  T_842;
  wire  s1_miss;
  wire  T_845;
  wire  T_846;
  wire  T_848;
  wire [31:0] GEN_1;
  wire [19:0] refill_tag;
  wire  FlowThroughSerializer_1_clk;
  wire  FlowThroughSerializer_1_reset;
  wire  FlowThroughSerializer_1_io_in_ready;
  wire  FlowThroughSerializer_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_io_out_ready;
  wire  FlowThroughSerializer_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_io_cnt;
  wire  FlowThroughSerializer_1_io_done;
  wire  T_849;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_10;
  wire  T_852;
  wire [3:0] T_854;
  wire [2:0] T_855;
  wire [2:0] GEN_2;
  wire  refill_wrap;
  wire  T_856;
  wire  refill_done;
  reg [15:0] T_859;
  reg [31:0] GEN_11;
  wire  T_860;
  wire  T_861;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_865;
  wire  T_866;
  wire [14:0] T_867;
  wire [15:0] T_868;
  wire [15:0] GEN_3;
  wire [1:0] repl_way;
  reg [19:0] tag_array_0 [0:63];
  reg [31:0] GEN_12;
  wire [19:0] tag_array_0_tag_rdata_data;
  wire [5:0] tag_array_0_tag_rdata_addr;
  wire  tag_array_0_tag_rdata_en;
  reg [5:0] GEN_13;
  reg [31:0] GEN_14;
  wire [19:0] tag_array_0_T_910_data;
  wire [5:0] tag_array_0_T_910_addr;
  wire  tag_array_0_T_910_mask;
  wire  tag_array_0_T_910_en;
  reg [19:0] tag_array_1 [0:63];
  reg [31:0] GEN_15;
  wire [19:0] tag_array_1_tag_rdata_data;
  wire [5:0] tag_array_1_tag_rdata_addr;
  wire  tag_array_1_tag_rdata_en;
  reg [5:0] GEN_16;
  reg [31:0] GEN_17;
  wire [19:0] tag_array_1_T_910_data;
  wire [5:0] tag_array_1_T_910_addr;
  wire  tag_array_1_T_910_mask;
  wire  tag_array_1_T_910_en;
  reg [19:0] tag_array_2 [0:63];
  reg [31:0] GEN_18;
  wire [19:0] tag_array_2_tag_rdata_data;
  wire [5:0] tag_array_2_tag_rdata_addr;
  wire  tag_array_2_tag_rdata_en;
  reg [5:0] GEN_19;
  reg [31:0] GEN_20;
  wire [19:0] tag_array_2_T_910_data;
  wire [5:0] tag_array_2_T_910_addr;
  wire  tag_array_2_T_910_mask;
  wire  tag_array_2_T_910_en;
  reg [19:0] tag_array_3 [0:63];
  reg [31:0] GEN_21;
  wire [19:0] tag_array_3_tag_rdata_data;
  wire [5:0] tag_array_3_tag_rdata_addr;
  wire  tag_array_3_tag_rdata_en;
  reg [5:0] GEN_22;
  reg [31:0] GEN_23;
  wire [19:0] tag_array_3_T_910_data;
  wire [5:0] tag_array_3_T_910_addr;
  wire  tag_array_3_T_910_mask;
  wire  tag_array_3_T_910_en;
  wire [5:0] T_877;
  wire  T_879;
  wire  T_880;
  wire [5:0] T_882;
  wire [19:0] T_891_0;
  wire [19:0] T_891_1;
  wire [19:0] T_891_2;
  wire [19:0] T_891_3;
  wire  T_894;
  wire  T_896;
  wire  T_898;
  wire  T_900;
  wire  T_906_0;
  wire  T_906_1;
  wire  T_906_2;
  wire  T_906_3;
  wire  GEN_26;
  wire  GEN_28;
  wire  GEN_30;
  wire  GEN_32;
  reg [255:0] vb_array;
  reg [255:0] GEN_24;
  wire  T_914;
  wire  T_915;
  wire [7:0] T_916;
  wire [255:0] T_919;
  wire [255:0] T_920;
  wire [255:0] T_921;
  wire [255:0] GEN_33;
  wire [255:0] GEN_34;
  wire  GEN_35;
  wire  s1_disparity_0;
  wire  s1_disparity_1;
  wire  s1_disparity_2;
  wire  s1_disparity_3;
  wire  T_934;
  wire [6:0] T_936;
  wire [127:0] T_939;
  wire [255:0] GEN_87;
  wire [255:0] T_942;
  wire [255:0] T_943;
  wire [255:0] GEN_36;
  wire  T_945;
  wire [6:0] T_947;
  wire [127:0] T_950;
  wire [255:0] GEN_89;
  wire [255:0] T_953;
  wire [255:0] T_954;
  wire [255:0] GEN_37;
  wire  T_956;
  wire [7:0] T_958;
  wire [255:0] T_961;
  wire [255:0] T_964;
  wire [255:0] T_965;
  wire [255:0] GEN_38;
  wire  T_967;
  wire [7:0] T_969;
  wire [255:0] T_972;
  wire [255:0] T_975;
  wire [255:0] T_976;
  wire [255:0] GEN_39;
  wire  s1_tag_match_0;
  wire  s1_tag_match_1;
  wire  s1_tag_match_2;
  wire  s1_tag_match_3;
  wire  s1_tag_hit_0;
  wire  s1_tag_hit_1;
  wire  s1_tag_hit_2;
  wire  s1_tag_hit_3;
  wire [63:0] s1_dout_0;
  wire [63:0] s1_dout_1;
  wire [63:0] s1_dout_2;
  wire [63:0] s1_dout_3;
  wire  T_1000;
  wire [255:0] T_1004;
  wire  T_1005;
  wire  T_1007;
  wire [19:0] T_1011;
  wire  T_1012;
  wire  T_1013;
  wire [255:0] T_1024;
  wire  T_1025;
  wire  T_1027;
  wire [19:0] T_1031;
  wire  T_1032;
  wire  T_1033;
  wire [255:0] T_1044;
  wire  T_1045;
  wire  T_1047;
  wire [19:0] T_1051;
  wire  T_1052;
  wire  T_1053;
  wire [255:0] T_1064;
  wire  T_1065;
  wire  T_1067;
  wire [19:0] T_1071;
  wire  T_1072;
  wire  T_1073;
  wire  T_1079;
  wire  T_1080;
  wire  T_1081;
  wire  T_1082;
  wire  T_1083;
  wire  T_1084;
  wire  T_1086;
  wire  T_1087;
  reg [63:0] T_1090 [0:511];
  reg [63:0] GEN_25;
  wire [63:0] T_1090_T_1103_data;
  wire [8:0] T_1090_T_1103_addr;
  wire  T_1090_T_1103_en;
  reg [8:0] GEN_27;
  reg [31:0] GEN_29;
  wire [63:0] T_1090_T_1096_data;
  wire [8:0] T_1090_T_1096_addr;
  wire  T_1090_T_1096_mask;
  wire  T_1090_T_1096_en;
  wire  T_1093;
  wire [8:0] GEN_91;
  wire [8:0] T_1094;
  wire [8:0] GEN_92;
  wire [8:0] T_1095;
  wire [63:0] GEN_43;
  wire [8:0] T_1097;
  wire  T_1099;
  wire  T_1100;
  wire [8:0] T_1102;
  reg [63:0] T_1106 [0:511];
  reg [63:0] GEN_31;
  wire [63:0] T_1106_T_1119_data;
  wire [8:0] T_1106_T_1119_addr;
  wire  T_1106_T_1119_en;
  reg [8:0] GEN_40;
  reg [31:0] GEN_41;
  wire [63:0] T_1106_T_1112_data;
  wire [8:0] T_1106_T_1112_addr;
  wire  T_1106_T_1112_mask;
  wire  T_1106_T_1112_en;
  wire  T_1109;
  wire  T_1115;
  wire  T_1116;
  wire [8:0] T_1118;
  reg [63:0] T_1122 [0:511];
  reg [63:0] GEN_42;
  wire [63:0] T_1122_T_1135_data;
  wire [8:0] T_1122_T_1135_addr;
  wire  T_1122_T_1135_en;
  reg [8:0] GEN_44;
  reg [31:0] GEN_45;
  wire [63:0] T_1122_T_1128_data;
  wire [8:0] T_1122_T_1128_addr;
  wire  T_1122_T_1128_mask;
  wire  T_1122_T_1128_en;
  wire  T_1125;
  wire  T_1131;
  wire  T_1132;
  wire [8:0] T_1134;
  reg [63:0] T_1138 [0:511];
  reg [63:0] GEN_46;
  wire [63:0] T_1138_T_1151_data;
  wire [8:0] T_1138_T_1151_addr;
  wire  T_1138_T_1151_en;
  reg [8:0] GEN_47;
  reg [31:0] GEN_48;
  wire [63:0] T_1138_T_1144_data;
  wire [8:0] T_1138_T_1144_addr;
  wire  T_1138_T_1144_mask;
  wire  T_1138_T_1144_en;
  wire  T_1141;
  wire  T_1147;
  wire  T_1148;
  wire [8:0] T_1150;
  wire  T_1153;
  reg  T_1154;
  reg [31:0] GEN_49;
  wire  GEN_68;
  reg  T_1159_0;
  reg [31:0] GEN_50;
  reg  T_1159_1;
  reg [31:0] GEN_51;
  reg  T_1159_2;
  reg [31:0] GEN_52;
  reg  T_1159_3;
  reg [31:0] GEN_53;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  reg [63:0] T_1165_0;
  reg [63:0] GEN_54;
  reg [63:0] T_1165_1;
  reg [63:0] GEN_55;
  reg [63:0] T_1165_2;
  reg [63:0] GEN_56;
  reg [63:0] T_1165_3;
  reg [63:0] GEN_57;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire [63:0] GEN_75;
  wire [63:0] GEN_76;
  wire [63:0] T_1168;
  wire [63:0] T_1170;
  wire [63:0] T_1172;
  wire [63:0] T_1174;
  wire [63:0] T_1176;
  wire [63:0] T_1177;
  wire [63:0] T_1178;
  wire [63:0] T_1179;
  wire  T_1180;
  wire  T_1182;
  wire  T_1183;
  wire [25:0] T_1184;
  wire [25:0] T_1308_addr_block;
  wire [1:0] T_1308_client_xact_id;
  wire [2:0] T_1308_addr_beat;
  wire  T_1308_is_builtin_type;
  wire [2:0] T_1308_a_type;
  wire [10:0] T_1308_union;
  wire [63:0] T_1308_data;
  wire  T_1336;
  wire [1:0] GEN_77;
  wire [1:0] GEN_78;
  wire  GEN_79;
  wire  T_1338;
  wire [1:0] GEN_80;
  wire [1:0] GEN_81;
  wire [1:0] GEN_82;
  wire  T_1339;
  wire [1:0] GEN_83;
  wire [1:0] GEN_84;
  wire  T_1340;
  wire [1:0] GEN_85;
  wire [1:0] GEN_86;
  wire [15:0] GEN_4;
  reg [31:0] GEN_58;
  FlowThroughSerializer FlowThroughSerializer_1 (
    .clk(FlowThroughSerializer_1_clk),
    .reset(FlowThroughSerializer_1_reset),
    .io_in_ready(FlowThroughSerializer_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_io_in_bits_data),
    .io_out_ready(FlowThroughSerializer_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_io_out_bits_data),
    .io_cnt(FlowThroughSerializer_1_io_cnt),
    .io_done(FlowThroughSerializer_1_io_done)
  );
  assign io_resp_valid = T_1154;
  assign io_resp_bits_data = GEN_4;
  assign io_resp_bits_datablock = T_1179;
  assign io_mem_acquire_valid = T_1183;
  assign io_mem_acquire_bits_addr_block = T_1308_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1308_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1308_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1308_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1308_a_type;
  assign io_mem_acquire_bits_union = T_1308_union;
  assign io_mem_acquire_bits_data = T_1308_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign stall = io_resp_ready == 1'h0;
  assign rdy = T_846;
  assign s1_any_tag_hit = T_1087;
  assign T_827 = s1_vaddr[11:0];
  assign s1_paddr = {io_s1_ppn,T_827};
  assign s1_tag = s1_paddr[31:12];
  assign T_828 = s1_valid & stall;
  assign s0_valid = io_req_valid | T_828;
  assign s0_vaddr = T_828 ? s1_vaddr : io_req_bits_addr;
  assign T_830 = io_req_valid & rdy;
  assign T_833 = io_s1_kill == 1'h0;
  assign T_834 = T_828 & T_833;
  assign T_835 = T_830 | T_834;
  assign GEN_0 = T_830 ? io_req_bits_addr : s1_vaddr;
  assign T_839 = s1_valid & T_833;
  assign T_840 = state == 2'h0;
  assign out_valid = T_839 & T_840;
  assign s1_idx = s1_vaddr[11:6];
  assign s1_hit = out_valid & s1_any_tag_hit;
  assign T_842 = s1_any_tag_hit == 1'h0;
  assign s1_miss = out_valid & T_842;
  assign T_845 = s1_miss == 1'h0;
  assign T_846 = T_840 & T_845;
  assign T_848 = s1_miss & T_840;
  assign GEN_1 = T_848 ? s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:12];
  assign FlowThroughSerializer_1_clk = clk;
  assign FlowThroughSerializer_1_reset = reset;
  assign FlowThroughSerializer_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_io_out_ready = 1'h1;
  assign T_849 = FlowThroughSerializer_1_io_out_ready & FlowThroughSerializer_1_io_out_valid;
  assign T_852 = refill_cnt == 3'h7;
  assign T_854 = refill_cnt + 3'h1;
  assign T_855 = T_854[2:0];
  assign GEN_2 = T_849 ? T_855 : refill_cnt;
  assign refill_wrap = T_849 & T_852;
  assign T_856 = state == 2'h3;
  assign refill_done = T_856 & refill_wrap;
  assign T_860 = T_859[0];
  assign T_861 = T_859[2];
  assign T_862 = T_860 ^ T_861;
  assign T_863 = T_859[3];
  assign T_864 = T_862 ^ T_863;
  assign T_865 = T_859[5];
  assign T_866 = T_864 ^ T_865;
  assign T_867 = T_859[15:1];
  assign T_868 = {T_866,T_867};
  assign GEN_3 = s1_miss ? T_868 : T_859;
  assign repl_way = T_859[1:0];
  assign tag_array_0_tag_rdata_addr = T_882;
  assign tag_array_0_tag_rdata_en = T_880;
  assign tag_array_0_tag_rdata_data = tag_array_0[GEN_13];
  assign tag_array_0_T_910_data = T_891_0;
  assign tag_array_0_T_910_addr = s1_idx;
  assign tag_array_0_T_910_mask = GEN_26;
  assign tag_array_0_T_910_en = refill_done;
  assign tag_array_1_tag_rdata_addr = T_882;
  assign tag_array_1_tag_rdata_en = T_880;
  assign tag_array_1_tag_rdata_data = tag_array_1[GEN_16];
  assign tag_array_1_T_910_data = T_891_1;
  assign tag_array_1_T_910_addr = s1_idx;
  assign tag_array_1_T_910_mask = GEN_28;
  assign tag_array_1_T_910_en = refill_done;
  assign tag_array_2_tag_rdata_addr = T_882;
  assign tag_array_2_tag_rdata_en = T_880;
  assign tag_array_2_tag_rdata_data = tag_array_2[GEN_19];
  assign tag_array_2_T_910_data = T_891_2;
  assign tag_array_2_T_910_addr = s1_idx;
  assign tag_array_2_T_910_mask = GEN_30;
  assign tag_array_2_T_910_en = refill_done;
  assign tag_array_3_tag_rdata_addr = T_882;
  assign tag_array_3_tag_rdata_en = T_880;
  assign tag_array_3_tag_rdata_data = tag_array_3[GEN_22];
  assign tag_array_3_T_910_data = T_891_3;
  assign tag_array_3_T_910_addr = s1_idx;
  assign tag_array_3_T_910_mask = GEN_32;
  assign tag_array_3_T_910_en = refill_done;
  assign T_877 = s0_vaddr[11:6];
  assign T_879 = refill_done == 1'h0;
  assign T_880 = T_879 & s0_valid;
  assign T_882 = T_877;
  assign T_891_0 = refill_tag;
  assign T_891_1 = refill_tag;
  assign T_891_2 = refill_tag;
  assign T_891_3 = refill_tag;
  assign T_894 = repl_way == 2'h0;
  assign T_896 = repl_way == 2'h1;
  assign T_898 = repl_way == 2'h2;
  assign T_900 = repl_way == 2'h3;
  assign T_906_0 = T_894;
  assign T_906_1 = T_896;
  assign T_906_2 = T_898;
  assign T_906_3 = T_900;
  assign GEN_26 = refill_done ? T_906_0 : 1'h0;
  assign GEN_28 = refill_done ? T_906_1 : 1'h0;
  assign GEN_30 = refill_done ? T_906_2 : 1'h0;
  assign GEN_32 = refill_done ? T_906_3 : 1'h0;
  assign T_914 = invalidated == 1'h0;
  assign T_915 = refill_done & T_914;
  assign T_916 = {repl_way,s1_idx};
  assign T_919 = 256'h1 << T_916;
  assign T_920 = vb_array | T_919;
  assign T_921 = ~ vb_array;
  assign GEN_33 = T_915 ? T_920 : vb_array;
  assign GEN_34 = io_invalidate ? 256'h0 : GEN_33;
  assign GEN_35 = io_invalidate ? 1'h1 : invalidated;
  assign s1_disparity_0 = 1'h0;
  assign s1_disparity_1 = 1'h0;
  assign s1_disparity_2 = 1'h0;
  assign s1_disparity_3 = 1'h0;
  assign T_934 = s1_valid & s1_disparity_0;
  assign T_936 = {1'h0,s1_idx};
  assign T_939 = 128'h1 << T_936;
  assign GEN_87 = {{128'd0}, T_939};
  assign T_942 = T_921 | GEN_87;
  assign T_943 = ~ T_942;
  assign GEN_36 = T_934 ? T_943 : GEN_34;
  assign T_945 = s1_valid & s1_disparity_1;
  assign T_947 = {1'h1,s1_idx};
  assign T_950 = 128'h1 << T_947;
  assign GEN_89 = {{128'd0}, T_950};
  assign T_953 = T_921 | GEN_89;
  assign T_954 = ~ T_953;
  assign GEN_37 = T_945 ? T_954 : GEN_36;
  assign T_956 = s1_valid & s1_disparity_2;
  assign T_958 = {2'h2,s1_idx};
  assign T_961 = 256'h1 << T_958;
  assign T_964 = T_921 | T_961;
  assign T_965 = ~ T_964;
  assign GEN_38 = T_956 ? T_965 : GEN_37;
  assign T_967 = s1_valid & s1_disparity_3;
  assign T_969 = {2'h3,s1_idx};
  assign T_972 = 256'h1 << T_969;
  assign T_975 = T_921 | T_972;
  assign T_976 = ~ T_975;
  assign GEN_39 = T_967 ? T_976 : GEN_38;
  assign s1_tag_match_0 = T_1012;
  assign s1_tag_match_1 = T_1032;
  assign s1_tag_match_2 = T_1052;
  assign s1_tag_match_3 = T_1072;
  assign s1_tag_hit_0 = T_1013;
  assign s1_tag_hit_1 = T_1033;
  assign s1_tag_hit_2 = T_1053;
  assign s1_tag_hit_3 = T_1073;
  assign s1_dout_0 = T_1090_T_1103_data;
  assign s1_dout_1 = T_1106_T_1119_data;
  assign s1_dout_2 = T_1122_T_1135_data;
  assign s1_dout_3 = T_1138_T_1151_data;
  assign T_1000 = io_invalidate == 1'h0;
  assign T_1004 = vb_array >> T_936;
  assign T_1005 = T_1004[0];
  assign T_1007 = T_1000 & T_1005;
  assign T_1011 = tag_array_0_tag_rdata_data;
  assign T_1012 = T_1011 == s1_tag;
  assign T_1013 = T_1007 & s1_tag_match_0;
  assign T_1024 = vb_array >> T_947;
  assign T_1025 = T_1024[0];
  assign T_1027 = T_1000 & T_1025;
  assign T_1031 = tag_array_1_tag_rdata_data;
  assign T_1032 = T_1031 == s1_tag;
  assign T_1033 = T_1027 & s1_tag_match_1;
  assign T_1044 = vb_array >> T_958;
  assign T_1045 = T_1044[0];
  assign T_1047 = T_1000 & T_1045;
  assign T_1051 = tag_array_2_tag_rdata_data;
  assign T_1052 = T_1051 == s1_tag;
  assign T_1053 = T_1047 & s1_tag_match_2;
  assign T_1064 = vb_array >> T_969;
  assign T_1065 = T_1064[0];
  assign T_1067 = T_1000 & T_1065;
  assign T_1071 = tag_array_3_tag_rdata_data;
  assign T_1072 = T_1071 == s1_tag;
  assign T_1073 = T_1067 & s1_tag_match_3;
  assign T_1079 = s1_tag_hit_0 | s1_tag_hit_1;
  assign T_1080 = T_1079 | s1_tag_hit_2;
  assign T_1081 = T_1080 | s1_tag_hit_3;
  assign T_1082 = s1_disparity_0 | s1_disparity_1;
  assign T_1083 = T_1082 | s1_disparity_2;
  assign T_1084 = T_1083 | s1_disparity_3;
  assign T_1086 = T_1084 == 1'h0;
  assign T_1087 = T_1081 & T_1086;
  assign T_1090_T_1103_addr = T_1102;
  assign T_1090_T_1103_en = T_1100;
  assign T_1090_T_1103_data = T_1090[GEN_27];
  assign T_1090_T_1096_data = GEN_43;
  assign T_1090_T_1096_addr = T_1095;
  assign T_1090_T_1096_mask = T_1093;
  assign T_1090_T_1096_en = T_1093;
  assign T_1093 = FlowThroughSerializer_1_io_out_valid & T_894;
  assign GEN_91 = {{3'd0}, s1_idx};
  assign T_1094 = GEN_91 << 3;
  assign GEN_92 = {{6'd0}, refill_cnt};
  assign T_1095 = T_1094 | GEN_92;
  assign GEN_43 = FlowThroughSerializer_1_io_out_bits_data;
  assign T_1097 = s0_vaddr[11:3];
  assign T_1099 = T_1093 == 1'h0;
  assign T_1100 = T_1099 & s0_valid;
  assign T_1102 = T_1097;
  assign T_1106_T_1119_addr = T_1118;
  assign T_1106_T_1119_en = T_1116;
  assign T_1106_T_1119_data = T_1106[GEN_40];
  assign T_1106_T_1112_data = GEN_43;
  assign T_1106_T_1112_addr = T_1095;
  assign T_1106_T_1112_mask = T_1109;
  assign T_1106_T_1112_en = T_1109;
  assign T_1109 = FlowThroughSerializer_1_io_out_valid & T_896;
  assign T_1115 = T_1109 == 1'h0;
  assign T_1116 = T_1115 & s0_valid;
  assign T_1118 = T_1097;
  assign T_1122_T_1135_addr = T_1134;
  assign T_1122_T_1135_en = T_1132;
  assign T_1122_T_1135_data = T_1122[GEN_44];
  assign T_1122_T_1128_data = GEN_43;
  assign T_1122_T_1128_addr = T_1095;
  assign T_1122_T_1128_mask = T_1125;
  assign T_1122_T_1128_en = T_1125;
  assign T_1125 = FlowThroughSerializer_1_io_out_valid & T_898;
  assign T_1131 = T_1125 == 1'h0;
  assign T_1132 = T_1131 & s0_valid;
  assign T_1134 = T_1097;
  assign T_1138_T_1151_addr = T_1150;
  assign T_1138_T_1151_en = T_1148;
  assign T_1138_T_1151_data = T_1138[GEN_47];
  assign T_1138_T_1144_data = GEN_43;
  assign T_1138_T_1144_addr = T_1095;
  assign T_1138_T_1144_mask = T_1141;
  assign T_1138_T_1144_en = T_1141;
  assign T_1141 = FlowThroughSerializer_1_io_out_valid & T_900;
  assign T_1147 = T_1141 == 1'h0;
  assign T_1148 = T_1147 & s0_valid;
  assign T_1150 = T_1097;
  assign T_1153 = stall == 1'h0;
  assign GEN_68 = T_1153 ? s1_hit : T_1154;
  assign GEN_69 = T_1153 ? s1_tag_hit_0 : T_1159_0;
  assign GEN_70 = T_1153 ? s1_tag_hit_1 : T_1159_1;
  assign GEN_71 = T_1153 ? s1_tag_hit_2 : T_1159_2;
  assign GEN_72 = T_1153 ? s1_tag_hit_3 : T_1159_3;
  assign GEN_73 = T_1153 ? s1_dout_0 : T_1165_0;
  assign GEN_74 = T_1153 ? s1_dout_1 : T_1165_1;
  assign GEN_75 = T_1153 ? s1_dout_2 : T_1165_2;
  assign GEN_76 = T_1153 ? s1_dout_3 : T_1165_3;
  assign T_1168 = T_1159_0 ? T_1165_0 : 64'h0;
  assign T_1170 = T_1159_1 ? T_1165_1 : 64'h0;
  assign T_1172 = T_1159_2 ? T_1165_2 : 64'h0;
  assign T_1174 = T_1159_3 ? T_1165_3 : 64'h0;
  assign T_1176 = T_1168 | T_1170;
  assign T_1177 = T_1176 | T_1172;
  assign T_1178 = T_1177 | T_1174;
  assign T_1179 = T_1178;
  assign T_1180 = state == 2'h1;
  assign T_1182 = io_s2_kill == 1'h0;
  assign T_1183 = T_1180 & T_1182;
  assign T_1184 = refill_addr[31:6];
  assign T_1308_addr_block = T_1184;
  assign T_1308_client_xact_id = 2'h0;
  assign T_1308_addr_beat = 3'h0;
  assign T_1308_is_builtin_type = 1'h1;
  assign T_1308_a_type = 3'h1;
  assign T_1308_union = 11'hc1;
  assign T_1308_data = 64'h0;
  assign T_1336 = 2'h0 == state;
  assign GEN_77 = s1_miss ? 2'h1 : state;
  assign GEN_78 = T_1336 ? GEN_77 : state;
  assign GEN_79 = T_1336 ? 1'h0 : GEN_35;
  assign T_1338 = 2'h1 == state;
  assign GEN_80 = io_mem_acquire_ready ? 2'h2 : GEN_78;
  assign GEN_81 = io_s2_kill ? 2'h0 : GEN_80;
  assign GEN_82 = T_1338 ? GEN_81 : GEN_78;
  assign T_1339 = 2'h2 == state;
  assign GEN_83 = io_mem_grant_valid ? 2'h3 : GEN_82;
  assign GEN_84 = T_1339 ? GEN_83 : GEN_82;
  assign T_1340 = 2'h3 == state;
  assign GEN_85 = refill_done ? 2'h0 : GEN_84;
  assign GEN_86 = T_1340 ? GEN_85 : GEN_84;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_58[15:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  state = GEN_5[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  invalidated = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  refill_addr = GEN_7[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  s1_valid = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {2{$random}};
  s1_vaddr = GEN_9[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  refill_cnt = GEN_10[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  T_859 = GEN_11[15:0];
  `endif
  GEN_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = GEN_12[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[5:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = GEN_15[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  GEN_16 = GEN_17[5:0];
  `endif
  GEN_18 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = GEN_18[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  GEN_19 = GEN_20[5:0];
  `endif
  GEN_21 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = GEN_21[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  GEN_22 = GEN_23[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_24 = {8{$random}};
  vb_array = GEN_24[255:0];
  `endif
  GEN_25 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1090[initvar] = GEN_25[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  GEN_27 = GEN_29[8:0];
  `endif
  GEN_31 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1106[initvar] = GEN_31[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  GEN_40 = GEN_41[8:0];
  `endif
  GEN_42 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1122[initvar] = GEN_42[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  GEN_44 = GEN_45[8:0];
  `endif
  GEN_46 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1138[initvar] = GEN_46[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  GEN_47 = GEN_48[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  T_1154 = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  T_1159_0 = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  T_1159_1 = GEN_51[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  T_1159_2 = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  T_1159_3 = GEN_53[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {2{$random}};
  T_1165_0 = GEN_54[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {2{$random}};
  T_1165_1 = GEN_55[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {2{$random}};
  T_1165_2 = GEN_56[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {2{$random}};
  T_1165_3 = GEN_57[63:0];
  `endif
  GEN_58 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(T_1340) begin
        if(refill_done) begin
          state <= 2'h0;
        end else begin
          if(T_1339) begin
            if(io_mem_grant_valid) begin
              state <= 2'h3;
            end else begin
              if(T_1338) begin
                if(io_s2_kill) begin
                  state <= 2'h0;
                end else begin
                  if(io_mem_acquire_ready) begin
                    state <= 2'h2;
                  end else begin
                    if(T_1336) begin
                      if(s1_miss) begin
                        state <= 2'h1;
                      end
                    end
                  end
                end
              end else begin
                if(T_1336) begin
                  if(s1_miss) begin
                    state <= 2'h1;
                  end
                end
              end
            end
          end else begin
            if(T_1338) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  if(T_1336) begin
                    if(s1_miss) begin
                      state <= 2'h1;
                    end
                  end
                end
              end
            end else begin
              if(T_1336) begin
                if(s1_miss) begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if(T_1339) begin
          if(io_mem_grant_valid) begin
            state <= 2'h3;
          end else begin
            if(T_1338) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  state <= GEN_78;
                end
              end
            end else begin
              state <= GEN_78;
            end
          end
        end else begin
          if(T_1338) begin
            if(io_s2_kill) begin
              state <= 2'h0;
            end else begin
              if(io_mem_acquire_ready) begin
                state <= 2'h2;
              end else begin
                state <= GEN_78;
              end
            end
          end else begin
            state <= GEN_78;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1336) begin
        invalidated <= 1'h0;
      end else begin
        if(io_invalidate) begin
          invalidated <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_848) begin
        refill_addr <= s1_paddr;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_835;
    end
    if(1'h0) begin
    end else begin
      if(T_830) begin
        s1_vaddr <= io_req_bits_addr;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_849) begin
        refill_cnt <= T_855;
      end
    end
    if(reset) begin
      T_859 <= 16'h1;
    end else begin
      if(s1_miss) begin
        T_859 <= T_868;
      end
    end
    if(tag_array_0_tag_rdata_en) begin
      GEN_13 <= tag_array_0_tag_rdata_addr;
    end
    if(tag_array_0_T_910_en & tag_array_0_T_910_mask) begin
      tag_array_0[tag_array_0_T_910_addr] <= tag_array_0_T_910_data;
    end
    if(tag_array_1_tag_rdata_en) begin
      GEN_16 <= tag_array_1_tag_rdata_addr;
    end
    if(tag_array_1_T_910_en & tag_array_1_T_910_mask) begin
      tag_array_1[tag_array_1_T_910_addr] <= tag_array_1_T_910_data;
    end
    if(tag_array_2_tag_rdata_en) begin
      GEN_19 <= tag_array_2_tag_rdata_addr;
    end
    if(tag_array_2_T_910_en & tag_array_2_T_910_mask) begin
      tag_array_2[tag_array_2_T_910_addr] <= tag_array_2_T_910_data;
    end
    if(tag_array_3_tag_rdata_en) begin
      GEN_22 <= tag_array_3_tag_rdata_addr;
    end
    if(tag_array_3_T_910_en & tag_array_3_T_910_mask) begin
      tag_array_3[tag_array_3_T_910_addr] <= tag_array_3_T_910_data;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else begin
      if(T_967) begin
        vb_array <= T_976;
      end else begin
        if(T_956) begin
          vb_array <= T_965;
        end else begin
          if(T_945) begin
            vb_array <= T_954;
          end else begin
            if(T_934) begin
              vb_array <= T_943;
            end else begin
              if(io_invalidate) begin
                vb_array <= 256'h0;
              end else begin
                if(T_915) begin
                  vb_array <= T_920;
                end
              end
            end
          end
        end
      end
    end
    if(T_1090_T_1103_en) begin
      GEN_27 <= T_1090_T_1103_addr;
    end
    if(T_1090_T_1096_en & T_1090_T_1096_mask) begin
      T_1090[T_1090_T_1096_addr] <= T_1090_T_1096_data;
    end
    if(T_1106_T_1119_en) begin
      GEN_40 <= T_1106_T_1119_addr;
    end
    if(T_1106_T_1112_en & T_1106_T_1112_mask) begin
      T_1106[T_1106_T_1112_addr] <= T_1106_T_1112_data;
    end
    if(T_1122_T_1135_en) begin
      GEN_44 <= T_1122_T_1135_addr;
    end
    if(T_1122_T_1128_en & T_1122_T_1128_mask) begin
      T_1122[T_1122_T_1128_addr] <= T_1122_T_1128_data;
    end
    if(T_1138_T_1151_en) begin
      GEN_47 <= T_1138_T_1151_addr;
    end
    if(T_1138_T_1144_en & T_1138_T_1144_mask) begin
      T_1138[T_1138_T_1144_addr] <= T_1138_T_1144_data;
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1154 <= s1_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1159_0 <= s1_tag_hit_0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1159_1 <= s1_tag_hit_1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1159_2 <= s1_tag_hit_2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1159_3 <= s1_tag_hit_3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1165_0 <= s1_dout_0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1165_1 <= s1_dout_1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1165_2 <= s1_dout_2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1153) begin
        T_1165_3 <= s1_dout_3;
      end
    end
  end
endmodule
module TLB(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [27:0] io_req_bits_vpn,
  input   io_req_bits_passthrough,
  input   io_req_bits_instruction,
  input   io_req_bits_store,
  output  io_resp_miss,
  output [19:0] io_resp_ppn,
  output  io_resp_xcpt_ld,
  output  io_resp_xcpt_st,
  output  io_resp_xcpt_if,
  output  io_resp_cacheable,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie
);
  reg [7:0] valid;
  reg [31:0] GEN_18;
  reg [19:0] ppns_0;
  reg [31:0] GEN_27;
  reg [19:0] ppns_1;
  reg [31:0] GEN_60;
  reg [19:0] ppns_2;
  reg [31:0] GEN_64;
  reg [19:0] ppns_3;
  reg [31:0] GEN_66;
  reg [19:0] ppns_4;
  reg [31:0] GEN_67;
  reg [19:0] ppns_5;
  reg [31:0] GEN_68;
  reg [19:0] ppns_6;
  reg [31:0] GEN_69;
  reg [19:0] ppns_7;
  reg [31:0] GEN_70;
  reg [33:0] tags_0;
  reg [63:0] GEN_71;
  reg [33:0] tags_1;
  reg [63:0] GEN_72;
  reg [33:0] tags_2;
  reg [63:0] GEN_73;
  reg [33:0] tags_3;
  reg [63:0] GEN_74;
  reg [33:0] tags_4;
  reg [63:0] GEN_75;
  reg [33:0] tags_5;
  reg [63:0] GEN_76;
  reg [33:0] tags_6;
  reg [63:0] GEN_77;
  reg [33:0] tags_7;
  reg [63:0] GEN_78;
  reg [1:0] state;
  reg [31:0] GEN_79;
  reg [33:0] r_refill_tag;
  reg [63:0] GEN_80;
  reg [2:0] r_refill_waddr;
  reg [31:0] GEN_81;
  reg [27:0] r_req_vpn;
  reg [31:0] GEN_82;
  reg  r_req_passthrough;
  reg [31:0] GEN_83;
  reg  r_req_instruction;
  reg [31:0] GEN_84;
  reg  r_req_store;
  reg [31:0] GEN_85;
  wire  T_217;
  wire  do_mprv;
  wire [1:0] priv;
  wire  priv_s;
  wire  T_220;
  wire  T_222;
  wire  priv_uses_vm;
  wire [19:0] passthrough_ppn;
  wire [19:0] refill_ppn;
  wire [19:0] mpu_ppn;
  wire [31:0] GEN_59;
  wire [31:0] T_224;
  wire  T_228;
  wire [2:0] T_232;
  wire  T_234;
  wire  T_236;
  wire  T_237;
  wire [2:0] T_240;
  wire  T_242;
  wire  T_244;
  wire  T_245;
  wire [2:0] T_248;
  wire  T_250;
  wire  T_252;
  wire  T_253;
  wire [2:0] T_256;
  wire  T_258;
  wire  T_260;
  wire  T_261;
  wire [2:0] T_264;
  wire [2:0] T_269;
  wire [2:0] T_270;
  wire [2:0] T_271;
  wire [2:0] T_272;
  wire  prot_x;
  wire  prot_w;
  wire  prot_r;
  wire  T_280;
  wire  T_281;
  wire  T_282;
  wire [26:0] T_290;
  wire [33:0] lookup_tag;
  wire  T_292;
  wire  T_294;
  wire  T_296;
  wire  vm_enabled;
  wire  T_297;
  wire  T_298;
  wire  T_299;
  wire  hitsVec_0;
  wire  T_300;
  wire  T_301;
  wire  T_302;
  wire  hitsVec_1;
  wire  T_303;
  wire  T_304;
  wire  T_305;
  wire  hitsVec_2;
  wire  T_306;
  wire  T_307;
  wire  T_308;
  wire  hitsVec_3;
  wire  T_309;
  wire  T_310;
  wire  T_311;
  wire  hitsVec_4;
  wire  T_312;
  wire  T_313;
  wire  T_314;
  wire  hitsVec_5;
  wire  T_315;
  wire  T_316;
  wire  T_317;
  wire  hitsVec_6;
  wire  T_318;
  wire  T_319;
  wire  T_320;
  wire  hitsVec_7;
  wire  hitsVec_8;
  wire [1:0] T_322;
  wire [1:0] T_323;
  wire [3:0] T_324;
  wire [1:0] T_325;
  wire [1:0] T_326;
  wire [2:0] T_327;
  wire [4:0] T_328;
  wire [8:0] hits;
  reg [15:0] pte_array_reserved_for_hardware;
  reg [31:0] GEN_86;
  reg [37:0] pte_array_ppn;
  reg [63:0] GEN_87;
  reg [1:0] pte_array_reserved_for_software;
  reg [31:0] GEN_88;
  reg  pte_array_d;
  reg [31:0] GEN_89;
  reg  pte_array_a;
  reg [31:0] GEN_90;
  reg  pte_array_g;
  reg [31:0] GEN_91;
  reg  pte_array_u;
  reg [31:0] GEN_92;
  reg  pte_array_x;
  reg [31:0] GEN_93;
  reg  pte_array_w;
  reg [31:0] GEN_94;
  reg  pte_array_r;
  reg [31:0] GEN_95;
  reg  pte_array_v;
  reg [31:0] GEN_96;
  reg [7:0] u_array;
  reg [31:0] GEN_97;
  reg [7:0] sw_array;
  reg [31:0] GEN_98;
  reg [7:0] sx_array;
  reg [31:0] GEN_99;
  reg [7:0] sr_array;
  reg [31:0] GEN_100;
  reg [7:0] xr_array;
  reg [31:0] GEN_101;
  reg [7:0] cash_array;
  reg [31:0] GEN_102;
  reg [7:0] dirty_array;
  reg [31:0] GEN_103;
  wire [19:0] GEN_0;
  wire [19:0] GEN_2;
  wire [19:0] GEN_3;
  wire [19:0] GEN_4;
  wire [19:0] GEN_5;
  wire [19:0] GEN_6;
  wire [19:0] GEN_7;
  wire [19:0] GEN_8;
  wire [19:0] GEN_9;
  wire [33:0] GEN_1;
  wire [33:0] GEN_10;
  wire [33:0] GEN_11;
  wire [33:0] GEN_12;
  wire [33:0] GEN_13;
  wire [33:0] GEN_14;
  wire [33:0] GEN_15;
  wire [33:0] GEN_16;
  wire [33:0] GEN_17;
  wire [7:0] T_360;
  wire [7:0] T_361;
  wire [7:0] T_362;
  wire [7:0] T_363;
  wire [7:0] T_364;
  wire [7:0] T_365;
  wire  T_367;
  wire  T_368;
  wire  T_369;
  wire  T_370;
  wire  T_371;
  wire  T_372;
  wire [7:0] T_373;
  wire [7:0] T_375;
  wire [7:0] T_376;
  wire  T_382;
  wire  T_383;
  wire [7:0] T_384;
  wire [7:0] T_386;
  wire [7:0] T_387;
  wire  T_393;
  wire  T_394;
  wire [7:0] T_395;
  wire [7:0] T_397;
  wire [7:0] T_398;
  wire  T_405;
  wire [7:0] T_406;
  wire [7:0] T_408;
  wire [7:0] T_409;
  wire [7:0] T_410;
  wire [7:0] T_412;
  wire [7:0] T_413;
  wire [7:0] T_414;
  wire [7:0] T_416;
  wire [7:0] T_417;
  wire [19:0] GEN_19;
  wire [19:0] GEN_20;
  wire [19:0] GEN_21;
  wire [19:0] GEN_22;
  wire [19:0] GEN_23;
  wire [19:0] GEN_24;
  wire [19:0] GEN_25;
  wire [19:0] GEN_26;
  wire [33:0] GEN_28;
  wire [33:0] GEN_29;
  wire [33:0] GEN_30;
  wire [33:0] GEN_31;
  wire [33:0] GEN_32;
  wire [33:0] GEN_33;
  wire [33:0] GEN_34;
  wire [33:0] GEN_35;
  wire [7:0] GEN_36;
  wire [7:0] GEN_37;
  wire [7:0] GEN_38;
  wire [7:0] GEN_39;
  wire [7:0] GEN_40;
  wire [7:0] GEN_41;
  wire [7:0] GEN_42;
  wire [7:0] GEN_43;
  reg [7:0] T_419;
  reg [31:0] GEN_104;
  wire [7:0] T_420;
  wire  T_422;
  wire  T_424;
  wire  T_426;
  wire  T_427;
  wire  T_428;
  wire  T_429;
  wire  T_430;
  wire  T_431;
  wire  T_432;
  wire [2:0] T_442;
  wire [2:0] T_443;
  wire [2:0] T_444;
  wire [2:0] T_445;
  wire [2:0] T_446;
  wire [2:0] T_447;
  wire [2:0] T_448;
  wire [7:0] T_450;
  wire  T_451;
  wire [1:0] T_452;
  wire [7:0] T_453;
  wire  T_454;
  wire [2:0] T_455;
  wire [7:0] T_456;
  wire  T_457;
  wire [3:0] T_458;
  wire [2:0] T_459;
  wire [2:0] repl_waddr;
  wire [7:0] T_461;
  wire [7:0] T_462;
  wire [7:0] priv_ok;
  wire [7:0] T_463;
  wire [8:0] w_array;
  wire [7:0] T_464;
  wire [8:0] x_array;
  wire [7:0] T_466;
  wire [7:0] T_467;
  wire [7:0] T_468;
  wire [8:0] r_array;
  wire [8:0] c_array;
  wire  T_469;
  wire  T_470;
  wire  bad_va;
  wire [7:0] T_471;
  wire [8:0] T_473;
  wire [8:0] T_474;
  wire [8:0] GEN_61;
  wire [8:0] T_475;
  wire [8:0] GEN_62;
  wire [8:0] tlb_hits;
  wire  tlb_hit;
  wire  T_478;
  wire  T_479;
  wire  T_481;
  wire  tlb_miss;
  wire  T_483;
  wire  T_484;
  wire [3:0] T_486;
  wire [3:0] T_487;
  wire  T_489;
  wire [3:0] T_490;
  wire [1:0] T_491;
  wire [1:0] T_492;
  wire  T_494;
  wire [1:0] T_495;
  wire  T_496;
  wire [1:0] T_497;
  wire [2:0] T_498;
  wire  T_500;
  wire  T_502;
  wire [1:0] T_504;
  wire [7:0] GEN_63;
  wire [7:0] T_505;
  wire [7:0] T_506;
  wire [7:0] T_507;
  wire [7:0] T_508;
  wire [7:0] T_509;
  wire [1:0] T_510;
  wire  T_511;
  wire  T_513;
  wire [3:0] T_515;
  wire [7:0] GEN_65;
  wire [7:0] T_516;
  wire [7:0] T_517;
  wire [7:0] T_518;
  wire [7:0] T_519;
  wire [7:0] T_520;
  wire [2:0] T_521;
  wire  T_522;
  wire  T_524;
  wire [7:0] T_526;
  wire [7:0] T_527;
  wire [7:0] T_528;
  wire [7:0] T_529;
  wire [7:0] T_530;
  wire [7:0] T_531;
  wire [7:0] GEN_44;
  wire  T_533;
  wire [8:0] T_534;
  wire [8:0] T_535;
  wire  T_537;
  wire  T_538;
  wire [8:0] T_539;
  wire [8:0] T_540;
  wire  T_542;
  wire  T_543;
  wire [8:0] T_544;
  wire [8:0] T_545;
  wire  T_547;
  wire  T_548;
  wire [8:0] T_549;
  wire  T_551;
  wire  T_552;
  wire [19:0] T_554;
  wire [19:0] T_556;
  wire [19:0] T_558;
  wire [19:0] T_560;
  wire [19:0] T_562;
  wire [19:0] T_564;
  wire [19:0] T_566;
  wire [19:0] T_568;
  wire [19:0] T_570;
  wire [19:0] T_572;
  wire [19:0] T_573;
  wire [19:0] T_574;
  wire [19:0] T_575;
  wire [19:0] T_576;
  wire [19:0] T_577;
  wire [19:0] T_578;
  wire [19:0] T_579;
  wire [19:0] T_580;
  wire  T_581;
  wire  T_582;
  wire  T_583;
  wire [1:0] GEN_45;
  wire [33:0] GEN_46;
  wire [2:0] GEN_47;
  wire [27:0] GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire [1:0] GEN_52;
  wire [1:0] GEN_53;
  wire [1:0] GEN_54;
  wire [1:0] GEN_55;
  wire  T_585;
  wire  T_586;
  wire [1:0] GEN_56;
  wire [1:0] GEN_57;
  wire [7:0] GEN_58;
  assign io_req_ready = T_533;
  assign io_resp_miss = T_552;
  assign io_resp_ppn = T_580;
  assign io_resp_xcpt_ld = T_538;
  assign io_resp_xcpt_st = T_543;
  assign io_resp_xcpt_if = T_548;
  assign io_resp_cacheable = T_551;
  assign io_ptw_req_valid = T_581;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_pum = io_ptw_status_pum;
  assign io_ptw_req_bits_mxr = io_ptw_status_mxr;
  assign io_ptw_req_bits_addr = r_refill_tag[26:0];
  assign io_ptw_req_bits_store = r_req_store;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign T_217 = io_req_bits_instruction == 1'h0;
  assign do_mprv = io_ptw_status_mprv & T_217;
  assign priv = do_mprv ? io_ptw_status_mpp : io_ptw_status_prv;
  assign priv_s = priv == 2'h1;
  assign T_220 = priv <= 2'h1;
  assign T_222 = io_ptw_status_debug == 1'h0;
  assign priv_uses_vm = T_220 & T_222;
  assign passthrough_ppn = io_req_bits_vpn[19:0];
  assign refill_ppn = io_ptw_resp_bits_pte_ppn[19:0];
  assign mpu_ppn = io_ptw_resp_valid ? refill_ppn : passthrough_ppn;
  assign GEN_59 = {{12'd0}, mpu_ppn};
  assign T_224 = GEN_59 << 12;
  assign T_228 = T_224 < 32'h1000;
  assign T_232 = T_228 ? 3'h7 : 3'h0;
  assign T_234 = 32'h1000 <= T_224;
  assign T_236 = T_224 < 32'h2000;
  assign T_237 = T_234 & T_236;
  assign T_240 = T_237 ? 3'h5 : 3'h0;
  assign T_242 = 32'h40000000 <= T_224;
  assign T_244 = T_224 < 32'h44000000;
  assign T_245 = T_242 & T_244;
  assign T_248 = T_245 ? 3'h3 : 3'h0;
  assign T_250 = 32'h44000000 <= T_224;
  assign T_252 = T_224 < 32'h48000000;
  assign T_253 = T_250 & T_252;
  assign T_256 = T_253 ? 3'h3 : 3'h0;
  assign T_258 = 32'h80000000 <= T_224;
  assign T_260 = T_224 < 32'h90000000;
  assign T_261 = T_258 & T_260;
  assign T_264 = T_261 ? 3'h7 : 3'h0;
  assign T_269 = T_232 | T_240;
  assign T_270 = T_269 | T_248;
  assign T_271 = T_270 | T_256;
  assign T_272 = T_271 | T_264;
  assign prot_x = T_282;
  assign prot_w = T_281;
  assign prot_r = T_280;
  assign T_280 = T_272[0];
  assign T_281 = T_272[1];
  assign T_282 = T_272[2];
  assign T_290 = io_req_bits_vpn[26:0];
  assign lookup_tag = {io_ptw_ptbr_asid,T_290};
  assign T_292 = io_ptw_status_vm[3];
  assign T_294 = T_292 & priv_uses_vm;
  assign T_296 = io_req_bits_passthrough == 1'h0;
  assign vm_enabled = T_294 & T_296;
  assign T_297 = valid[0];
  assign T_298 = T_297 & vm_enabled;
  assign T_299 = tags_0 == lookup_tag;
  assign hitsVec_0 = T_298 & T_299;
  assign T_300 = valid[1];
  assign T_301 = T_300 & vm_enabled;
  assign T_302 = tags_1 == lookup_tag;
  assign hitsVec_1 = T_301 & T_302;
  assign T_303 = valid[2];
  assign T_304 = T_303 & vm_enabled;
  assign T_305 = tags_2 == lookup_tag;
  assign hitsVec_2 = T_304 & T_305;
  assign T_306 = valid[3];
  assign T_307 = T_306 & vm_enabled;
  assign T_308 = tags_3 == lookup_tag;
  assign hitsVec_3 = T_307 & T_308;
  assign T_309 = valid[4];
  assign T_310 = T_309 & vm_enabled;
  assign T_311 = tags_4 == lookup_tag;
  assign hitsVec_4 = T_310 & T_311;
  assign T_312 = valid[5];
  assign T_313 = T_312 & vm_enabled;
  assign T_314 = tags_5 == lookup_tag;
  assign hitsVec_5 = T_313 & T_314;
  assign T_315 = valid[6];
  assign T_316 = T_315 & vm_enabled;
  assign T_317 = tags_6 == lookup_tag;
  assign hitsVec_6 = T_316 & T_317;
  assign T_318 = valid[7];
  assign T_319 = T_318 & vm_enabled;
  assign T_320 = tags_7 == lookup_tag;
  assign hitsVec_7 = T_319 & T_320;
  assign hitsVec_8 = vm_enabled == 1'h0;
  assign T_322 = {hitsVec_1,hitsVec_0};
  assign T_323 = {hitsVec_3,hitsVec_2};
  assign T_324 = {T_323,T_322};
  assign T_325 = {hitsVec_5,hitsVec_4};
  assign T_326 = {hitsVec_8,hitsVec_7};
  assign T_327 = {T_326,hitsVec_6};
  assign T_328 = {T_327,T_325};
  assign hits = {T_328,T_324};
  assign GEN_0 = io_ptw_resp_bits_pte_ppn[19:0];
  assign GEN_2 = 3'h0 == r_refill_waddr ? GEN_0 : ppns_0;
  assign GEN_3 = 3'h1 == r_refill_waddr ? GEN_0 : ppns_1;
  assign GEN_4 = 3'h2 == r_refill_waddr ? GEN_0 : ppns_2;
  assign GEN_5 = 3'h3 == r_refill_waddr ? GEN_0 : ppns_3;
  assign GEN_6 = 3'h4 == r_refill_waddr ? GEN_0 : ppns_4;
  assign GEN_7 = 3'h5 == r_refill_waddr ? GEN_0 : ppns_5;
  assign GEN_8 = 3'h6 == r_refill_waddr ? GEN_0 : ppns_6;
  assign GEN_9 = 3'h7 == r_refill_waddr ? GEN_0 : ppns_7;
  assign GEN_1 = r_refill_tag;
  assign GEN_10 = 3'h0 == r_refill_waddr ? GEN_1 : tags_0;
  assign GEN_11 = 3'h1 == r_refill_waddr ? GEN_1 : tags_1;
  assign GEN_12 = 3'h2 == r_refill_waddr ? GEN_1 : tags_2;
  assign GEN_13 = 3'h3 == r_refill_waddr ? GEN_1 : tags_3;
  assign GEN_14 = 3'h4 == r_refill_waddr ? GEN_1 : tags_4;
  assign GEN_15 = 3'h5 == r_refill_waddr ? GEN_1 : tags_5;
  assign GEN_16 = 3'h6 == r_refill_waddr ? GEN_1 : tags_6;
  assign GEN_17 = 3'h7 == r_refill_waddr ? GEN_1 : tags_7;
  assign T_360 = 8'h1 << r_refill_waddr;
  assign T_361 = valid | T_360;
  assign T_362 = u_array | T_360;
  assign T_363 = ~ T_360;
  assign T_364 = u_array & T_363;
  assign T_365 = io_ptw_resp_bits_pte_u ? T_362 : T_364;
  assign T_367 = io_ptw_resp_bits_pte_w == 1'h0;
  assign T_368 = io_ptw_resp_bits_pte_x & T_367;
  assign T_369 = io_ptw_resp_bits_pte_r | T_368;
  assign T_370 = io_ptw_resp_bits_pte_v & T_369;
  assign T_371 = T_370 & io_ptw_resp_bits_pte_w;
  assign T_372 = T_371 & prot_w;
  assign T_373 = sw_array | T_360;
  assign T_375 = sw_array & T_363;
  assign T_376 = T_372 ? T_373 : T_375;
  assign T_382 = T_370 & io_ptw_resp_bits_pte_x;
  assign T_383 = T_382 & prot_x;
  assign T_384 = sx_array | T_360;
  assign T_386 = sx_array & T_363;
  assign T_387 = T_383 ? T_384 : T_386;
  assign T_393 = T_370 & io_ptw_resp_bits_pte_r;
  assign T_394 = T_393 & prot_r;
  assign T_395 = sr_array | T_360;
  assign T_397 = sr_array & T_363;
  assign T_398 = T_394 ? T_395 : T_397;
  assign T_405 = T_382 & prot_r;
  assign T_406 = xr_array | T_360;
  assign T_408 = xr_array & T_363;
  assign T_409 = T_405 ? T_406 : T_408;
  assign T_410 = cash_array | T_360;
  assign T_412 = cash_array & T_363;
  assign T_413 = T_261 ? T_410 : T_412;
  assign T_414 = dirty_array | T_360;
  assign T_416 = dirty_array & T_363;
  assign T_417 = io_ptw_resp_bits_pte_d ? T_414 : T_416;
  assign GEN_19 = io_ptw_resp_valid ? GEN_2 : ppns_0;
  assign GEN_20 = io_ptw_resp_valid ? GEN_3 : ppns_1;
  assign GEN_21 = io_ptw_resp_valid ? GEN_4 : ppns_2;
  assign GEN_22 = io_ptw_resp_valid ? GEN_5 : ppns_3;
  assign GEN_23 = io_ptw_resp_valid ? GEN_6 : ppns_4;
  assign GEN_24 = io_ptw_resp_valid ? GEN_7 : ppns_5;
  assign GEN_25 = io_ptw_resp_valid ? GEN_8 : ppns_6;
  assign GEN_26 = io_ptw_resp_valid ? GEN_9 : ppns_7;
  assign GEN_28 = io_ptw_resp_valid ? GEN_10 : tags_0;
  assign GEN_29 = io_ptw_resp_valid ? GEN_11 : tags_1;
  assign GEN_30 = io_ptw_resp_valid ? GEN_12 : tags_2;
  assign GEN_31 = io_ptw_resp_valid ? GEN_13 : tags_3;
  assign GEN_32 = io_ptw_resp_valid ? GEN_14 : tags_4;
  assign GEN_33 = io_ptw_resp_valid ? GEN_15 : tags_5;
  assign GEN_34 = io_ptw_resp_valid ? GEN_16 : tags_6;
  assign GEN_35 = io_ptw_resp_valid ? GEN_17 : tags_7;
  assign GEN_36 = io_ptw_resp_valid ? T_361 : valid;
  assign GEN_37 = io_ptw_resp_valid ? T_365 : u_array;
  assign GEN_38 = io_ptw_resp_valid ? T_376 : sw_array;
  assign GEN_39 = io_ptw_resp_valid ? T_387 : sx_array;
  assign GEN_40 = io_ptw_resp_valid ? T_398 : sr_array;
  assign GEN_41 = io_ptw_resp_valid ? T_409 : xr_array;
  assign GEN_42 = io_ptw_resp_valid ? T_413 : cash_array;
  assign GEN_43 = io_ptw_resp_valid ? T_417 : dirty_array;
  assign T_420 = ~ valid;
  assign T_422 = T_420 == 8'h0;
  assign T_424 = T_422 == 1'h0;
  assign T_426 = T_420[0];
  assign T_427 = T_420[1];
  assign T_428 = T_420[2];
  assign T_429 = T_420[3];
  assign T_430 = T_420[4];
  assign T_431 = T_420[5];
  assign T_432 = T_420[6];
  assign T_442 = T_432 ? 3'h6 : 3'h7;
  assign T_443 = T_431 ? 3'h5 : T_442;
  assign T_444 = T_430 ? 3'h4 : T_443;
  assign T_445 = T_429 ? 3'h3 : T_444;
  assign T_446 = T_428 ? 3'h2 : T_445;
  assign T_447 = T_427 ? 3'h1 : T_446;
  assign T_448 = T_426 ? 3'h0 : T_447;
  assign T_450 = T_419 >> 1'h1;
  assign T_451 = T_450[0];
  assign T_452 = {1'h1,T_451};
  assign T_453 = T_419 >> T_452;
  assign T_454 = T_453[0];
  assign T_455 = {T_452,T_454};
  assign T_456 = T_419 >> T_455;
  assign T_457 = T_456[0];
  assign T_458 = {T_455,T_457};
  assign T_459 = T_458[2:0];
  assign repl_waddr = T_424 ? T_448 : T_459;
  assign T_461 = io_ptw_status_pum ? u_array : 8'h0;
  assign T_462 = ~ T_461;
  assign priv_ok = priv_s ? T_462 : u_array;
  assign T_463 = priv_ok & sw_array;
  assign w_array = {prot_w,T_463};
  assign T_464 = priv_ok & sx_array;
  assign x_array = {prot_x,T_464};
  assign T_466 = io_ptw_status_mxr ? xr_array : 8'h0;
  assign T_467 = sr_array | T_466;
  assign T_468 = priv_ok & T_467;
  assign r_array = {prot_r,T_468};
  assign c_array = {T_261,cash_array};
  assign T_469 = io_req_bits_vpn[27];
  assign T_470 = io_req_bits_vpn[26];
  assign bad_va = T_469 != T_470;
  assign T_471 = hits[7:0];
  assign T_473 = io_req_bits_store ? w_array : 9'h0;
  assign T_474 = ~ T_473;
  assign GEN_61 = {{1'd0}, dirty_array};
  assign T_475 = GEN_61 | T_474;
  assign GEN_62 = {{1'd0}, T_471};
  assign tlb_hits = GEN_62 & T_475;
  assign tlb_hit = tlb_hits != 9'h0;
  assign T_478 = bad_va == 1'h0;
  assign T_479 = vm_enabled & T_478;
  assign T_481 = tlb_hit == 1'h0;
  assign tlb_miss = T_479 & T_481;
  assign T_483 = tlb_miss == 1'h0;
  assign T_484 = io_req_valid & T_483;
  assign T_486 = T_471[7:4];
  assign T_487 = T_471[3:0];
  assign T_489 = T_486 != 4'h0;
  assign T_490 = T_486 | T_487;
  assign T_491 = T_490[3:2];
  assign T_492 = T_490[1:0];
  assign T_494 = T_491 != 2'h0;
  assign T_495 = T_491 | T_492;
  assign T_496 = T_495[1];
  assign T_497 = {T_494,T_496};
  assign T_498 = {T_489,T_497};
  assign T_500 = T_498[2];
  assign T_502 = T_500 == 1'h0;
  assign T_504 = 2'h1 << 1'h1;
  assign GEN_63 = {{6'd0}, T_504};
  assign T_505 = T_419 | GEN_63;
  assign T_506 = ~ T_419;
  assign T_507 = T_506 | GEN_63;
  assign T_508 = ~ T_507;
  assign T_509 = T_502 ? T_505 : T_508;
  assign T_510 = {1'h1,T_500};
  assign T_511 = T_498[1];
  assign T_513 = T_511 == 1'h0;
  assign T_515 = 4'h1 << T_510;
  assign GEN_65 = {{4'd0}, T_515};
  assign T_516 = T_509 | GEN_65;
  assign T_517 = ~ T_509;
  assign T_518 = T_517 | GEN_65;
  assign T_519 = ~ T_518;
  assign T_520 = T_513 ? T_516 : T_519;
  assign T_521 = {T_510,T_511};
  assign T_522 = T_498[0];
  assign T_524 = T_522 == 1'h0;
  assign T_526 = 8'h1 << T_521;
  assign T_527 = T_520 | T_526;
  assign T_528 = ~ T_520;
  assign T_529 = T_528 | T_526;
  assign T_530 = ~ T_529;
  assign T_531 = T_524 ? T_527 : T_530;
  assign GEN_44 = T_484 ? T_531 : T_419;
  assign T_533 = state == 2'h0;
  assign T_534 = ~ r_array;
  assign T_535 = T_534 & hits;
  assign T_537 = T_535 != 9'h0;
  assign T_538 = bad_va | T_537;
  assign T_539 = ~ w_array;
  assign T_540 = T_539 & hits;
  assign T_542 = T_540 != 9'h0;
  assign T_543 = bad_va | T_542;
  assign T_544 = ~ x_array;
  assign T_545 = T_544 & hits;
  assign T_547 = T_545 != 9'h0;
  assign T_548 = bad_va | T_547;
  assign T_549 = c_array & hits;
  assign T_551 = T_549 != 9'h0;
  assign T_552 = io_ptw_resp_valid | tlb_miss;
  assign T_554 = hitsVec_0 ? ppns_0 : 20'h0;
  assign T_556 = hitsVec_1 ? ppns_1 : 20'h0;
  assign T_558 = hitsVec_2 ? ppns_2 : 20'h0;
  assign T_560 = hitsVec_3 ? ppns_3 : 20'h0;
  assign T_562 = hitsVec_4 ? ppns_4 : 20'h0;
  assign T_564 = hitsVec_5 ? ppns_5 : 20'h0;
  assign T_566 = hitsVec_6 ? ppns_6 : 20'h0;
  assign T_568 = hitsVec_7 ? ppns_7 : 20'h0;
  assign T_570 = hitsVec_8 ? passthrough_ppn : 20'h0;
  assign T_572 = T_554 | T_556;
  assign T_573 = T_572 | T_558;
  assign T_574 = T_573 | T_560;
  assign T_575 = T_574 | T_562;
  assign T_576 = T_575 | T_564;
  assign T_577 = T_576 | T_566;
  assign T_578 = T_577 | T_568;
  assign T_579 = T_578 | T_570;
  assign T_580 = T_579;
  assign T_581 = state == 2'h1;
  assign T_582 = io_req_ready & io_req_valid;
  assign T_583 = T_582 & tlb_miss;
  assign GEN_45 = T_583 ? 2'h1 : state;
  assign GEN_46 = T_583 ? lookup_tag : r_refill_tag;
  assign GEN_47 = T_583 ? repl_waddr : r_refill_waddr;
  assign GEN_48 = T_583 ? io_req_bits_vpn : r_req_vpn;
  assign GEN_49 = T_583 ? io_req_bits_passthrough : r_req_passthrough;
  assign GEN_50 = T_583 ? io_req_bits_instruction : r_req_instruction;
  assign GEN_51 = T_583 ? io_req_bits_store : r_req_store;
  assign GEN_52 = io_ptw_invalidate ? 2'h0 : GEN_45;
  assign GEN_53 = io_ptw_invalidate ? 2'h3 : 2'h2;
  assign GEN_54 = io_ptw_req_ready ? GEN_53 : GEN_52;
  assign GEN_55 = T_581 ? GEN_54 : GEN_45;
  assign T_585 = state == 2'h2;
  assign T_586 = T_585 & io_ptw_invalidate;
  assign GEN_56 = T_586 ? 2'h3 : GEN_55;
  assign GEN_57 = io_ptw_resp_valid ? 2'h0 : GEN_56;
  assign GEN_58 = io_ptw_invalidate ? 8'h0 : GEN_36;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  valid = GEN_18[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  ppns_0 = GEN_27[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {1{$random}};
  ppns_1 = GEN_60[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_64 = {1{$random}};
  ppns_2 = GEN_64[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_66 = {1{$random}};
  ppns_3 = GEN_66[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_67 = {1{$random}};
  ppns_4 = GEN_67[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_68 = {1{$random}};
  ppns_5 = GEN_68[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_69 = {1{$random}};
  ppns_6 = GEN_69[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_70 = {1{$random}};
  ppns_7 = GEN_70[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_71 = {2{$random}};
  tags_0 = GEN_71[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_72 = {2{$random}};
  tags_1 = GEN_72[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_73 = {2{$random}};
  tags_2 = GEN_73[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_74 = {2{$random}};
  tags_3 = GEN_74[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_75 = {2{$random}};
  tags_4 = GEN_75[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_76 = {2{$random}};
  tags_5 = GEN_76[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_77 = {2{$random}};
  tags_6 = GEN_77[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {2{$random}};
  tags_7 = GEN_78[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  state = GEN_79[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {2{$random}};
  r_refill_tag = GEN_80[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  r_refill_waddr = GEN_81[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  r_req_vpn = GEN_82[27:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  r_req_passthrough = GEN_83[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  r_req_instruction = GEN_84[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  r_req_store = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pte_array_reserved_for_hardware = GEN_86[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {2{$random}};
  pte_array_ppn = GEN_87[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  pte_array_reserved_for_software = GEN_88[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {1{$random}};
  pte_array_d = GEN_89[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  pte_array_a = GEN_90[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {1{$random}};
  pte_array_g = GEN_91[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {1{$random}};
  pte_array_u = GEN_92[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {1{$random}};
  pte_array_x = GEN_93[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {1{$random}};
  pte_array_w = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {1{$random}};
  pte_array_r = GEN_95[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {1{$random}};
  pte_array_v = GEN_96[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  u_array = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  sw_array = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  sx_array = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  sr_array = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  xr_array = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  cash_array = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  dirty_array = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  T_419 = GEN_104[7:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      valid <= 8'h0;
    end else begin
      if(io_ptw_invalidate) begin
        valid <= 8'h0;
      end else begin
        if(io_ptw_resp_valid) begin
          valid <= T_361;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h0 == r_refill_waddr) begin
          ppns_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h1 == r_refill_waddr) begin
          ppns_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h2 == r_refill_waddr) begin
          ppns_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h3 == r_refill_waddr) begin
          ppns_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          ppns_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          ppns_5 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          ppns_6 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          ppns_7 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h0 == r_refill_waddr) begin
          tags_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h1 == r_refill_waddr) begin
          tags_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h2 == r_refill_waddr) begin
          tags_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h3 == r_refill_waddr) begin
          tags_3 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h4 == r_refill_waddr) begin
          tags_4 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h5 == r_refill_waddr) begin
          tags_5 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h6 == r_refill_waddr) begin
          tags_6 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(3'h7 == r_refill_waddr) begin
          tags_7 <= GEN_1;
        end
      end
    end
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(io_ptw_resp_valid) begin
        state <= 2'h0;
      end else begin
        if(T_586) begin
          state <= 2'h3;
        end else begin
          if(T_581) begin
            if(io_ptw_req_ready) begin
              if(io_ptw_invalidate) begin
                state <= 2'h3;
              end else begin
                state <= 2'h2;
              end
            end else begin
              if(io_ptw_invalidate) begin
                state <= 2'h0;
              end else begin
                if(T_583) begin
                  state <= 2'h1;
                end
              end
            end
          end else begin
            if(T_583) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        r_refill_tag <= lookup_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        if(T_424) begin
          if(T_426) begin
            r_refill_waddr <= 3'h0;
          end else begin
            if(T_427) begin
              r_refill_waddr <= 3'h1;
            end else begin
              if(T_428) begin
                r_refill_waddr <= 3'h2;
              end else begin
                if(T_429) begin
                  r_refill_waddr <= 3'h3;
                end else begin
                  if(T_430) begin
                    r_refill_waddr <= 3'h4;
                  end else begin
                    if(T_431) begin
                      r_refill_waddr <= 3'h5;
                    end else begin
                      if(T_432) begin
                        r_refill_waddr <= 3'h6;
                      end else begin
                        r_refill_waddr <= 3'h7;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          r_refill_waddr <= T_459;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        r_req_vpn <= io_req_bits_vpn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        r_req_passthrough <= io_req_bits_passthrough;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        r_req_instruction <= io_req_bits_instruction;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_583) begin
        r_req_store <= io_req_bits_store;
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(io_ptw_resp_bits_pte_u) begin
          u_array <= T_362;
        end else begin
          u_array <= T_364;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_372) begin
          sw_array <= T_373;
        end else begin
          sw_array <= T_375;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_383) begin
          sx_array <= T_384;
        end else begin
          sx_array <= T_386;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_394) begin
          sr_array <= T_395;
        end else begin
          sr_array <= T_397;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_405) begin
          xr_array <= T_406;
        end else begin
          xr_array <= T_408;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_261) begin
          cash_array <= T_410;
        end else begin
          cash_array <= T_412;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(io_ptw_resp_bits_pte_d) begin
          dirty_array <= T_414;
        end else begin
          dirty_array <= T_416;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_484) begin
        if(T_524) begin
          T_419 <= T_527;
        end else begin
          T_419 <= T_530;
        end
      end
    end
  end
endmodule
module BTB(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  output  io_resp_valid,
  output  io_resp_bits_taken,
  output [1:0] io_resp_bits_mask,
  output  io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [5:0] io_resp_bits_entry,
  output [6:0] io_resp_bits_bht_history,
  output [1:0] io_resp_bits_bht_value,
  input   io_btb_update_valid,
  input   io_btb_update_bits_prediction_valid,
  input   io_btb_update_bits_prediction_bits_taken,
  input  [1:0] io_btb_update_bits_prediction_bits_mask,
  input   io_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_btb_update_bits_prediction_bits_target,
  input  [5:0] io_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_btb_update_bits_pc,
  input  [38:0] io_btb_update_bits_target,
  input   io_btb_update_bits_taken,
  input   io_btb_update_bits_isValid,
  input   io_btb_update_bits_isJump,
  input   io_btb_update_bits_isReturn,
  input  [38:0] io_btb_update_bits_br_pc,
  input   io_bht_update_valid,
  input   io_bht_update_bits_prediction_valid,
  input   io_bht_update_bits_prediction_bits_taken,
  input  [1:0] io_bht_update_bits_prediction_bits_mask,
  input   io_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_bht_update_bits_prediction_bits_target,
  input  [5:0] io_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_bht_update_bits_pc,
  input   io_bht_update_bits_taken,
  input   io_bht_update_bits_mispredict,
  input   io_ras_update_valid,
  input   io_ras_update_bits_isCall,
  input   io_ras_update_bits_isReturn,
  input  [38:0] io_ras_update_bits_returnAddr,
  input   io_ras_update_bits_prediction_valid,
  input   io_ras_update_bits_prediction_bits_taken,
  input  [1:0] io_ras_update_bits_prediction_bits_mask,
  input   io_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_ras_update_bits_prediction_bits_target,
  input  [5:0] io_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_ras_update_bits_prediction_bits_bht_value
);
  reg [10:0] idxs_0;
  reg [31:0] GEN_231;
  reg [10:0] idxs_1;
  reg [31:0] GEN_272;
  reg [10:0] idxs_2;
  reg [31:0] GEN_313;
  reg [10:0] idxs_3;
  reg [31:0] GEN_354;
  reg [10:0] idxs_4;
  reg [31:0] GEN_398;
  reg [10:0] idxs_5;
  reg [31:0] GEN_448;
  reg [10:0] idxs_6;
  reg [31:0] GEN_449;
  reg [10:0] idxs_7;
  reg [31:0] GEN_450;
  reg [10:0] idxs_8;
  reg [31:0] GEN_451;
  reg [10:0] idxs_9;
  reg [31:0] GEN_452;
  reg [10:0] idxs_10;
  reg [31:0] GEN_456;
  reg [10:0] idxs_11;
  reg [31:0] GEN_463;
  reg [10:0] idxs_12;
  reg [31:0] GEN_473;
  reg [10:0] idxs_13;
  reg [31:0] GEN_480;
  reg [10:0] idxs_14;
  reg [31:0] GEN_482;
  reg [10:0] idxs_15;
  reg [31:0] GEN_484;
  reg [10:0] idxs_16;
  reg [31:0] GEN_490;
  reg [10:0] idxs_17;
  reg [31:0] GEN_491;
  reg [10:0] idxs_18;
  reg [31:0] GEN_492;
  reg [10:0] idxs_19;
  reg [31:0] GEN_493;
  reg [10:0] idxs_20;
  reg [31:0] GEN_494;
  reg [10:0] idxs_21;
  reg [31:0] GEN_495;
  reg [10:0] idxs_22;
  reg [31:0] GEN_496;
  reg [10:0] idxs_23;
  reg [31:0] GEN_497;
  reg [10:0] idxs_24;
  reg [31:0] GEN_498;
  reg [10:0] idxs_25;
  reg [31:0] GEN_499;
  reg [10:0] idxs_26;
  reg [31:0] GEN_500;
  reg [10:0] idxs_27;
  reg [31:0] GEN_501;
  reg [10:0] idxs_28;
  reg [31:0] GEN_502;
  reg [10:0] idxs_29;
  reg [31:0] GEN_503;
  reg [10:0] idxs_30;
  reg [31:0] GEN_504;
  reg [10:0] idxs_31;
  reg [31:0] GEN_505;
  reg [10:0] idxs_32;
  reg [31:0] GEN_506;
  reg [10:0] idxs_33;
  reg [31:0] GEN_507;
  reg [10:0] idxs_34;
  reg [31:0] GEN_508;
  reg [10:0] idxs_35;
  reg [31:0] GEN_509;
  reg [10:0] idxs_36;
  reg [31:0] GEN_510;
  reg [10:0] idxs_37;
  reg [31:0] GEN_511;
  reg [10:0] idxs_38;
  reg [31:0] GEN_512;
  reg [10:0] idxs_39;
  reg [31:0] GEN_513;
  reg [2:0] idxPages_0;
  reg [31:0] GEN_514;
  reg [2:0] idxPages_1;
  reg [31:0] GEN_515;
  reg [2:0] idxPages_2;
  reg [31:0] GEN_516;
  reg [2:0] idxPages_3;
  reg [31:0] GEN_517;
  reg [2:0] idxPages_4;
  reg [31:0] GEN_518;
  reg [2:0] idxPages_5;
  reg [31:0] GEN_519;
  reg [2:0] idxPages_6;
  reg [31:0] GEN_520;
  reg [2:0] idxPages_7;
  reg [31:0] GEN_521;
  reg [2:0] idxPages_8;
  reg [31:0] GEN_522;
  reg [2:0] idxPages_9;
  reg [31:0] GEN_523;
  reg [2:0] idxPages_10;
  reg [31:0] GEN_524;
  reg [2:0] idxPages_11;
  reg [31:0] GEN_525;
  reg [2:0] idxPages_12;
  reg [31:0] GEN_526;
  reg [2:0] idxPages_13;
  reg [31:0] GEN_527;
  reg [2:0] idxPages_14;
  reg [31:0] GEN_528;
  reg [2:0] idxPages_15;
  reg [31:0] GEN_529;
  reg [2:0] idxPages_16;
  reg [31:0] GEN_530;
  reg [2:0] idxPages_17;
  reg [31:0] GEN_531;
  reg [2:0] idxPages_18;
  reg [31:0] GEN_532;
  reg [2:0] idxPages_19;
  reg [31:0] GEN_533;
  reg [2:0] idxPages_20;
  reg [31:0] GEN_534;
  reg [2:0] idxPages_21;
  reg [31:0] GEN_535;
  reg [2:0] idxPages_22;
  reg [31:0] GEN_536;
  reg [2:0] idxPages_23;
  reg [31:0] GEN_537;
  reg [2:0] idxPages_24;
  reg [31:0] GEN_538;
  reg [2:0] idxPages_25;
  reg [31:0] GEN_539;
  reg [2:0] idxPages_26;
  reg [31:0] GEN_540;
  reg [2:0] idxPages_27;
  reg [31:0] GEN_541;
  reg [2:0] idxPages_28;
  reg [31:0] GEN_542;
  reg [2:0] idxPages_29;
  reg [31:0] GEN_543;
  reg [2:0] idxPages_30;
  reg [31:0] GEN_544;
  reg [2:0] idxPages_31;
  reg [31:0] GEN_545;
  reg [2:0] idxPages_32;
  reg [31:0] GEN_546;
  reg [2:0] idxPages_33;
  reg [31:0] GEN_547;
  reg [2:0] idxPages_34;
  reg [31:0] GEN_548;
  reg [2:0] idxPages_35;
  reg [31:0] GEN_549;
  reg [2:0] idxPages_36;
  reg [31:0] GEN_550;
  reg [2:0] idxPages_37;
  reg [31:0] GEN_551;
  reg [2:0] idxPages_38;
  reg [31:0] GEN_552;
  reg [2:0] idxPages_39;
  reg [31:0] GEN_553;
  reg [10:0] tgts_0;
  reg [31:0] GEN_554;
  reg [10:0] tgts_1;
  reg [31:0] GEN_555;
  reg [10:0] tgts_2;
  reg [31:0] GEN_556;
  reg [10:0] tgts_3;
  reg [31:0] GEN_557;
  reg [10:0] tgts_4;
  reg [31:0] GEN_558;
  reg [10:0] tgts_5;
  reg [31:0] GEN_559;
  reg [10:0] tgts_6;
  reg [31:0] GEN_560;
  reg [10:0] tgts_7;
  reg [31:0] GEN_561;
  reg [10:0] tgts_8;
  reg [31:0] GEN_562;
  reg [10:0] tgts_9;
  reg [31:0] GEN_563;
  reg [10:0] tgts_10;
  reg [31:0] GEN_564;
  reg [10:0] tgts_11;
  reg [31:0] GEN_565;
  reg [10:0] tgts_12;
  reg [31:0] GEN_566;
  reg [10:0] tgts_13;
  reg [31:0] GEN_567;
  reg [10:0] tgts_14;
  reg [31:0] GEN_568;
  reg [10:0] tgts_15;
  reg [31:0] GEN_569;
  reg [10:0] tgts_16;
  reg [31:0] GEN_570;
  reg [10:0] tgts_17;
  reg [31:0] GEN_571;
  reg [10:0] tgts_18;
  reg [31:0] GEN_572;
  reg [10:0] tgts_19;
  reg [31:0] GEN_573;
  reg [10:0] tgts_20;
  reg [31:0] GEN_574;
  reg [10:0] tgts_21;
  reg [31:0] GEN_575;
  reg [10:0] tgts_22;
  reg [31:0] GEN_576;
  reg [10:0] tgts_23;
  reg [31:0] GEN_577;
  reg [10:0] tgts_24;
  reg [31:0] GEN_578;
  reg [10:0] tgts_25;
  reg [31:0] GEN_579;
  reg [10:0] tgts_26;
  reg [31:0] GEN_580;
  reg [10:0] tgts_27;
  reg [31:0] GEN_581;
  reg [10:0] tgts_28;
  reg [31:0] GEN_582;
  reg [10:0] tgts_29;
  reg [31:0] GEN_583;
  reg [10:0] tgts_30;
  reg [31:0] GEN_584;
  reg [10:0] tgts_31;
  reg [31:0] GEN_585;
  reg [10:0] tgts_32;
  reg [31:0] GEN_586;
  reg [10:0] tgts_33;
  reg [31:0] GEN_587;
  reg [10:0] tgts_34;
  reg [31:0] GEN_588;
  reg [10:0] tgts_35;
  reg [31:0] GEN_589;
  reg [10:0] tgts_36;
  reg [31:0] GEN_590;
  reg [10:0] tgts_37;
  reg [31:0] GEN_591;
  reg [10:0] tgts_38;
  reg [31:0] GEN_592;
  reg [10:0] tgts_39;
  reg [31:0] GEN_593;
  reg [2:0] tgtPages_0;
  reg [31:0] GEN_594;
  reg [2:0] tgtPages_1;
  reg [31:0] GEN_595;
  reg [2:0] tgtPages_2;
  reg [31:0] GEN_596;
  reg [2:0] tgtPages_3;
  reg [31:0] GEN_597;
  reg [2:0] tgtPages_4;
  reg [31:0] GEN_598;
  reg [2:0] tgtPages_5;
  reg [31:0] GEN_599;
  reg [2:0] tgtPages_6;
  reg [31:0] GEN_600;
  reg [2:0] tgtPages_7;
  reg [31:0] GEN_601;
  reg [2:0] tgtPages_8;
  reg [31:0] GEN_602;
  reg [2:0] tgtPages_9;
  reg [31:0] GEN_603;
  reg [2:0] tgtPages_10;
  reg [31:0] GEN_604;
  reg [2:0] tgtPages_11;
  reg [31:0] GEN_605;
  reg [2:0] tgtPages_12;
  reg [31:0] GEN_606;
  reg [2:0] tgtPages_13;
  reg [31:0] GEN_607;
  reg [2:0] tgtPages_14;
  reg [31:0] GEN_608;
  reg [2:0] tgtPages_15;
  reg [31:0] GEN_609;
  reg [2:0] tgtPages_16;
  reg [31:0] GEN_610;
  reg [2:0] tgtPages_17;
  reg [31:0] GEN_611;
  reg [2:0] tgtPages_18;
  reg [31:0] GEN_612;
  reg [2:0] tgtPages_19;
  reg [31:0] GEN_613;
  reg [2:0] tgtPages_20;
  reg [31:0] GEN_614;
  reg [2:0] tgtPages_21;
  reg [31:0] GEN_615;
  reg [2:0] tgtPages_22;
  reg [31:0] GEN_616;
  reg [2:0] tgtPages_23;
  reg [31:0] GEN_617;
  reg [2:0] tgtPages_24;
  reg [31:0] GEN_618;
  reg [2:0] tgtPages_25;
  reg [31:0] GEN_619;
  reg [2:0] tgtPages_26;
  reg [31:0] GEN_620;
  reg [2:0] tgtPages_27;
  reg [31:0] GEN_621;
  reg [2:0] tgtPages_28;
  reg [31:0] GEN_622;
  reg [2:0] tgtPages_29;
  reg [31:0] GEN_623;
  reg [2:0] tgtPages_30;
  reg [31:0] GEN_624;
  reg [2:0] tgtPages_31;
  reg [31:0] GEN_625;
  reg [2:0] tgtPages_32;
  reg [31:0] GEN_626;
  reg [2:0] tgtPages_33;
  reg [31:0] GEN_627;
  reg [2:0] tgtPages_34;
  reg [31:0] GEN_628;
  reg [2:0] tgtPages_35;
  reg [31:0] GEN_629;
  reg [2:0] tgtPages_36;
  reg [31:0] GEN_630;
  reg [2:0] tgtPages_37;
  reg [31:0] GEN_631;
  reg [2:0] tgtPages_38;
  reg [31:0] GEN_632;
  reg [2:0] tgtPages_39;
  reg [31:0] GEN_633;
  reg [26:0] pages_0;
  reg [31:0] GEN_634;
  reg [26:0] pages_1;
  reg [31:0] GEN_635;
  reg [26:0] pages_2;
  reg [31:0] GEN_636;
  reg [26:0] pages_3;
  reg [31:0] GEN_637;
  reg [26:0] pages_4;
  reg [31:0] GEN_638;
  reg [26:0] pages_5;
  reg [31:0] GEN_639;
  reg [5:0] pageValid;
  reg [31:0] GEN_640;
  wire [7:0] T_606;
  wire [5:0] idxPagesOH_0;
  wire [7:0] T_608;
  wire [5:0] idxPagesOH_1;
  wire [7:0] T_610;
  wire [5:0] idxPagesOH_2;
  wire [7:0] T_612;
  wire [5:0] idxPagesOH_3;
  wire [7:0] T_614;
  wire [5:0] idxPagesOH_4;
  wire [7:0] T_616;
  wire [5:0] idxPagesOH_5;
  wire [7:0] T_618;
  wire [5:0] idxPagesOH_6;
  wire [7:0] T_620;
  wire [5:0] idxPagesOH_7;
  wire [7:0] T_622;
  wire [5:0] idxPagesOH_8;
  wire [7:0] T_624;
  wire [5:0] idxPagesOH_9;
  wire [7:0] T_626;
  wire [5:0] idxPagesOH_10;
  wire [7:0] T_628;
  wire [5:0] idxPagesOH_11;
  wire [7:0] T_630;
  wire [5:0] idxPagesOH_12;
  wire [7:0] T_632;
  wire [5:0] idxPagesOH_13;
  wire [7:0] T_634;
  wire [5:0] idxPagesOH_14;
  wire [7:0] T_636;
  wire [5:0] idxPagesOH_15;
  wire [7:0] T_638;
  wire [5:0] idxPagesOH_16;
  wire [7:0] T_640;
  wire [5:0] idxPagesOH_17;
  wire [7:0] T_642;
  wire [5:0] idxPagesOH_18;
  wire [7:0] T_644;
  wire [5:0] idxPagesOH_19;
  wire [7:0] T_646;
  wire [5:0] idxPagesOH_20;
  wire [7:0] T_648;
  wire [5:0] idxPagesOH_21;
  wire [7:0] T_650;
  wire [5:0] idxPagesOH_22;
  wire [7:0] T_652;
  wire [5:0] idxPagesOH_23;
  wire [7:0] T_654;
  wire [5:0] idxPagesOH_24;
  wire [7:0] T_656;
  wire [5:0] idxPagesOH_25;
  wire [7:0] T_658;
  wire [5:0] idxPagesOH_26;
  wire [7:0] T_660;
  wire [5:0] idxPagesOH_27;
  wire [7:0] T_662;
  wire [5:0] idxPagesOH_28;
  wire [7:0] T_664;
  wire [5:0] idxPagesOH_29;
  wire [7:0] T_666;
  wire [5:0] idxPagesOH_30;
  wire [7:0] T_668;
  wire [5:0] idxPagesOH_31;
  wire [7:0] T_670;
  wire [5:0] idxPagesOH_32;
  wire [7:0] T_672;
  wire [5:0] idxPagesOH_33;
  wire [7:0] T_674;
  wire [5:0] idxPagesOH_34;
  wire [7:0] T_676;
  wire [5:0] idxPagesOH_35;
  wire [7:0] T_678;
  wire [5:0] idxPagesOH_36;
  wire [7:0] T_680;
  wire [5:0] idxPagesOH_37;
  wire [7:0] T_682;
  wire [5:0] idxPagesOH_38;
  wire [7:0] T_684;
  wire [5:0] idxPagesOH_39;
  wire [7:0] T_686;
  wire [5:0] tgtPagesOH_0;
  wire [7:0] T_688;
  wire [5:0] tgtPagesOH_1;
  wire [7:0] T_690;
  wire [5:0] tgtPagesOH_2;
  wire [7:0] T_692;
  wire [5:0] tgtPagesOH_3;
  wire [7:0] T_694;
  wire [5:0] tgtPagesOH_4;
  wire [7:0] T_696;
  wire [5:0] tgtPagesOH_5;
  wire [7:0] T_698;
  wire [5:0] tgtPagesOH_6;
  wire [7:0] T_700;
  wire [5:0] tgtPagesOH_7;
  wire [7:0] T_702;
  wire [5:0] tgtPagesOH_8;
  wire [7:0] T_704;
  wire [5:0] tgtPagesOH_9;
  wire [7:0] T_706;
  wire [5:0] tgtPagesOH_10;
  wire [7:0] T_708;
  wire [5:0] tgtPagesOH_11;
  wire [7:0] T_710;
  wire [5:0] tgtPagesOH_12;
  wire [7:0] T_712;
  wire [5:0] tgtPagesOH_13;
  wire [7:0] T_714;
  wire [5:0] tgtPagesOH_14;
  wire [7:0] T_716;
  wire [5:0] tgtPagesOH_15;
  wire [7:0] T_718;
  wire [5:0] tgtPagesOH_16;
  wire [7:0] T_720;
  wire [5:0] tgtPagesOH_17;
  wire [7:0] T_722;
  wire [5:0] tgtPagesOH_18;
  wire [7:0] T_724;
  wire [5:0] tgtPagesOH_19;
  wire [7:0] T_726;
  wire [5:0] tgtPagesOH_20;
  wire [7:0] T_728;
  wire [5:0] tgtPagesOH_21;
  wire [7:0] T_730;
  wire [5:0] tgtPagesOH_22;
  wire [7:0] T_732;
  wire [5:0] tgtPagesOH_23;
  wire [7:0] T_734;
  wire [5:0] tgtPagesOH_24;
  wire [7:0] T_736;
  wire [5:0] tgtPagesOH_25;
  wire [7:0] T_738;
  wire [5:0] tgtPagesOH_26;
  wire [7:0] T_740;
  wire [5:0] tgtPagesOH_27;
  wire [7:0] T_742;
  wire [5:0] tgtPagesOH_28;
  wire [7:0] T_744;
  wire [5:0] tgtPagesOH_29;
  wire [7:0] T_746;
  wire [5:0] tgtPagesOH_30;
  wire [7:0] T_748;
  wire [5:0] tgtPagesOH_31;
  wire [7:0] T_750;
  wire [5:0] tgtPagesOH_32;
  wire [7:0] T_752;
  wire [5:0] tgtPagesOH_33;
  wire [7:0] T_754;
  wire [5:0] tgtPagesOH_34;
  wire [7:0] T_756;
  wire [5:0] tgtPagesOH_35;
  wire [7:0] T_758;
  wire [5:0] tgtPagesOH_36;
  wire [7:0] T_760;
  wire [5:0] tgtPagesOH_37;
  wire [7:0] T_762;
  wire [5:0] tgtPagesOH_38;
  wire [7:0] T_764;
  wire [5:0] tgtPagesOH_39;
  reg [39:0] isValid;
  reg [63:0] GEN_641;
  reg [39:0] isReturn;
  reg [63:0] GEN_642;
  reg [39:0] isJump;
  reg [63:0] GEN_643;
  reg  brIdx_0;
  reg [31:0] GEN_644;
  reg  brIdx_1;
  reg [31:0] GEN_645;
  reg  brIdx_2;
  reg [31:0] GEN_646;
  reg  brIdx_3;
  reg [31:0] GEN_647;
  reg  brIdx_4;
  reg [31:0] GEN_648;
  reg  brIdx_5;
  reg [31:0] GEN_649;
  reg  brIdx_6;
  reg [31:0] GEN_650;
  reg  brIdx_7;
  reg [31:0] GEN_651;
  reg  brIdx_8;
  reg [31:0] GEN_652;
  reg  brIdx_9;
  reg [31:0] GEN_653;
  reg  brIdx_10;
  reg [31:0] GEN_654;
  reg  brIdx_11;
  reg [31:0] GEN_655;
  reg  brIdx_12;
  reg [31:0] GEN_656;
  reg  brIdx_13;
  reg [31:0] GEN_657;
  reg  brIdx_14;
  reg [31:0] GEN_658;
  reg  brIdx_15;
  reg [31:0] GEN_659;
  reg  brIdx_16;
  reg [31:0] GEN_660;
  reg  brIdx_17;
  reg [31:0] GEN_661;
  reg  brIdx_18;
  reg [31:0] GEN_662;
  reg  brIdx_19;
  reg [31:0] GEN_663;
  reg  brIdx_20;
  reg [31:0] GEN_664;
  reg  brIdx_21;
  reg [31:0] GEN_665;
  reg  brIdx_22;
  reg [31:0] GEN_666;
  reg  brIdx_23;
  reg [31:0] GEN_667;
  reg  brIdx_24;
  reg [31:0] GEN_668;
  reg  brIdx_25;
  reg [31:0] GEN_669;
  reg  brIdx_26;
  reg [31:0] GEN_670;
  reg  brIdx_27;
  reg [31:0] GEN_671;
  reg  brIdx_28;
  reg [31:0] GEN_672;
  reg  brIdx_29;
  reg [31:0] GEN_673;
  reg  brIdx_30;
  reg [31:0] GEN_674;
  reg  brIdx_31;
  reg [31:0] GEN_675;
  reg  brIdx_32;
  reg [31:0] GEN_676;
  reg  brIdx_33;
  reg [31:0] GEN_677;
  reg  brIdx_34;
  reg [31:0] GEN_678;
  reg  brIdx_35;
  reg [31:0] GEN_679;
  reg  brIdx_36;
  reg [31:0] GEN_680;
  reg  brIdx_37;
  reg [31:0] GEN_681;
  reg  brIdx_38;
  reg [31:0] GEN_682;
  reg  brIdx_39;
  reg [31:0] GEN_683;
  reg  T_777;
  reg [31:0] GEN_684;
  reg  T_778_prediction_valid;
  reg [31:0] GEN_685;
  reg  T_778_prediction_bits_taken;
  reg [31:0] GEN_686;
  reg [1:0] T_778_prediction_bits_mask;
  reg [31:0] GEN_687;
  reg  T_778_prediction_bits_bridx;
  reg [31:0] GEN_688;
  reg [38:0] T_778_prediction_bits_target;
  reg [63:0] GEN_689;
  reg [5:0] T_778_prediction_bits_entry;
  reg [31:0] GEN_690;
  reg [6:0] T_778_prediction_bits_bht_history;
  reg [31:0] GEN_691;
  reg [1:0] T_778_prediction_bits_bht_value;
  reg [31:0] GEN_692;
  reg [38:0] T_778_pc;
  reg [63:0] GEN_693;
  reg [38:0] T_778_target;
  reg [63:0] GEN_694;
  reg  T_778_taken;
  reg [31:0] GEN_695;
  reg  T_778_isValid;
  reg [31:0] GEN_696;
  reg  T_778_isJump;
  reg [31:0] GEN_697;
  reg  T_778_isReturn;
  reg [31:0] GEN_698;
  reg [38:0] T_778_br_pc;
  reg [63:0] GEN_699;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] GEN_9;
  wire  GEN_10;
  wire [38:0] GEN_11;
  wire [5:0] GEN_12;
  wire [6:0] GEN_13;
  wire [1:0] GEN_14;
  wire [38:0] GEN_15;
  wire [38:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [38:0] GEN_21;
  wire  r_btb_update_valid;
  wire  r_btb_update_bits_prediction_valid;
  wire  r_btb_update_bits_prediction_bits_taken;
  wire [1:0] r_btb_update_bits_prediction_bits_mask;
  wire  r_btb_update_bits_prediction_bits_bridx;
  wire [38:0] r_btb_update_bits_prediction_bits_target;
  wire [5:0] r_btb_update_bits_prediction_bits_entry;
  wire [6:0] r_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] r_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] r_btb_update_bits_pc;
  wire [38:0] r_btb_update_bits_target;
  wire  r_btb_update_bits_taken;
  wire  r_btb_update_bits_isValid;
  wire  r_btb_update_bits_isJump;
  wire  r_btb_update_bits_isReturn;
  wire [38:0] r_btb_update_bits_br_pc;
  wire [26:0] T_964;
  wire  T_965;
  wire  T_966;
  wire  T_967;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire [1:0] T_971;
  wire [2:0] T_972;
  wire [1:0] T_973;
  wire [2:0] T_974;
  wire [5:0] T_975;
  wire [5:0] pageHit;
  wire [10:0] T_976;
  wire  T_977;
  wire  T_979;
  wire  T_981;
  wire  T_983;
  wire  T_985;
  wire  T_987;
  wire  T_989;
  wire  T_991;
  wire  T_993;
  wire  T_995;
  wire  T_997;
  wire  T_999;
  wire  T_1001;
  wire  T_1003;
  wire  T_1005;
  wire  T_1007;
  wire  T_1009;
  wire  T_1011;
  wire  T_1013;
  wire  T_1015;
  wire  T_1017;
  wire  T_1019;
  wire  T_1021;
  wire  T_1023;
  wire  T_1025;
  wire  T_1027;
  wire  T_1029;
  wire  T_1031;
  wire  T_1033;
  wire  T_1035;
  wire  T_1037;
  wire  T_1039;
  wire  T_1041;
  wire  T_1043;
  wire  T_1045;
  wire  T_1047;
  wire  T_1049;
  wire  T_1051;
  wire  T_1053;
  wire  T_1055;
  wire [1:0] T_1056;
  wire [1:0] T_1057;
  wire [2:0] T_1058;
  wire [4:0] T_1059;
  wire [1:0] T_1060;
  wire [1:0] T_1061;
  wire [2:0] T_1062;
  wire [4:0] T_1063;
  wire [9:0] T_1064;
  wire [1:0] T_1065;
  wire [1:0] T_1066;
  wire [2:0] T_1067;
  wire [4:0] T_1068;
  wire [1:0] T_1069;
  wire [1:0] T_1070;
  wire [2:0] T_1071;
  wire [4:0] T_1072;
  wire [9:0] T_1073;
  wire [19:0] T_1074;
  wire [1:0] T_1075;
  wire [1:0] T_1076;
  wire [2:0] T_1077;
  wire [4:0] T_1078;
  wire [1:0] T_1079;
  wire [1:0] T_1080;
  wire [2:0] T_1081;
  wire [4:0] T_1082;
  wire [9:0] T_1083;
  wire [1:0] T_1084;
  wire [1:0] T_1085;
  wire [2:0] T_1086;
  wire [4:0] T_1087;
  wire [1:0] T_1088;
  wire [1:0] T_1089;
  wire [2:0] T_1090;
  wire [4:0] T_1091;
  wire [9:0] T_1092;
  wire [19:0] T_1093;
  wire [39:0] T_1094;
  wire [5:0] T_1095;
  wire [5:0] T_1096;
  wire [5:0] T_1097;
  wire [5:0] T_1098;
  wire [5:0] T_1099;
  wire [5:0] T_1100;
  wire [5:0] T_1101;
  wire [5:0] T_1102;
  wire [5:0] T_1103;
  wire [5:0] T_1104;
  wire [5:0] T_1105;
  wire [5:0] T_1106;
  wire [5:0] T_1107;
  wire [5:0] T_1108;
  wire [5:0] T_1109;
  wire [5:0] T_1110;
  wire [5:0] T_1111;
  wire [5:0] T_1112;
  wire [5:0] T_1113;
  wire [5:0] T_1114;
  wire [5:0] T_1115;
  wire [5:0] T_1116;
  wire [5:0] T_1117;
  wire [5:0] T_1118;
  wire [5:0] T_1119;
  wire [5:0] T_1120;
  wire [5:0] T_1121;
  wire [5:0] T_1122;
  wire [5:0] T_1123;
  wire [5:0] T_1124;
  wire [5:0] T_1125;
  wire [5:0] T_1126;
  wire [5:0] T_1127;
  wire [5:0] T_1128;
  wire [5:0] T_1129;
  wire [5:0] T_1130;
  wire [5:0] T_1131;
  wire [5:0] T_1132;
  wire [5:0] T_1133;
  wire [5:0] T_1134;
  wire  T_1136;
  wire  T_1138;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1146;
  wire  T_1148;
  wire  T_1150;
  wire  T_1152;
  wire  T_1154;
  wire  T_1156;
  wire  T_1158;
  wire  T_1160;
  wire  T_1162;
  wire  T_1164;
  wire  T_1166;
  wire  T_1168;
  wire  T_1170;
  wire  T_1172;
  wire  T_1174;
  wire  T_1176;
  wire  T_1178;
  wire  T_1180;
  wire  T_1182;
  wire  T_1184;
  wire  T_1186;
  wire  T_1188;
  wire  T_1190;
  wire  T_1192;
  wire  T_1194;
  wire  T_1196;
  wire  T_1198;
  wire  T_1200;
  wire  T_1202;
  wire  T_1204;
  wire  T_1206;
  wire  T_1208;
  wire  T_1210;
  wire  T_1212;
  wire  T_1214;
  wire [1:0] T_1215;
  wire [1:0] T_1216;
  wire [2:0] T_1217;
  wire [4:0] T_1218;
  wire [1:0] T_1219;
  wire [1:0] T_1220;
  wire [2:0] T_1221;
  wire [4:0] T_1222;
  wire [9:0] T_1223;
  wire [1:0] T_1224;
  wire [1:0] T_1225;
  wire [2:0] T_1226;
  wire [4:0] T_1227;
  wire [1:0] T_1228;
  wire [1:0] T_1229;
  wire [2:0] T_1230;
  wire [4:0] T_1231;
  wire [9:0] T_1232;
  wire [19:0] T_1233;
  wire [1:0] T_1234;
  wire [1:0] T_1235;
  wire [2:0] T_1236;
  wire [4:0] T_1237;
  wire [1:0] T_1238;
  wire [1:0] T_1239;
  wire [2:0] T_1240;
  wire [4:0] T_1241;
  wire [9:0] T_1242;
  wire [1:0] T_1243;
  wire [1:0] T_1244;
  wire [2:0] T_1245;
  wire [4:0] T_1246;
  wire [1:0] T_1247;
  wire [1:0] T_1248;
  wire [2:0] T_1249;
  wire [4:0] T_1250;
  wire [9:0] T_1251;
  wire [19:0] T_1252;
  wire [39:0] T_1253;
  wire [39:0] T_1254;
  wire [39:0] hitsVec;
  wire [26:0] T_1255;
  wire  T_1256;
  wire  T_1257;
  wire  T_1258;
  wire  T_1259;
  wire  T_1260;
  wire  T_1261;
  wire [1:0] T_1262;
  wire [2:0] T_1263;
  wire [1:0] T_1264;
  wire [2:0] T_1265;
  wire [5:0] T_1266;
  wire [5:0] updatePageHit;
  wire [10:0] T_1267;
  wire  T_1547;
  wire  T_1548;
  reg [5:0] nextRepl;
  reg [31:0] GEN_700;
  wire  T_1551;
  wire [6:0] T_1553;
  wire [5:0] T_1554;
  wire [5:0] GEN_22;
  wire [5:0] GEN_23;
  wire  useUpdatePageHit;
  wire  usePageHit;
  wire  doIdxPageRepl;
  reg [2:0] nextPageRepl;
  reg [31:0] GEN_701;
  wire [4:0] T_1561;
  wire  T_1562;
  wire [5:0] T_1563;
  wire [7:0] T_1565;
  wire [7:0] idxPageRepl;
  wire [7:0] idxPageUpdateOH;
  wire [3:0] T_1566;
  wire [3:0] T_1567;
  wire  T_1569;
  wire [3:0] T_1570;
  wire [1:0] T_1571;
  wire [1:0] T_1572;
  wire  T_1574;
  wire [1:0] T_1575;
  wire  T_1576;
  wire [1:0] T_1577;
  wire [2:0] idxPageUpdate;
  wire [7:0] idxPageReplEn;
  wire  samePage;
  wire  T_1582;
  wire  T_1584;
  wire  doTgtPageRepl;
  wire [4:0] T_1585;
  wire  T_1586;
  wire [5:0] T_1587;
  wire [7:0] tgtPageRepl;
  wire [7:0] T_1588;
  wire [3:0] T_1589;
  wire [3:0] T_1590;
  wire  T_1592;
  wire [3:0] T_1593;
  wire [1:0] T_1594;
  wire [1:0] T_1595;
  wire  T_1597;
  wire [1:0] T_1598;
  wire  T_1599;
  wire [1:0] T_1600;
  wire [2:0] tgtPageUpdate;
  wire [7:0] tgtPageReplEn;
  wire  T_1602;
  wire  T_1603;
  wire  T_1604;
  wire [1:0] T_1607;
  wire [2:0] GEN_478;
  wire [3:0] T_1608;
  wire [2:0] T_1609;
  wire  T_1611;
  wire  T_1612;
  wire [2:0] T_1614;
  wire [2:0] GEN_24;
  wire [5:0] T_1615;
  wire [63:0] T_1617;
  wire [10:0] GEN_0;
  wire [10:0] GEN_25;
  wire [10:0] GEN_26;
  wire [10:0] GEN_27;
  wire [10:0] GEN_28;
  wire [10:0] GEN_29;
  wire [10:0] GEN_30;
  wire [10:0] GEN_31;
  wire [10:0] GEN_32;
  wire [10:0] GEN_33;
  wire [10:0] GEN_34;
  wire [10:0] GEN_35;
  wire [10:0] GEN_36;
  wire [10:0] GEN_37;
  wire [10:0] GEN_38;
  wire [10:0] GEN_39;
  wire [10:0] GEN_40;
  wire [10:0] GEN_41;
  wire [10:0] GEN_42;
  wire [10:0] GEN_43;
  wire [10:0] GEN_44;
  wire [10:0] GEN_45;
  wire [10:0] GEN_46;
  wire [10:0] GEN_47;
  wire [10:0] GEN_48;
  wire [10:0] GEN_49;
  wire [10:0] GEN_50;
  wire [10:0] GEN_51;
  wire [10:0] GEN_52;
  wire [10:0] GEN_53;
  wire [10:0] GEN_54;
  wire [10:0] GEN_55;
  wire [10:0] GEN_56;
  wire [10:0] GEN_57;
  wire [10:0] GEN_58;
  wire [10:0] GEN_59;
  wire [10:0] GEN_60;
  wire [10:0] GEN_61;
  wire [10:0] GEN_62;
  wire [10:0] GEN_63;
  wire [10:0] GEN_64;
  wire [10:0] GEN_1;
  wire [10:0] GEN_65;
  wire [10:0] GEN_66;
  wire [10:0] GEN_67;
  wire [10:0] GEN_68;
  wire [10:0] GEN_69;
  wire [10:0] GEN_70;
  wire [10:0] GEN_71;
  wire [10:0] GEN_72;
  wire [10:0] GEN_73;
  wire [10:0] GEN_74;
  wire [10:0] GEN_75;
  wire [10:0] GEN_76;
  wire [10:0] GEN_77;
  wire [10:0] GEN_78;
  wire [10:0] GEN_79;
  wire [10:0] GEN_80;
  wire [10:0] GEN_81;
  wire [10:0] GEN_82;
  wire [10:0] GEN_83;
  wire [10:0] GEN_84;
  wire [10:0] GEN_85;
  wire [10:0] GEN_86;
  wire [10:0] GEN_87;
  wire [10:0] GEN_88;
  wire [10:0] GEN_89;
  wire [10:0] GEN_90;
  wire [10:0] GEN_91;
  wire [10:0] GEN_92;
  wire [10:0] GEN_93;
  wire [10:0] GEN_94;
  wire [10:0] GEN_95;
  wire [10:0] GEN_96;
  wire [10:0] GEN_97;
  wire [10:0] GEN_98;
  wire [10:0] GEN_99;
  wire [10:0] GEN_100;
  wire [10:0] GEN_101;
  wire [10:0] GEN_102;
  wire [10:0] GEN_103;
  wire [10:0] GEN_104;
  wire [2:0] GEN_2;
  wire [2:0] GEN_105;
  wire [2:0] GEN_106;
  wire [2:0] GEN_107;
  wire [2:0] GEN_108;
  wire [2:0] GEN_109;
  wire [2:0] GEN_110;
  wire [2:0] GEN_111;
  wire [2:0] GEN_112;
  wire [2:0] GEN_113;
  wire [2:0] GEN_114;
  wire [2:0] GEN_115;
  wire [2:0] GEN_116;
  wire [2:0] GEN_117;
  wire [2:0] GEN_118;
  wire [2:0] GEN_119;
  wire [2:0] GEN_120;
  wire [2:0] GEN_121;
  wire [2:0] GEN_122;
  wire [2:0] GEN_123;
  wire [2:0] GEN_124;
  wire [2:0] GEN_125;
  wire [2:0] GEN_126;
  wire [2:0] GEN_127;
  wire [2:0] GEN_128;
  wire [2:0] GEN_129;
  wire [2:0] GEN_130;
  wire [2:0] GEN_131;
  wire [2:0] GEN_132;
  wire [2:0] GEN_133;
  wire [2:0] GEN_134;
  wire [2:0] GEN_135;
  wire [2:0] GEN_136;
  wire [2:0] GEN_137;
  wire [2:0] GEN_138;
  wire [2:0] GEN_139;
  wire [2:0] GEN_140;
  wire [2:0] GEN_141;
  wire [2:0] GEN_142;
  wire [2:0] GEN_143;
  wire [2:0] GEN_144;
  wire [2:0] GEN_3;
  wire [2:0] GEN_145;
  wire [2:0] GEN_146;
  wire [2:0] GEN_147;
  wire [2:0] GEN_148;
  wire [2:0] GEN_149;
  wire [2:0] GEN_150;
  wire [2:0] GEN_151;
  wire [2:0] GEN_152;
  wire [2:0] GEN_153;
  wire [2:0] GEN_154;
  wire [2:0] GEN_155;
  wire [2:0] GEN_156;
  wire [2:0] GEN_157;
  wire [2:0] GEN_158;
  wire [2:0] GEN_159;
  wire [2:0] GEN_160;
  wire [2:0] GEN_161;
  wire [2:0] GEN_162;
  wire [2:0] GEN_163;
  wire [2:0] GEN_164;
  wire [2:0] GEN_165;
  wire [2:0] GEN_166;
  wire [2:0] GEN_167;
  wire [2:0] GEN_168;
  wire [2:0] GEN_169;
  wire [2:0] GEN_170;
  wire [2:0] GEN_171;
  wire [2:0] GEN_172;
  wire [2:0] GEN_173;
  wire [2:0] GEN_174;
  wire [2:0] GEN_175;
  wire [2:0] GEN_176;
  wire [2:0] GEN_177;
  wire [2:0] GEN_178;
  wire [2:0] GEN_179;
  wire [2:0] GEN_180;
  wire [2:0] GEN_181;
  wire [2:0] GEN_182;
  wire [2:0] GEN_183;
  wire [2:0] GEN_184;
  wire [63:0] GEN_479;
  wire [63:0] T_1620;
  wire [63:0] T_1621;
  wire [63:0] T_1622;
  wire [63:0] T_1623;
  wire [63:0] GEN_481;
  wire [63:0] T_1624;
  wire [63:0] T_1626;
  wire [63:0] T_1627;
  wire [63:0] GEN_483;
  wire [63:0] T_1628;
  wire [63:0] T_1630;
  wire [63:0] T_1631;
  wire [37:0] T_1632;
  wire  GEN_4;
  wire  GEN_185;
  wire  GEN_186;
  wire  GEN_187;
  wire  GEN_188;
  wire  GEN_189;
  wire  GEN_190;
  wire  GEN_191;
  wire  GEN_192;
  wire  GEN_193;
  wire  GEN_194;
  wire  GEN_195;
  wire  GEN_196;
  wire  GEN_197;
  wire  GEN_198;
  wire  GEN_199;
  wire  GEN_200;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  T_1633;
  wire  T_1635;
  wire [7:0] T_1636;
  wire [26:0] T_1639;
  wire  T_1640;
  wire [26:0] GEN_225;
  wire  T_1641;
  wire [26:0] GEN_226;
  wire  T_1642;
  wire [26:0] GEN_227;
  wire [7:0] T_1643;
  wire [26:0] T_1646;
  wire  T_1647;
  wire [26:0] GEN_228;
  wire  T_1648;
  wire [26:0] GEN_229;
  wire  T_1649;
  wire [26:0] GEN_230;
  wire [7:0] GEN_485;
  wire [7:0] T_1650;
  wire [7:0] T_1651;
  wire [10:0] GEN_232;
  wire [10:0] GEN_233;
  wire [10:0] GEN_234;
  wire [10:0] GEN_235;
  wire [10:0] GEN_236;
  wire [10:0] GEN_237;
  wire [10:0] GEN_238;
  wire [10:0] GEN_239;
  wire [10:0] GEN_240;
  wire [10:0] GEN_241;
  wire [10:0] GEN_242;
  wire [10:0] GEN_243;
  wire [10:0] GEN_244;
  wire [10:0] GEN_245;
  wire [10:0] GEN_246;
  wire [10:0] GEN_247;
  wire [10:0] GEN_248;
  wire [10:0] GEN_249;
  wire [10:0] GEN_250;
  wire [10:0] GEN_251;
  wire [10:0] GEN_252;
  wire [10:0] GEN_253;
  wire [10:0] GEN_254;
  wire [10:0] GEN_255;
  wire [10:0] GEN_256;
  wire [10:0] GEN_257;
  wire [10:0] GEN_258;
  wire [10:0] GEN_259;
  wire [10:0] GEN_260;
  wire [10:0] GEN_261;
  wire [10:0] GEN_262;
  wire [10:0] GEN_263;
  wire [10:0] GEN_264;
  wire [10:0] GEN_265;
  wire [10:0] GEN_266;
  wire [10:0] GEN_267;
  wire [10:0] GEN_268;
  wire [10:0] GEN_269;
  wire [10:0] GEN_270;
  wire [10:0] GEN_271;
  wire [10:0] GEN_273;
  wire [10:0] GEN_274;
  wire [10:0] GEN_275;
  wire [10:0] GEN_276;
  wire [10:0] GEN_277;
  wire [10:0] GEN_278;
  wire [10:0] GEN_279;
  wire [10:0] GEN_280;
  wire [10:0] GEN_281;
  wire [10:0] GEN_282;
  wire [10:0] GEN_283;
  wire [10:0] GEN_284;
  wire [10:0] GEN_285;
  wire [10:0] GEN_286;
  wire [10:0] GEN_287;
  wire [10:0] GEN_288;
  wire [10:0] GEN_289;
  wire [10:0] GEN_290;
  wire [10:0] GEN_291;
  wire [10:0] GEN_292;
  wire [10:0] GEN_293;
  wire [10:0] GEN_294;
  wire [10:0] GEN_295;
  wire [10:0] GEN_296;
  wire [10:0] GEN_297;
  wire [10:0] GEN_298;
  wire [10:0] GEN_299;
  wire [10:0] GEN_300;
  wire [10:0] GEN_301;
  wire [10:0] GEN_302;
  wire [10:0] GEN_303;
  wire [10:0] GEN_304;
  wire [10:0] GEN_305;
  wire [10:0] GEN_306;
  wire [10:0] GEN_307;
  wire [10:0] GEN_308;
  wire [10:0] GEN_309;
  wire [10:0] GEN_310;
  wire [10:0] GEN_311;
  wire [10:0] GEN_312;
  wire [2:0] GEN_314;
  wire [2:0] GEN_315;
  wire [2:0] GEN_316;
  wire [2:0] GEN_317;
  wire [2:0] GEN_318;
  wire [2:0] GEN_319;
  wire [2:0] GEN_320;
  wire [2:0] GEN_321;
  wire [2:0] GEN_322;
  wire [2:0] GEN_323;
  wire [2:0] GEN_324;
  wire [2:0] GEN_325;
  wire [2:0] GEN_326;
  wire [2:0] GEN_327;
  wire [2:0] GEN_328;
  wire [2:0] GEN_329;
  wire [2:0] GEN_330;
  wire [2:0] GEN_331;
  wire [2:0] GEN_332;
  wire [2:0] GEN_333;
  wire [2:0] GEN_334;
  wire [2:0] GEN_335;
  wire [2:0] GEN_336;
  wire [2:0] GEN_337;
  wire [2:0] GEN_338;
  wire [2:0] GEN_339;
  wire [2:0] GEN_340;
  wire [2:0] GEN_341;
  wire [2:0] GEN_342;
  wire [2:0] GEN_343;
  wire [2:0] GEN_344;
  wire [2:0] GEN_345;
  wire [2:0] GEN_346;
  wire [2:0] GEN_347;
  wire [2:0] GEN_348;
  wire [2:0] GEN_349;
  wire [2:0] GEN_350;
  wire [2:0] GEN_351;
  wire [2:0] GEN_352;
  wire [2:0] GEN_353;
  wire [2:0] GEN_355;
  wire [2:0] GEN_356;
  wire [2:0] GEN_357;
  wire [2:0] GEN_358;
  wire [2:0] GEN_359;
  wire [2:0] GEN_360;
  wire [2:0] GEN_361;
  wire [2:0] GEN_362;
  wire [2:0] GEN_363;
  wire [2:0] GEN_364;
  wire [2:0] GEN_365;
  wire [2:0] GEN_366;
  wire [2:0] GEN_367;
  wire [2:0] GEN_368;
  wire [2:0] GEN_369;
  wire [2:0] GEN_370;
  wire [2:0] GEN_371;
  wire [2:0] GEN_372;
  wire [2:0] GEN_373;
  wire [2:0] GEN_374;
  wire [2:0] GEN_375;
  wire [2:0] GEN_376;
  wire [2:0] GEN_377;
  wire [2:0] GEN_378;
  wire [2:0] GEN_379;
  wire [2:0] GEN_380;
  wire [2:0] GEN_381;
  wire [2:0] GEN_382;
  wire [2:0] GEN_383;
  wire [2:0] GEN_384;
  wire [2:0] GEN_385;
  wire [2:0] GEN_386;
  wire [2:0] GEN_387;
  wire [2:0] GEN_388;
  wire [2:0] GEN_389;
  wire [2:0] GEN_390;
  wire [2:0] GEN_391;
  wire [2:0] GEN_392;
  wire [2:0] GEN_393;
  wire [2:0] GEN_394;
  wire [63:0] GEN_395;
  wire [63:0] GEN_396;
  wire [63:0] GEN_397;
  wire  GEN_399;
  wire  GEN_400;
  wire  GEN_401;
  wire  GEN_402;
  wire  GEN_403;
  wire  GEN_404;
  wire  GEN_405;
  wire  GEN_406;
  wire  GEN_407;
  wire  GEN_408;
  wire  GEN_409;
  wire  GEN_410;
  wire  GEN_411;
  wire  GEN_412;
  wire  GEN_413;
  wire  GEN_414;
  wire  GEN_415;
  wire  GEN_416;
  wire  GEN_417;
  wire  GEN_418;
  wire  GEN_419;
  wire  GEN_420;
  wire  GEN_421;
  wire  GEN_422;
  wire  GEN_423;
  wire  GEN_424;
  wire  GEN_425;
  wire  GEN_426;
  wire  GEN_427;
  wire  GEN_428;
  wire  GEN_429;
  wire  GEN_430;
  wire  GEN_431;
  wire  GEN_432;
  wire  GEN_433;
  wire  GEN_434;
  wire  GEN_435;
  wire  GEN_436;
  wire  GEN_437;
  wire  GEN_438;
  wire [26:0] GEN_439;
  wire [26:0] GEN_440;
  wire [26:0] GEN_441;
  wire [26:0] GEN_442;
  wire [26:0] GEN_443;
  wire [26:0] GEN_444;
  wire [7:0] GEN_445;
  wire  T_1653;
  wire  T_1655;
  wire  T_1656;
  wire  T_1657;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1662;
  wire  T_1663;
  wire  T_1664;
  wire  T_1665;
  wire  T_1666;
  wire  T_1667;
  wire  T_1668;
  wire  T_1669;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1673;
  wire  T_1674;
  wire  T_1675;
  wire  T_1676;
  wire  T_1677;
  wire  T_1678;
  wire  T_1679;
  wire  T_1680;
  wire  T_1681;
  wire  T_1682;
  wire  T_1683;
  wire  T_1684;
  wire  T_1685;
  wire  T_1686;
  wire  T_1687;
  wire  T_1688;
  wire  T_1689;
  wire  T_1690;
  wire  T_1691;
  wire  T_1692;
  wire  T_1693;
  wire  T_1694;
  wire [5:0] T_1696;
  wire [5:0] T_1698;
  wire [5:0] T_1700;
  wire [5:0] T_1702;
  wire [5:0] T_1704;
  wire [5:0] T_1706;
  wire [5:0] T_1708;
  wire [5:0] T_1710;
  wire [5:0] T_1712;
  wire [5:0] T_1714;
  wire [5:0] T_1716;
  wire [5:0] T_1718;
  wire [5:0] T_1720;
  wire [5:0] T_1722;
  wire [5:0] T_1724;
  wire [5:0] T_1726;
  wire [5:0] T_1728;
  wire [5:0] T_1730;
  wire [5:0] T_1732;
  wire [5:0] T_1734;
  wire [5:0] T_1736;
  wire [5:0] T_1738;
  wire [5:0] T_1740;
  wire [5:0] T_1742;
  wire [5:0] T_1744;
  wire [5:0] T_1746;
  wire [5:0] T_1748;
  wire [5:0] T_1750;
  wire [5:0] T_1752;
  wire [5:0] T_1754;
  wire [5:0] T_1756;
  wire [5:0] T_1758;
  wire [5:0] T_1760;
  wire [5:0] T_1762;
  wire [5:0] T_1764;
  wire [5:0] T_1766;
  wire [5:0] T_1768;
  wire [5:0] T_1770;
  wire [5:0] T_1772;
  wire [5:0] T_1774;
  wire [5:0] T_1776;
  wire [5:0] T_1777;
  wire [5:0] T_1778;
  wire [5:0] T_1779;
  wire [5:0] T_1780;
  wire [5:0] T_1781;
  wire [5:0] T_1782;
  wire [5:0] T_1783;
  wire [5:0] T_1784;
  wire [5:0] T_1785;
  wire [5:0] T_1786;
  wire [5:0] T_1787;
  wire [5:0] T_1788;
  wire [5:0] T_1789;
  wire [5:0] T_1790;
  wire [5:0] T_1791;
  wire [5:0] T_1792;
  wire [5:0] T_1793;
  wire [5:0] T_1794;
  wire [5:0] T_1795;
  wire [5:0] T_1796;
  wire [5:0] T_1797;
  wire [5:0] T_1798;
  wire [5:0] T_1799;
  wire [5:0] T_1800;
  wire [5:0] T_1801;
  wire [5:0] T_1802;
  wire [5:0] T_1803;
  wire [5:0] T_1804;
  wire [5:0] T_1805;
  wire [5:0] T_1806;
  wire [5:0] T_1807;
  wire [5:0] T_1808;
  wire [5:0] T_1809;
  wire [5:0] T_1810;
  wire [5:0] T_1811;
  wire [5:0] T_1812;
  wire [5:0] T_1813;
  wire [5:0] T_1814;
  wire [5:0] T_1815;
  wire  T_1816;
  wire  T_1817;
  wire  T_1818;
  wire  T_1819;
  wire  T_1820;
  wire  T_1821;
  wire [26:0] T_1823;
  wire [26:0] T_1825;
  wire [26:0] T_1827;
  wire [26:0] T_1829;
  wire [26:0] T_1831;
  wire [26:0] T_1833;
  wire [26:0] T_1835;
  wire [26:0] T_1836;
  wire [26:0] T_1837;
  wire [26:0] T_1838;
  wire [26:0] T_1839;
  wire [26:0] T_1840;
  wire [10:0] T_1882;
  wire [10:0] T_1884;
  wire [10:0] T_1886;
  wire [10:0] T_1888;
  wire [10:0] T_1890;
  wire [10:0] T_1892;
  wire [10:0] T_1894;
  wire [10:0] T_1896;
  wire [10:0] T_1898;
  wire [10:0] T_1900;
  wire [10:0] T_1902;
  wire [10:0] T_1904;
  wire [10:0] T_1906;
  wire [10:0] T_1908;
  wire [10:0] T_1910;
  wire [10:0] T_1912;
  wire [10:0] T_1914;
  wire [10:0] T_1916;
  wire [10:0] T_1918;
  wire [10:0] T_1920;
  wire [10:0] T_1922;
  wire [10:0] T_1924;
  wire [10:0] T_1926;
  wire [10:0] T_1928;
  wire [10:0] T_1930;
  wire [10:0] T_1932;
  wire [10:0] T_1934;
  wire [10:0] T_1936;
  wire [10:0] T_1938;
  wire [10:0] T_1940;
  wire [10:0] T_1942;
  wire [10:0] T_1944;
  wire [10:0] T_1946;
  wire [10:0] T_1948;
  wire [10:0] T_1950;
  wire [10:0] T_1952;
  wire [10:0] T_1954;
  wire [10:0] T_1956;
  wire [10:0] T_1958;
  wire [10:0] T_1960;
  wire [10:0] T_1962;
  wire [10:0] T_1963;
  wire [10:0] T_1964;
  wire [10:0] T_1965;
  wire [10:0] T_1966;
  wire [10:0] T_1967;
  wire [10:0] T_1968;
  wire [10:0] T_1969;
  wire [10:0] T_1970;
  wire [10:0] T_1971;
  wire [10:0] T_1972;
  wire [10:0] T_1973;
  wire [10:0] T_1974;
  wire [10:0] T_1975;
  wire [10:0] T_1976;
  wire [10:0] T_1977;
  wire [10:0] T_1978;
  wire [10:0] T_1979;
  wire [10:0] T_1980;
  wire [10:0] T_1981;
  wire [10:0] T_1982;
  wire [10:0] T_1983;
  wire [10:0] T_1984;
  wire [10:0] T_1985;
  wire [10:0] T_1986;
  wire [10:0] T_1987;
  wire [10:0] T_1988;
  wire [10:0] T_1989;
  wire [10:0] T_1990;
  wire [10:0] T_1991;
  wire [10:0] T_1992;
  wire [10:0] T_1993;
  wire [10:0] T_1994;
  wire [10:0] T_1995;
  wire [10:0] T_1996;
  wire [10:0] T_1997;
  wire [10:0] T_1998;
  wire [10:0] T_1999;
  wire [10:0] T_2000;
  wire [10:0] T_2001;
  wire [11:0] GEN_486;
  wire [11:0] T_2002;
  wire [38:0] T_2003;
  wire [7:0] T_2004;
  wire [31:0] T_2005;
  wire  T_2007;
  wire [31:0] GEN_487;
  wire [31:0] T_2008;
  wire [15:0] T_2009;
  wire [15:0] T_2010;
  wire  T_2012;
  wire [15:0] T_2013;
  wire [7:0] T_2014;
  wire [7:0] T_2015;
  wire  T_2017;
  wire [7:0] T_2018;
  wire [3:0] T_2019;
  wire [3:0] T_2020;
  wire  T_2022;
  wire [3:0] T_2023;
  wire [1:0] T_2024;
  wire [1:0] T_2025;
  wire  T_2027;
  wire [1:0] T_2028;
  wire  T_2029;
  wire [1:0] T_2030;
  wire [2:0] T_2031;
  wire [3:0] T_2032;
  wire [4:0] T_2033;
  wire [5:0] T_2034;
  wire  T_2076;
  wire  T_2078;
  wire  T_2080;
  wire  T_2082;
  wire  T_2084;
  wire  T_2086;
  wire  T_2088;
  wire  T_2090;
  wire  T_2092;
  wire  T_2094;
  wire  T_2096;
  wire  T_2098;
  wire  T_2100;
  wire  T_2102;
  wire  T_2104;
  wire  T_2106;
  wire  T_2108;
  wire  T_2110;
  wire  T_2112;
  wire  T_2114;
  wire  T_2116;
  wire  T_2118;
  wire  T_2120;
  wire  T_2122;
  wire  T_2124;
  wire  T_2126;
  wire  T_2128;
  wire  T_2130;
  wire  T_2132;
  wire  T_2134;
  wire  T_2136;
  wire  T_2138;
  wire  T_2140;
  wire  T_2142;
  wire  T_2144;
  wire  T_2146;
  wire  T_2148;
  wire  T_2150;
  wire  T_2152;
  wire  T_2154;
  wire  T_2156;
  wire  T_2157;
  wire  T_2158;
  wire  T_2159;
  wire  T_2160;
  wire  T_2161;
  wire  T_2162;
  wire  T_2163;
  wire  T_2164;
  wire  T_2165;
  wire  T_2166;
  wire  T_2167;
  wire  T_2168;
  wire  T_2169;
  wire  T_2170;
  wire  T_2171;
  wire  T_2172;
  wire  T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2176;
  wire  T_2177;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire  T_2182;
  wire  T_2183;
  wire  T_2184;
  wire  T_2185;
  wire  T_2186;
  wire  T_2187;
  wire  T_2188;
  wire  T_2189;
  wire  T_2190;
  wire  T_2191;
  wire  T_2192;
  wire  T_2193;
  wire  T_2194;
  wire  T_2195;
  wire  T_2197;
  wire  T_2199;
  wire  T_2200;
  wire [1:0] T_2201;
  wire [2:0] T_2203;
  wire [1:0] T_2204;
  wire [2:0] T_2206;
  reg [1:0] T_2209 [0:127];
  reg [31:0] GEN_702;
  wire [1:0] T_2209_T_2227_data;
  wire [6:0] T_2209_T_2227_addr;
  wire  T_2209_T_2227_en;
  wire [1:0] T_2209_T_2234_data;
  wire [6:0] T_2209_T_2234_addr;
  wire  T_2209_T_2234_mask;
  wire  T_2209_T_2234_en;
  reg [6:0] T_2211;
  reg [31:0] GEN_703;
  wire [39:0] T_2212;
  wire  T_2214;
  wire  T_2216;
  wire  T_2217;
  wire  T_2218;
  wire [6:0] T_2222_history;
  wire [1:0] T_2222_value;
  wire [7:0] T_2225;
  wire [7:0] GEN_488;
  wire [7:0] T_2226;
  wire  T_2228;
  wire [5:0] T_2229;
  wire [6:0] T_2230;
  wire [6:0] GEN_446;
  wire  T_2231;
  wire [7:0] T_2232;
  wire [7:0] GEN_489;
  wire [7:0] T_2233;
  wire  T_2235;
  wire  T_2236;
  wire  T_2237;
  wire  T_2240;
  wire  T_2241;
  wire  T_2242;
  wire [1:0] T_2243;
  wire [5:0] T_2244;
  wire [6:0] T_2245;
  wire [6:0] GEN_447;
  wire [6:0] GEN_453;
  wire  T_2248;
  wire  T_2249;
  wire  GEN_454;
  reg [1:0] T_2252;
  reg [31:0] GEN_704;
  reg  T_2254;
  reg [31:0] GEN_705;
  reg [38:0] T_2261_0;
  reg [63:0] GEN_706;
  reg [38:0] T_2261_1;
  reg [63:0] GEN_707;
  wire [39:0] T_2263;
  wire  T_2265;
  wire  T_2267;
  wire  T_2269;
  wire  T_2270;
  wire [38:0] GEN_5;
  wire [38:0] GEN_455;
  wire [38:0] GEN_457;
  wire  T_2272;
  wire [2:0] T_2274;
  wire [1:0] T_2275;
  wire [1:0] GEN_458;
  wire [1:0] T_2281;
  wire  T_2282;
  wire [38:0] GEN_6;
  wire [38:0] GEN_459;
  wire [38:0] GEN_460;
  wire [38:0] GEN_461;
  wire [1:0] GEN_462;
  wire [38:0] GEN_464;
  wire [38:0] GEN_465;
  wire  GEN_466;
  wire [38:0] GEN_467;
  wire  T_2285;
  wire  T_2287;
  wire  T_2288;
  wire [2:0] T_2294;
  wire [1:0] T_2295;
  wire [1:0] T_2301;
  wire  T_2302;
  wire [1:0] GEN_468;
  wire  GEN_469;
  wire [1:0] GEN_470;
  wire  GEN_471;
  wire [1:0] GEN_472;
  wire [38:0] GEN_474;
  wire [38:0] GEN_475;
  wire  GEN_476;
  wire [38:0] GEN_477;
  assign io_resp_valid = T_1653;
  assign io_resp_bits_taken = GEN_454;
  assign io_resp_bits_mask = T_2206[1:0];
  assign io_resp_bits_bridx = T_2195;
  assign io_resp_bits_target = GEN_477;
  assign io_resp_bits_entry = T_2034;
  assign io_resp_bits_bht_history = T_2222_history;
  assign io_resp_bits_bht_value = T_2222_value;
  assign T_606 = 8'h1 << idxPages_0;
  assign idxPagesOH_0 = T_606[5:0];
  assign T_608 = 8'h1 << idxPages_1;
  assign idxPagesOH_1 = T_608[5:0];
  assign T_610 = 8'h1 << idxPages_2;
  assign idxPagesOH_2 = T_610[5:0];
  assign T_612 = 8'h1 << idxPages_3;
  assign idxPagesOH_3 = T_612[5:0];
  assign T_614 = 8'h1 << idxPages_4;
  assign idxPagesOH_4 = T_614[5:0];
  assign T_616 = 8'h1 << idxPages_5;
  assign idxPagesOH_5 = T_616[5:0];
  assign T_618 = 8'h1 << idxPages_6;
  assign idxPagesOH_6 = T_618[5:0];
  assign T_620 = 8'h1 << idxPages_7;
  assign idxPagesOH_7 = T_620[5:0];
  assign T_622 = 8'h1 << idxPages_8;
  assign idxPagesOH_8 = T_622[5:0];
  assign T_624 = 8'h1 << idxPages_9;
  assign idxPagesOH_9 = T_624[5:0];
  assign T_626 = 8'h1 << idxPages_10;
  assign idxPagesOH_10 = T_626[5:0];
  assign T_628 = 8'h1 << idxPages_11;
  assign idxPagesOH_11 = T_628[5:0];
  assign T_630 = 8'h1 << idxPages_12;
  assign idxPagesOH_12 = T_630[5:0];
  assign T_632 = 8'h1 << idxPages_13;
  assign idxPagesOH_13 = T_632[5:0];
  assign T_634 = 8'h1 << idxPages_14;
  assign idxPagesOH_14 = T_634[5:0];
  assign T_636 = 8'h1 << idxPages_15;
  assign idxPagesOH_15 = T_636[5:0];
  assign T_638 = 8'h1 << idxPages_16;
  assign idxPagesOH_16 = T_638[5:0];
  assign T_640 = 8'h1 << idxPages_17;
  assign idxPagesOH_17 = T_640[5:0];
  assign T_642 = 8'h1 << idxPages_18;
  assign idxPagesOH_18 = T_642[5:0];
  assign T_644 = 8'h1 << idxPages_19;
  assign idxPagesOH_19 = T_644[5:0];
  assign T_646 = 8'h1 << idxPages_20;
  assign idxPagesOH_20 = T_646[5:0];
  assign T_648 = 8'h1 << idxPages_21;
  assign idxPagesOH_21 = T_648[5:0];
  assign T_650 = 8'h1 << idxPages_22;
  assign idxPagesOH_22 = T_650[5:0];
  assign T_652 = 8'h1 << idxPages_23;
  assign idxPagesOH_23 = T_652[5:0];
  assign T_654 = 8'h1 << idxPages_24;
  assign idxPagesOH_24 = T_654[5:0];
  assign T_656 = 8'h1 << idxPages_25;
  assign idxPagesOH_25 = T_656[5:0];
  assign T_658 = 8'h1 << idxPages_26;
  assign idxPagesOH_26 = T_658[5:0];
  assign T_660 = 8'h1 << idxPages_27;
  assign idxPagesOH_27 = T_660[5:0];
  assign T_662 = 8'h1 << idxPages_28;
  assign idxPagesOH_28 = T_662[5:0];
  assign T_664 = 8'h1 << idxPages_29;
  assign idxPagesOH_29 = T_664[5:0];
  assign T_666 = 8'h1 << idxPages_30;
  assign idxPagesOH_30 = T_666[5:0];
  assign T_668 = 8'h1 << idxPages_31;
  assign idxPagesOH_31 = T_668[5:0];
  assign T_670 = 8'h1 << idxPages_32;
  assign idxPagesOH_32 = T_670[5:0];
  assign T_672 = 8'h1 << idxPages_33;
  assign idxPagesOH_33 = T_672[5:0];
  assign T_674 = 8'h1 << idxPages_34;
  assign idxPagesOH_34 = T_674[5:0];
  assign T_676 = 8'h1 << idxPages_35;
  assign idxPagesOH_35 = T_676[5:0];
  assign T_678 = 8'h1 << idxPages_36;
  assign idxPagesOH_36 = T_678[5:0];
  assign T_680 = 8'h1 << idxPages_37;
  assign idxPagesOH_37 = T_680[5:0];
  assign T_682 = 8'h1 << idxPages_38;
  assign idxPagesOH_38 = T_682[5:0];
  assign T_684 = 8'h1 << idxPages_39;
  assign idxPagesOH_39 = T_684[5:0];
  assign T_686 = 8'h1 << tgtPages_0;
  assign tgtPagesOH_0 = T_686[5:0];
  assign T_688 = 8'h1 << tgtPages_1;
  assign tgtPagesOH_1 = T_688[5:0];
  assign T_690 = 8'h1 << tgtPages_2;
  assign tgtPagesOH_2 = T_690[5:0];
  assign T_692 = 8'h1 << tgtPages_3;
  assign tgtPagesOH_3 = T_692[5:0];
  assign T_694 = 8'h1 << tgtPages_4;
  assign tgtPagesOH_4 = T_694[5:0];
  assign T_696 = 8'h1 << tgtPages_5;
  assign tgtPagesOH_5 = T_696[5:0];
  assign T_698 = 8'h1 << tgtPages_6;
  assign tgtPagesOH_6 = T_698[5:0];
  assign T_700 = 8'h1 << tgtPages_7;
  assign tgtPagesOH_7 = T_700[5:0];
  assign T_702 = 8'h1 << tgtPages_8;
  assign tgtPagesOH_8 = T_702[5:0];
  assign T_704 = 8'h1 << tgtPages_9;
  assign tgtPagesOH_9 = T_704[5:0];
  assign T_706 = 8'h1 << tgtPages_10;
  assign tgtPagesOH_10 = T_706[5:0];
  assign T_708 = 8'h1 << tgtPages_11;
  assign tgtPagesOH_11 = T_708[5:0];
  assign T_710 = 8'h1 << tgtPages_12;
  assign tgtPagesOH_12 = T_710[5:0];
  assign T_712 = 8'h1 << tgtPages_13;
  assign tgtPagesOH_13 = T_712[5:0];
  assign T_714 = 8'h1 << tgtPages_14;
  assign tgtPagesOH_14 = T_714[5:0];
  assign T_716 = 8'h1 << tgtPages_15;
  assign tgtPagesOH_15 = T_716[5:0];
  assign T_718 = 8'h1 << tgtPages_16;
  assign tgtPagesOH_16 = T_718[5:0];
  assign T_720 = 8'h1 << tgtPages_17;
  assign tgtPagesOH_17 = T_720[5:0];
  assign T_722 = 8'h1 << tgtPages_18;
  assign tgtPagesOH_18 = T_722[5:0];
  assign T_724 = 8'h1 << tgtPages_19;
  assign tgtPagesOH_19 = T_724[5:0];
  assign T_726 = 8'h1 << tgtPages_20;
  assign tgtPagesOH_20 = T_726[5:0];
  assign T_728 = 8'h1 << tgtPages_21;
  assign tgtPagesOH_21 = T_728[5:0];
  assign T_730 = 8'h1 << tgtPages_22;
  assign tgtPagesOH_22 = T_730[5:0];
  assign T_732 = 8'h1 << tgtPages_23;
  assign tgtPagesOH_23 = T_732[5:0];
  assign T_734 = 8'h1 << tgtPages_24;
  assign tgtPagesOH_24 = T_734[5:0];
  assign T_736 = 8'h1 << tgtPages_25;
  assign tgtPagesOH_25 = T_736[5:0];
  assign T_738 = 8'h1 << tgtPages_26;
  assign tgtPagesOH_26 = T_738[5:0];
  assign T_740 = 8'h1 << tgtPages_27;
  assign tgtPagesOH_27 = T_740[5:0];
  assign T_742 = 8'h1 << tgtPages_28;
  assign tgtPagesOH_28 = T_742[5:0];
  assign T_744 = 8'h1 << tgtPages_29;
  assign tgtPagesOH_29 = T_744[5:0];
  assign T_746 = 8'h1 << tgtPages_30;
  assign tgtPagesOH_30 = T_746[5:0];
  assign T_748 = 8'h1 << tgtPages_31;
  assign tgtPagesOH_31 = T_748[5:0];
  assign T_750 = 8'h1 << tgtPages_32;
  assign tgtPagesOH_32 = T_750[5:0];
  assign T_752 = 8'h1 << tgtPages_33;
  assign tgtPagesOH_33 = T_752[5:0];
  assign T_754 = 8'h1 << tgtPages_34;
  assign tgtPagesOH_34 = T_754[5:0];
  assign T_756 = 8'h1 << tgtPages_35;
  assign tgtPagesOH_35 = T_756[5:0];
  assign T_758 = 8'h1 << tgtPages_36;
  assign tgtPagesOH_36 = T_758[5:0];
  assign T_760 = 8'h1 << tgtPages_37;
  assign tgtPagesOH_37 = T_760[5:0];
  assign T_762 = 8'h1 << tgtPages_38;
  assign tgtPagesOH_38 = T_762[5:0];
  assign T_764 = 8'h1 << tgtPages_39;
  assign tgtPagesOH_39 = T_764[5:0];
  assign GEN_7 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : T_778_prediction_valid;
  assign GEN_8 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_taken : T_778_prediction_bits_taken;
  assign GEN_9 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_mask : T_778_prediction_bits_mask;
  assign GEN_10 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bridx : T_778_prediction_bits_bridx;
  assign GEN_11 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_target : T_778_prediction_bits_target;
  assign GEN_12 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : T_778_prediction_bits_entry;
  assign GEN_13 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_history : T_778_prediction_bits_bht_history;
  assign GEN_14 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_value : T_778_prediction_bits_bht_value;
  assign GEN_15 = io_btb_update_valid ? io_btb_update_bits_pc : T_778_pc;
  assign GEN_16 = io_btb_update_valid ? io_btb_update_bits_target : T_778_target;
  assign GEN_17 = io_btb_update_valid ? io_btb_update_bits_taken : T_778_taken;
  assign GEN_18 = io_btb_update_valid ? io_btb_update_bits_isValid : T_778_isValid;
  assign GEN_19 = io_btb_update_valid ? io_btb_update_bits_isJump : T_778_isJump;
  assign GEN_20 = io_btb_update_valid ? io_btb_update_bits_isReturn : T_778_isReturn;
  assign GEN_21 = io_btb_update_valid ? io_btb_update_bits_br_pc : T_778_br_pc;
  assign r_btb_update_valid = T_777;
  assign r_btb_update_bits_prediction_valid = T_778_prediction_valid;
  assign r_btb_update_bits_prediction_bits_taken = T_778_prediction_bits_taken;
  assign r_btb_update_bits_prediction_bits_mask = T_778_prediction_bits_mask;
  assign r_btb_update_bits_prediction_bits_bridx = T_778_prediction_bits_bridx;
  assign r_btb_update_bits_prediction_bits_target = T_778_prediction_bits_target;
  assign r_btb_update_bits_prediction_bits_entry = T_778_prediction_bits_entry;
  assign r_btb_update_bits_prediction_bits_bht_history = T_778_prediction_bits_bht_history;
  assign r_btb_update_bits_prediction_bits_bht_value = T_778_prediction_bits_bht_value;
  assign r_btb_update_bits_pc = T_778_pc;
  assign r_btb_update_bits_target = T_778_target;
  assign r_btb_update_bits_taken = T_778_taken;
  assign r_btb_update_bits_isValid = T_778_isValid;
  assign r_btb_update_bits_isJump = T_778_isJump;
  assign r_btb_update_bits_isReturn = T_778_isReturn;
  assign r_btb_update_bits_br_pc = T_778_br_pc;
  assign T_964 = io_req_bits_addr[38:12];
  assign T_965 = pages_0 == T_964;
  assign T_966 = pages_1 == T_964;
  assign T_967 = pages_2 == T_964;
  assign T_968 = pages_3 == T_964;
  assign T_969 = pages_4 == T_964;
  assign T_970 = pages_5 == T_964;
  assign T_971 = {T_967,T_966};
  assign T_972 = {T_971,T_965};
  assign T_973 = {T_970,T_969};
  assign T_974 = {T_973,T_968};
  assign T_975 = {T_974,T_972};
  assign pageHit = pageValid & T_975;
  assign T_976 = io_req_bits_addr[11:1];
  assign T_977 = idxs_0 == T_976;
  assign T_979 = idxs_1 == T_976;
  assign T_981 = idxs_2 == T_976;
  assign T_983 = idxs_3 == T_976;
  assign T_985 = idxs_4 == T_976;
  assign T_987 = idxs_5 == T_976;
  assign T_989 = idxs_6 == T_976;
  assign T_991 = idxs_7 == T_976;
  assign T_993 = idxs_8 == T_976;
  assign T_995 = idxs_9 == T_976;
  assign T_997 = idxs_10 == T_976;
  assign T_999 = idxs_11 == T_976;
  assign T_1001 = idxs_12 == T_976;
  assign T_1003 = idxs_13 == T_976;
  assign T_1005 = idxs_14 == T_976;
  assign T_1007 = idxs_15 == T_976;
  assign T_1009 = idxs_16 == T_976;
  assign T_1011 = idxs_17 == T_976;
  assign T_1013 = idxs_18 == T_976;
  assign T_1015 = idxs_19 == T_976;
  assign T_1017 = idxs_20 == T_976;
  assign T_1019 = idxs_21 == T_976;
  assign T_1021 = idxs_22 == T_976;
  assign T_1023 = idxs_23 == T_976;
  assign T_1025 = idxs_24 == T_976;
  assign T_1027 = idxs_25 == T_976;
  assign T_1029 = idxs_26 == T_976;
  assign T_1031 = idxs_27 == T_976;
  assign T_1033 = idxs_28 == T_976;
  assign T_1035 = idxs_29 == T_976;
  assign T_1037 = idxs_30 == T_976;
  assign T_1039 = idxs_31 == T_976;
  assign T_1041 = idxs_32 == T_976;
  assign T_1043 = idxs_33 == T_976;
  assign T_1045 = idxs_34 == T_976;
  assign T_1047 = idxs_35 == T_976;
  assign T_1049 = idxs_36 == T_976;
  assign T_1051 = idxs_37 == T_976;
  assign T_1053 = idxs_38 == T_976;
  assign T_1055 = idxs_39 == T_976;
  assign T_1056 = {T_979,T_977};
  assign T_1057 = {T_985,T_983};
  assign T_1058 = {T_1057,T_981};
  assign T_1059 = {T_1058,T_1056};
  assign T_1060 = {T_989,T_987};
  assign T_1061 = {T_995,T_993};
  assign T_1062 = {T_1061,T_991};
  assign T_1063 = {T_1062,T_1060};
  assign T_1064 = {T_1063,T_1059};
  assign T_1065 = {T_999,T_997};
  assign T_1066 = {T_1005,T_1003};
  assign T_1067 = {T_1066,T_1001};
  assign T_1068 = {T_1067,T_1065};
  assign T_1069 = {T_1009,T_1007};
  assign T_1070 = {T_1015,T_1013};
  assign T_1071 = {T_1070,T_1011};
  assign T_1072 = {T_1071,T_1069};
  assign T_1073 = {T_1072,T_1068};
  assign T_1074 = {T_1073,T_1064};
  assign T_1075 = {T_1019,T_1017};
  assign T_1076 = {T_1025,T_1023};
  assign T_1077 = {T_1076,T_1021};
  assign T_1078 = {T_1077,T_1075};
  assign T_1079 = {T_1029,T_1027};
  assign T_1080 = {T_1035,T_1033};
  assign T_1081 = {T_1080,T_1031};
  assign T_1082 = {T_1081,T_1079};
  assign T_1083 = {T_1082,T_1078};
  assign T_1084 = {T_1039,T_1037};
  assign T_1085 = {T_1045,T_1043};
  assign T_1086 = {T_1085,T_1041};
  assign T_1087 = {T_1086,T_1084};
  assign T_1088 = {T_1049,T_1047};
  assign T_1089 = {T_1055,T_1053};
  assign T_1090 = {T_1089,T_1051};
  assign T_1091 = {T_1090,T_1088};
  assign T_1092 = {T_1091,T_1087};
  assign T_1093 = {T_1092,T_1083};
  assign T_1094 = {T_1093,T_1074};
  assign T_1095 = idxPagesOH_0 & pageHit;
  assign T_1096 = idxPagesOH_1 & pageHit;
  assign T_1097 = idxPagesOH_2 & pageHit;
  assign T_1098 = idxPagesOH_3 & pageHit;
  assign T_1099 = idxPagesOH_4 & pageHit;
  assign T_1100 = idxPagesOH_5 & pageHit;
  assign T_1101 = idxPagesOH_6 & pageHit;
  assign T_1102 = idxPagesOH_7 & pageHit;
  assign T_1103 = idxPagesOH_8 & pageHit;
  assign T_1104 = idxPagesOH_9 & pageHit;
  assign T_1105 = idxPagesOH_10 & pageHit;
  assign T_1106 = idxPagesOH_11 & pageHit;
  assign T_1107 = idxPagesOH_12 & pageHit;
  assign T_1108 = idxPagesOH_13 & pageHit;
  assign T_1109 = idxPagesOH_14 & pageHit;
  assign T_1110 = idxPagesOH_15 & pageHit;
  assign T_1111 = idxPagesOH_16 & pageHit;
  assign T_1112 = idxPagesOH_17 & pageHit;
  assign T_1113 = idxPagesOH_18 & pageHit;
  assign T_1114 = idxPagesOH_19 & pageHit;
  assign T_1115 = idxPagesOH_20 & pageHit;
  assign T_1116 = idxPagesOH_21 & pageHit;
  assign T_1117 = idxPagesOH_22 & pageHit;
  assign T_1118 = idxPagesOH_23 & pageHit;
  assign T_1119 = idxPagesOH_24 & pageHit;
  assign T_1120 = idxPagesOH_25 & pageHit;
  assign T_1121 = idxPagesOH_26 & pageHit;
  assign T_1122 = idxPagesOH_27 & pageHit;
  assign T_1123 = idxPagesOH_28 & pageHit;
  assign T_1124 = idxPagesOH_29 & pageHit;
  assign T_1125 = idxPagesOH_30 & pageHit;
  assign T_1126 = idxPagesOH_31 & pageHit;
  assign T_1127 = idxPagesOH_32 & pageHit;
  assign T_1128 = idxPagesOH_33 & pageHit;
  assign T_1129 = idxPagesOH_34 & pageHit;
  assign T_1130 = idxPagesOH_35 & pageHit;
  assign T_1131 = idxPagesOH_36 & pageHit;
  assign T_1132 = idxPagesOH_37 & pageHit;
  assign T_1133 = idxPagesOH_38 & pageHit;
  assign T_1134 = idxPagesOH_39 & pageHit;
  assign T_1136 = T_1095 != 6'h0;
  assign T_1138 = T_1096 != 6'h0;
  assign T_1140 = T_1097 != 6'h0;
  assign T_1142 = T_1098 != 6'h0;
  assign T_1144 = T_1099 != 6'h0;
  assign T_1146 = T_1100 != 6'h0;
  assign T_1148 = T_1101 != 6'h0;
  assign T_1150 = T_1102 != 6'h0;
  assign T_1152 = T_1103 != 6'h0;
  assign T_1154 = T_1104 != 6'h0;
  assign T_1156 = T_1105 != 6'h0;
  assign T_1158 = T_1106 != 6'h0;
  assign T_1160 = T_1107 != 6'h0;
  assign T_1162 = T_1108 != 6'h0;
  assign T_1164 = T_1109 != 6'h0;
  assign T_1166 = T_1110 != 6'h0;
  assign T_1168 = T_1111 != 6'h0;
  assign T_1170 = T_1112 != 6'h0;
  assign T_1172 = T_1113 != 6'h0;
  assign T_1174 = T_1114 != 6'h0;
  assign T_1176 = T_1115 != 6'h0;
  assign T_1178 = T_1116 != 6'h0;
  assign T_1180 = T_1117 != 6'h0;
  assign T_1182 = T_1118 != 6'h0;
  assign T_1184 = T_1119 != 6'h0;
  assign T_1186 = T_1120 != 6'h0;
  assign T_1188 = T_1121 != 6'h0;
  assign T_1190 = T_1122 != 6'h0;
  assign T_1192 = T_1123 != 6'h0;
  assign T_1194 = T_1124 != 6'h0;
  assign T_1196 = T_1125 != 6'h0;
  assign T_1198 = T_1126 != 6'h0;
  assign T_1200 = T_1127 != 6'h0;
  assign T_1202 = T_1128 != 6'h0;
  assign T_1204 = T_1129 != 6'h0;
  assign T_1206 = T_1130 != 6'h0;
  assign T_1208 = T_1131 != 6'h0;
  assign T_1210 = T_1132 != 6'h0;
  assign T_1212 = T_1133 != 6'h0;
  assign T_1214 = T_1134 != 6'h0;
  assign T_1215 = {T_1138,T_1136};
  assign T_1216 = {T_1144,T_1142};
  assign T_1217 = {T_1216,T_1140};
  assign T_1218 = {T_1217,T_1215};
  assign T_1219 = {T_1148,T_1146};
  assign T_1220 = {T_1154,T_1152};
  assign T_1221 = {T_1220,T_1150};
  assign T_1222 = {T_1221,T_1219};
  assign T_1223 = {T_1222,T_1218};
  assign T_1224 = {T_1158,T_1156};
  assign T_1225 = {T_1164,T_1162};
  assign T_1226 = {T_1225,T_1160};
  assign T_1227 = {T_1226,T_1224};
  assign T_1228 = {T_1168,T_1166};
  assign T_1229 = {T_1174,T_1172};
  assign T_1230 = {T_1229,T_1170};
  assign T_1231 = {T_1230,T_1228};
  assign T_1232 = {T_1231,T_1227};
  assign T_1233 = {T_1232,T_1223};
  assign T_1234 = {T_1178,T_1176};
  assign T_1235 = {T_1184,T_1182};
  assign T_1236 = {T_1235,T_1180};
  assign T_1237 = {T_1236,T_1234};
  assign T_1238 = {T_1188,T_1186};
  assign T_1239 = {T_1194,T_1192};
  assign T_1240 = {T_1239,T_1190};
  assign T_1241 = {T_1240,T_1238};
  assign T_1242 = {T_1241,T_1237};
  assign T_1243 = {T_1198,T_1196};
  assign T_1244 = {T_1204,T_1202};
  assign T_1245 = {T_1244,T_1200};
  assign T_1246 = {T_1245,T_1243};
  assign T_1247 = {T_1208,T_1206};
  assign T_1248 = {T_1214,T_1212};
  assign T_1249 = {T_1248,T_1210};
  assign T_1250 = {T_1249,T_1247};
  assign T_1251 = {T_1250,T_1246};
  assign T_1252 = {T_1251,T_1242};
  assign T_1253 = {T_1252,T_1233};
  assign T_1254 = T_1094 & T_1253;
  assign hitsVec = T_1254 & isValid;
  assign T_1255 = r_btb_update_bits_pc[38:12];
  assign T_1256 = pages_0 == T_1255;
  assign T_1257 = pages_1 == T_1255;
  assign T_1258 = pages_2 == T_1255;
  assign T_1259 = pages_3 == T_1255;
  assign T_1260 = pages_4 == T_1255;
  assign T_1261 = pages_5 == T_1255;
  assign T_1262 = {T_1258,T_1257};
  assign T_1263 = {T_1262,T_1256};
  assign T_1264 = {T_1261,T_1260};
  assign T_1265 = {T_1264,T_1259};
  assign T_1266 = {T_1265,T_1263};
  assign updatePageHit = pageValid & T_1266;
  assign T_1267 = r_btb_update_bits_pc[11:1];
  assign T_1547 = r_btb_update_bits_prediction_valid == 1'h0;
  assign T_1548 = r_btb_update_valid & T_1547;
  assign T_1551 = nextRepl == 6'h27;
  assign T_1553 = nextRepl + 6'h1;
  assign T_1554 = T_1553[5:0];
  assign GEN_22 = T_1551 ? 6'h0 : T_1554;
  assign GEN_23 = T_1548 ? GEN_22 : nextRepl;
  assign useUpdatePageHit = updatePageHit != 6'h0;
  assign usePageHit = pageHit != 6'h0;
  assign doIdxPageRepl = useUpdatePageHit == 1'h0;
  assign T_1561 = pageHit[4:0];
  assign T_1562 = pageHit[5];
  assign T_1563 = {T_1561,T_1562};
  assign T_1565 = 8'h1 << nextPageRepl;
  assign idxPageRepl = usePageHit ? {{2'd0}, T_1563} : T_1565;
  assign idxPageUpdateOH = useUpdatePageHit ? {{2'd0}, updatePageHit} : idxPageRepl;
  assign T_1566 = idxPageUpdateOH[7:4];
  assign T_1567 = idxPageUpdateOH[3:0];
  assign T_1569 = T_1566 != 4'h0;
  assign T_1570 = T_1566 | T_1567;
  assign T_1571 = T_1570[3:2];
  assign T_1572 = T_1570[1:0];
  assign T_1574 = T_1571 != 2'h0;
  assign T_1575 = T_1571 | T_1572;
  assign T_1576 = T_1575[1];
  assign T_1577 = {T_1574,T_1576};
  assign idxPageUpdate = {T_1569,T_1577};
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 8'h0;
  assign samePage = T_1255 == T_964;
  assign T_1582 = samePage == 1'h0;
  assign T_1584 = usePageHit == 1'h0;
  assign doTgtPageRepl = T_1582 & T_1584;
  assign T_1585 = idxPageUpdateOH[4:0];
  assign T_1586 = idxPageUpdateOH[5];
  assign T_1587 = {T_1585,T_1586};
  assign tgtPageRepl = samePage ? idxPageUpdateOH : {{2'd0}, T_1587};
  assign T_1588 = usePageHit ? {{2'd0}, pageHit} : tgtPageRepl;
  assign T_1589 = T_1588[7:4];
  assign T_1590 = T_1588[3:0];
  assign T_1592 = T_1589 != 4'h0;
  assign T_1593 = T_1589 | T_1590;
  assign T_1594 = T_1593[3:2];
  assign T_1595 = T_1593[1:0];
  assign T_1597 = T_1594 != 2'h0;
  assign T_1598 = T_1594 | T_1595;
  assign T_1599 = T_1598[1];
  assign T_1600 = {T_1597,T_1599};
  assign tgtPageUpdate = {T_1592,T_1600};
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 8'h0;
  assign T_1602 = doIdxPageRepl | doTgtPageRepl;
  assign T_1603 = r_btb_update_valid & T_1602;
  assign T_1604 = doIdxPageRepl & doTgtPageRepl;
  assign T_1607 = T_1604 ? 2'h2 : 2'h1;
  assign GEN_478 = {{1'd0}, T_1607};
  assign T_1608 = nextPageRepl + GEN_478;
  assign T_1609 = T_1608[2:0];
  assign T_1611 = T_1609 >= 3'h6;
  assign T_1612 = T_1609[0];
  assign T_1614 = T_1611 ? {{2'd0}, T_1612} : T_1609;
  assign GEN_24 = T_1603 ? T_1614 : nextPageRepl;
  assign T_1615 = r_btb_update_bits_prediction_valid ? r_btb_update_bits_prediction_bits_entry : nextRepl;
  assign T_1617 = 64'h1 << T_1615;
  assign GEN_0 = T_1267;
  assign GEN_25 = 6'h0 == T_1615 ? GEN_0 : idxs_0;
  assign GEN_26 = 6'h1 == T_1615 ? GEN_0 : idxs_1;
  assign GEN_27 = 6'h2 == T_1615 ? GEN_0 : idxs_2;
  assign GEN_28 = 6'h3 == T_1615 ? GEN_0 : idxs_3;
  assign GEN_29 = 6'h4 == T_1615 ? GEN_0 : idxs_4;
  assign GEN_30 = 6'h5 == T_1615 ? GEN_0 : idxs_5;
  assign GEN_31 = 6'h6 == T_1615 ? GEN_0 : idxs_6;
  assign GEN_32 = 6'h7 == T_1615 ? GEN_0 : idxs_7;
  assign GEN_33 = 6'h8 == T_1615 ? GEN_0 : idxs_8;
  assign GEN_34 = 6'h9 == T_1615 ? GEN_0 : idxs_9;
  assign GEN_35 = 6'ha == T_1615 ? GEN_0 : idxs_10;
  assign GEN_36 = 6'hb == T_1615 ? GEN_0 : idxs_11;
  assign GEN_37 = 6'hc == T_1615 ? GEN_0 : idxs_12;
  assign GEN_38 = 6'hd == T_1615 ? GEN_0 : idxs_13;
  assign GEN_39 = 6'he == T_1615 ? GEN_0 : idxs_14;
  assign GEN_40 = 6'hf == T_1615 ? GEN_0 : idxs_15;
  assign GEN_41 = 6'h10 == T_1615 ? GEN_0 : idxs_16;
  assign GEN_42 = 6'h11 == T_1615 ? GEN_0 : idxs_17;
  assign GEN_43 = 6'h12 == T_1615 ? GEN_0 : idxs_18;
  assign GEN_44 = 6'h13 == T_1615 ? GEN_0 : idxs_19;
  assign GEN_45 = 6'h14 == T_1615 ? GEN_0 : idxs_20;
  assign GEN_46 = 6'h15 == T_1615 ? GEN_0 : idxs_21;
  assign GEN_47 = 6'h16 == T_1615 ? GEN_0 : idxs_22;
  assign GEN_48 = 6'h17 == T_1615 ? GEN_0 : idxs_23;
  assign GEN_49 = 6'h18 == T_1615 ? GEN_0 : idxs_24;
  assign GEN_50 = 6'h19 == T_1615 ? GEN_0 : idxs_25;
  assign GEN_51 = 6'h1a == T_1615 ? GEN_0 : idxs_26;
  assign GEN_52 = 6'h1b == T_1615 ? GEN_0 : idxs_27;
  assign GEN_53 = 6'h1c == T_1615 ? GEN_0 : idxs_28;
  assign GEN_54 = 6'h1d == T_1615 ? GEN_0 : idxs_29;
  assign GEN_55 = 6'h1e == T_1615 ? GEN_0 : idxs_30;
  assign GEN_56 = 6'h1f == T_1615 ? GEN_0 : idxs_31;
  assign GEN_57 = 6'h20 == T_1615 ? GEN_0 : idxs_32;
  assign GEN_58 = 6'h21 == T_1615 ? GEN_0 : idxs_33;
  assign GEN_59 = 6'h22 == T_1615 ? GEN_0 : idxs_34;
  assign GEN_60 = 6'h23 == T_1615 ? GEN_0 : idxs_35;
  assign GEN_61 = 6'h24 == T_1615 ? GEN_0 : idxs_36;
  assign GEN_62 = 6'h25 == T_1615 ? GEN_0 : idxs_37;
  assign GEN_63 = 6'h26 == T_1615 ? GEN_0 : idxs_38;
  assign GEN_64 = 6'h27 == T_1615 ? GEN_0 : idxs_39;
  assign GEN_1 = T_976;
  assign GEN_65 = 6'h0 == T_1615 ? GEN_1 : tgts_0;
  assign GEN_66 = 6'h1 == T_1615 ? GEN_1 : tgts_1;
  assign GEN_67 = 6'h2 == T_1615 ? GEN_1 : tgts_2;
  assign GEN_68 = 6'h3 == T_1615 ? GEN_1 : tgts_3;
  assign GEN_69 = 6'h4 == T_1615 ? GEN_1 : tgts_4;
  assign GEN_70 = 6'h5 == T_1615 ? GEN_1 : tgts_5;
  assign GEN_71 = 6'h6 == T_1615 ? GEN_1 : tgts_6;
  assign GEN_72 = 6'h7 == T_1615 ? GEN_1 : tgts_7;
  assign GEN_73 = 6'h8 == T_1615 ? GEN_1 : tgts_8;
  assign GEN_74 = 6'h9 == T_1615 ? GEN_1 : tgts_9;
  assign GEN_75 = 6'ha == T_1615 ? GEN_1 : tgts_10;
  assign GEN_76 = 6'hb == T_1615 ? GEN_1 : tgts_11;
  assign GEN_77 = 6'hc == T_1615 ? GEN_1 : tgts_12;
  assign GEN_78 = 6'hd == T_1615 ? GEN_1 : tgts_13;
  assign GEN_79 = 6'he == T_1615 ? GEN_1 : tgts_14;
  assign GEN_80 = 6'hf == T_1615 ? GEN_1 : tgts_15;
  assign GEN_81 = 6'h10 == T_1615 ? GEN_1 : tgts_16;
  assign GEN_82 = 6'h11 == T_1615 ? GEN_1 : tgts_17;
  assign GEN_83 = 6'h12 == T_1615 ? GEN_1 : tgts_18;
  assign GEN_84 = 6'h13 == T_1615 ? GEN_1 : tgts_19;
  assign GEN_85 = 6'h14 == T_1615 ? GEN_1 : tgts_20;
  assign GEN_86 = 6'h15 == T_1615 ? GEN_1 : tgts_21;
  assign GEN_87 = 6'h16 == T_1615 ? GEN_1 : tgts_22;
  assign GEN_88 = 6'h17 == T_1615 ? GEN_1 : tgts_23;
  assign GEN_89 = 6'h18 == T_1615 ? GEN_1 : tgts_24;
  assign GEN_90 = 6'h19 == T_1615 ? GEN_1 : tgts_25;
  assign GEN_91 = 6'h1a == T_1615 ? GEN_1 : tgts_26;
  assign GEN_92 = 6'h1b == T_1615 ? GEN_1 : tgts_27;
  assign GEN_93 = 6'h1c == T_1615 ? GEN_1 : tgts_28;
  assign GEN_94 = 6'h1d == T_1615 ? GEN_1 : tgts_29;
  assign GEN_95 = 6'h1e == T_1615 ? GEN_1 : tgts_30;
  assign GEN_96 = 6'h1f == T_1615 ? GEN_1 : tgts_31;
  assign GEN_97 = 6'h20 == T_1615 ? GEN_1 : tgts_32;
  assign GEN_98 = 6'h21 == T_1615 ? GEN_1 : tgts_33;
  assign GEN_99 = 6'h22 == T_1615 ? GEN_1 : tgts_34;
  assign GEN_100 = 6'h23 == T_1615 ? GEN_1 : tgts_35;
  assign GEN_101 = 6'h24 == T_1615 ? GEN_1 : tgts_36;
  assign GEN_102 = 6'h25 == T_1615 ? GEN_1 : tgts_37;
  assign GEN_103 = 6'h26 == T_1615 ? GEN_1 : tgts_38;
  assign GEN_104 = 6'h27 == T_1615 ? GEN_1 : tgts_39;
  assign GEN_2 = idxPageUpdate;
  assign GEN_105 = 6'h0 == T_1615 ? GEN_2 : idxPages_0;
  assign GEN_106 = 6'h1 == T_1615 ? GEN_2 : idxPages_1;
  assign GEN_107 = 6'h2 == T_1615 ? GEN_2 : idxPages_2;
  assign GEN_108 = 6'h3 == T_1615 ? GEN_2 : idxPages_3;
  assign GEN_109 = 6'h4 == T_1615 ? GEN_2 : idxPages_4;
  assign GEN_110 = 6'h5 == T_1615 ? GEN_2 : idxPages_5;
  assign GEN_111 = 6'h6 == T_1615 ? GEN_2 : idxPages_6;
  assign GEN_112 = 6'h7 == T_1615 ? GEN_2 : idxPages_7;
  assign GEN_113 = 6'h8 == T_1615 ? GEN_2 : idxPages_8;
  assign GEN_114 = 6'h9 == T_1615 ? GEN_2 : idxPages_9;
  assign GEN_115 = 6'ha == T_1615 ? GEN_2 : idxPages_10;
  assign GEN_116 = 6'hb == T_1615 ? GEN_2 : idxPages_11;
  assign GEN_117 = 6'hc == T_1615 ? GEN_2 : idxPages_12;
  assign GEN_118 = 6'hd == T_1615 ? GEN_2 : idxPages_13;
  assign GEN_119 = 6'he == T_1615 ? GEN_2 : idxPages_14;
  assign GEN_120 = 6'hf == T_1615 ? GEN_2 : idxPages_15;
  assign GEN_121 = 6'h10 == T_1615 ? GEN_2 : idxPages_16;
  assign GEN_122 = 6'h11 == T_1615 ? GEN_2 : idxPages_17;
  assign GEN_123 = 6'h12 == T_1615 ? GEN_2 : idxPages_18;
  assign GEN_124 = 6'h13 == T_1615 ? GEN_2 : idxPages_19;
  assign GEN_125 = 6'h14 == T_1615 ? GEN_2 : idxPages_20;
  assign GEN_126 = 6'h15 == T_1615 ? GEN_2 : idxPages_21;
  assign GEN_127 = 6'h16 == T_1615 ? GEN_2 : idxPages_22;
  assign GEN_128 = 6'h17 == T_1615 ? GEN_2 : idxPages_23;
  assign GEN_129 = 6'h18 == T_1615 ? GEN_2 : idxPages_24;
  assign GEN_130 = 6'h19 == T_1615 ? GEN_2 : idxPages_25;
  assign GEN_131 = 6'h1a == T_1615 ? GEN_2 : idxPages_26;
  assign GEN_132 = 6'h1b == T_1615 ? GEN_2 : idxPages_27;
  assign GEN_133 = 6'h1c == T_1615 ? GEN_2 : idxPages_28;
  assign GEN_134 = 6'h1d == T_1615 ? GEN_2 : idxPages_29;
  assign GEN_135 = 6'h1e == T_1615 ? GEN_2 : idxPages_30;
  assign GEN_136 = 6'h1f == T_1615 ? GEN_2 : idxPages_31;
  assign GEN_137 = 6'h20 == T_1615 ? GEN_2 : idxPages_32;
  assign GEN_138 = 6'h21 == T_1615 ? GEN_2 : idxPages_33;
  assign GEN_139 = 6'h22 == T_1615 ? GEN_2 : idxPages_34;
  assign GEN_140 = 6'h23 == T_1615 ? GEN_2 : idxPages_35;
  assign GEN_141 = 6'h24 == T_1615 ? GEN_2 : idxPages_36;
  assign GEN_142 = 6'h25 == T_1615 ? GEN_2 : idxPages_37;
  assign GEN_143 = 6'h26 == T_1615 ? GEN_2 : idxPages_38;
  assign GEN_144 = 6'h27 == T_1615 ? GEN_2 : idxPages_39;
  assign GEN_3 = tgtPageUpdate;
  assign GEN_145 = 6'h0 == T_1615 ? GEN_3 : tgtPages_0;
  assign GEN_146 = 6'h1 == T_1615 ? GEN_3 : tgtPages_1;
  assign GEN_147 = 6'h2 == T_1615 ? GEN_3 : tgtPages_2;
  assign GEN_148 = 6'h3 == T_1615 ? GEN_3 : tgtPages_3;
  assign GEN_149 = 6'h4 == T_1615 ? GEN_3 : tgtPages_4;
  assign GEN_150 = 6'h5 == T_1615 ? GEN_3 : tgtPages_5;
  assign GEN_151 = 6'h6 == T_1615 ? GEN_3 : tgtPages_6;
  assign GEN_152 = 6'h7 == T_1615 ? GEN_3 : tgtPages_7;
  assign GEN_153 = 6'h8 == T_1615 ? GEN_3 : tgtPages_8;
  assign GEN_154 = 6'h9 == T_1615 ? GEN_3 : tgtPages_9;
  assign GEN_155 = 6'ha == T_1615 ? GEN_3 : tgtPages_10;
  assign GEN_156 = 6'hb == T_1615 ? GEN_3 : tgtPages_11;
  assign GEN_157 = 6'hc == T_1615 ? GEN_3 : tgtPages_12;
  assign GEN_158 = 6'hd == T_1615 ? GEN_3 : tgtPages_13;
  assign GEN_159 = 6'he == T_1615 ? GEN_3 : tgtPages_14;
  assign GEN_160 = 6'hf == T_1615 ? GEN_3 : tgtPages_15;
  assign GEN_161 = 6'h10 == T_1615 ? GEN_3 : tgtPages_16;
  assign GEN_162 = 6'h11 == T_1615 ? GEN_3 : tgtPages_17;
  assign GEN_163 = 6'h12 == T_1615 ? GEN_3 : tgtPages_18;
  assign GEN_164 = 6'h13 == T_1615 ? GEN_3 : tgtPages_19;
  assign GEN_165 = 6'h14 == T_1615 ? GEN_3 : tgtPages_20;
  assign GEN_166 = 6'h15 == T_1615 ? GEN_3 : tgtPages_21;
  assign GEN_167 = 6'h16 == T_1615 ? GEN_3 : tgtPages_22;
  assign GEN_168 = 6'h17 == T_1615 ? GEN_3 : tgtPages_23;
  assign GEN_169 = 6'h18 == T_1615 ? GEN_3 : tgtPages_24;
  assign GEN_170 = 6'h19 == T_1615 ? GEN_3 : tgtPages_25;
  assign GEN_171 = 6'h1a == T_1615 ? GEN_3 : tgtPages_26;
  assign GEN_172 = 6'h1b == T_1615 ? GEN_3 : tgtPages_27;
  assign GEN_173 = 6'h1c == T_1615 ? GEN_3 : tgtPages_28;
  assign GEN_174 = 6'h1d == T_1615 ? GEN_3 : tgtPages_29;
  assign GEN_175 = 6'h1e == T_1615 ? GEN_3 : tgtPages_30;
  assign GEN_176 = 6'h1f == T_1615 ? GEN_3 : tgtPages_31;
  assign GEN_177 = 6'h20 == T_1615 ? GEN_3 : tgtPages_32;
  assign GEN_178 = 6'h21 == T_1615 ? GEN_3 : tgtPages_33;
  assign GEN_179 = 6'h22 == T_1615 ? GEN_3 : tgtPages_34;
  assign GEN_180 = 6'h23 == T_1615 ? GEN_3 : tgtPages_35;
  assign GEN_181 = 6'h24 == T_1615 ? GEN_3 : tgtPages_36;
  assign GEN_182 = 6'h25 == T_1615 ? GEN_3 : tgtPages_37;
  assign GEN_183 = 6'h26 == T_1615 ? GEN_3 : tgtPages_38;
  assign GEN_184 = 6'h27 == T_1615 ? GEN_3 : tgtPages_39;
  assign GEN_479 = {{24'd0}, isValid};
  assign T_1620 = GEN_479 | T_1617;
  assign T_1621 = ~ T_1617;
  assign T_1622 = GEN_479 & T_1621;
  assign T_1623 = r_btb_update_bits_isValid ? T_1620 : T_1622;
  assign GEN_481 = {{24'd0}, isReturn};
  assign T_1624 = GEN_481 | T_1617;
  assign T_1626 = GEN_481 & T_1621;
  assign T_1627 = r_btb_update_bits_isReturn ? T_1624 : T_1626;
  assign GEN_483 = {{24'd0}, isJump};
  assign T_1628 = GEN_483 | T_1617;
  assign T_1630 = GEN_483 & T_1621;
  assign T_1631 = r_btb_update_bits_isJump ? T_1628 : T_1630;
  assign T_1632 = r_btb_update_bits_br_pc[38:1];
  assign GEN_4 = T_1632[0];
  assign GEN_185 = 6'h0 == T_1615 ? GEN_4 : brIdx_0;
  assign GEN_186 = 6'h1 == T_1615 ? GEN_4 : brIdx_1;
  assign GEN_187 = 6'h2 == T_1615 ? GEN_4 : brIdx_2;
  assign GEN_188 = 6'h3 == T_1615 ? GEN_4 : brIdx_3;
  assign GEN_189 = 6'h4 == T_1615 ? GEN_4 : brIdx_4;
  assign GEN_190 = 6'h5 == T_1615 ? GEN_4 : brIdx_5;
  assign GEN_191 = 6'h6 == T_1615 ? GEN_4 : brIdx_6;
  assign GEN_192 = 6'h7 == T_1615 ? GEN_4 : brIdx_7;
  assign GEN_193 = 6'h8 == T_1615 ? GEN_4 : brIdx_8;
  assign GEN_194 = 6'h9 == T_1615 ? GEN_4 : brIdx_9;
  assign GEN_195 = 6'ha == T_1615 ? GEN_4 : brIdx_10;
  assign GEN_196 = 6'hb == T_1615 ? GEN_4 : brIdx_11;
  assign GEN_197 = 6'hc == T_1615 ? GEN_4 : brIdx_12;
  assign GEN_198 = 6'hd == T_1615 ? GEN_4 : brIdx_13;
  assign GEN_199 = 6'he == T_1615 ? GEN_4 : brIdx_14;
  assign GEN_200 = 6'hf == T_1615 ? GEN_4 : brIdx_15;
  assign GEN_201 = 6'h10 == T_1615 ? GEN_4 : brIdx_16;
  assign GEN_202 = 6'h11 == T_1615 ? GEN_4 : brIdx_17;
  assign GEN_203 = 6'h12 == T_1615 ? GEN_4 : brIdx_18;
  assign GEN_204 = 6'h13 == T_1615 ? GEN_4 : brIdx_19;
  assign GEN_205 = 6'h14 == T_1615 ? GEN_4 : brIdx_20;
  assign GEN_206 = 6'h15 == T_1615 ? GEN_4 : brIdx_21;
  assign GEN_207 = 6'h16 == T_1615 ? GEN_4 : brIdx_22;
  assign GEN_208 = 6'h17 == T_1615 ? GEN_4 : brIdx_23;
  assign GEN_209 = 6'h18 == T_1615 ? GEN_4 : brIdx_24;
  assign GEN_210 = 6'h19 == T_1615 ? GEN_4 : brIdx_25;
  assign GEN_211 = 6'h1a == T_1615 ? GEN_4 : brIdx_26;
  assign GEN_212 = 6'h1b == T_1615 ? GEN_4 : brIdx_27;
  assign GEN_213 = 6'h1c == T_1615 ? GEN_4 : brIdx_28;
  assign GEN_214 = 6'h1d == T_1615 ? GEN_4 : brIdx_29;
  assign GEN_215 = 6'h1e == T_1615 ? GEN_4 : brIdx_30;
  assign GEN_216 = 6'h1f == T_1615 ? GEN_4 : brIdx_31;
  assign GEN_217 = 6'h20 == T_1615 ? GEN_4 : brIdx_32;
  assign GEN_218 = 6'h21 == T_1615 ? GEN_4 : brIdx_33;
  assign GEN_219 = 6'h22 == T_1615 ? GEN_4 : brIdx_34;
  assign GEN_220 = 6'h23 == T_1615 ? GEN_4 : brIdx_35;
  assign GEN_221 = 6'h24 == T_1615 ? GEN_4 : brIdx_36;
  assign GEN_222 = 6'h25 == T_1615 ? GEN_4 : brIdx_37;
  assign GEN_223 = 6'h26 == T_1615 ? GEN_4 : brIdx_38;
  assign GEN_224 = 6'h27 == T_1615 ? GEN_4 : brIdx_39;
  assign T_1633 = idxPageUpdate[0];
  assign T_1635 = T_1633 == 1'h0;
  assign T_1636 = T_1635 ? idxPageReplEn : tgtPageReplEn;
  assign T_1639 = T_1635 ? T_1255 : T_964;
  assign T_1640 = T_1636[0];
  assign GEN_225 = T_1640 ? T_1639 : pages_0;
  assign T_1641 = T_1636[2];
  assign GEN_226 = T_1641 ? T_1639 : pages_2;
  assign T_1642 = T_1636[4];
  assign GEN_227 = T_1642 ? T_1639 : pages_4;
  assign T_1643 = T_1635 ? tgtPageReplEn : idxPageReplEn;
  assign T_1646 = T_1635 ? T_964 : T_1255;
  assign T_1647 = T_1643[1];
  assign GEN_228 = T_1647 ? T_1646 : pages_1;
  assign T_1648 = T_1643[3];
  assign GEN_229 = T_1648 ? T_1646 : pages_3;
  assign T_1649 = T_1643[5];
  assign GEN_230 = T_1649 ? T_1646 : pages_5;
  assign GEN_485 = {{2'd0}, pageValid};
  assign T_1650 = GEN_485 | tgtPageReplEn;
  assign T_1651 = T_1650 | idxPageReplEn;
  assign GEN_232 = r_btb_update_valid ? GEN_25 : idxs_0;
  assign GEN_233 = r_btb_update_valid ? GEN_26 : idxs_1;
  assign GEN_234 = r_btb_update_valid ? GEN_27 : idxs_2;
  assign GEN_235 = r_btb_update_valid ? GEN_28 : idxs_3;
  assign GEN_236 = r_btb_update_valid ? GEN_29 : idxs_4;
  assign GEN_237 = r_btb_update_valid ? GEN_30 : idxs_5;
  assign GEN_238 = r_btb_update_valid ? GEN_31 : idxs_6;
  assign GEN_239 = r_btb_update_valid ? GEN_32 : idxs_7;
  assign GEN_240 = r_btb_update_valid ? GEN_33 : idxs_8;
  assign GEN_241 = r_btb_update_valid ? GEN_34 : idxs_9;
  assign GEN_242 = r_btb_update_valid ? GEN_35 : idxs_10;
  assign GEN_243 = r_btb_update_valid ? GEN_36 : idxs_11;
  assign GEN_244 = r_btb_update_valid ? GEN_37 : idxs_12;
  assign GEN_245 = r_btb_update_valid ? GEN_38 : idxs_13;
  assign GEN_246 = r_btb_update_valid ? GEN_39 : idxs_14;
  assign GEN_247 = r_btb_update_valid ? GEN_40 : idxs_15;
  assign GEN_248 = r_btb_update_valid ? GEN_41 : idxs_16;
  assign GEN_249 = r_btb_update_valid ? GEN_42 : idxs_17;
  assign GEN_250 = r_btb_update_valid ? GEN_43 : idxs_18;
  assign GEN_251 = r_btb_update_valid ? GEN_44 : idxs_19;
  assign GEN_252 = r_btb_update_valid ? GEN_45 : idxs_20;
  assign GEN_253 = r_btb_update_valid ? GEN_46 : idxs_21;
  assign GEN_254 = r_btb_update_valid ? GEN_47 : idxs_22;
  assign GEN_255 = r_btb_update_valid ? GEN_48 : idxs_23;
  assign GEN_256 = r_btb_update_valid ? GEN_49 : idxs_24;
  assign GEN_257 = r_btb_update_valid ? GEN_50 : idxs_25;
  assign GEN_258 = r_btb_update_valid ? GEN_51 : idxs_26;
  assign GEN_259 = r_btb_update_valid ? GEN_52 : idxs_27;
  assign GEN_260 = r_btb_update_valid ? GEN_53 : idxs_28;
  assign GEN_261 = r_btb_update_valid ? GEN_54 : idxs_29;
  assign GEN_262 = r_btb_update_valid ? GEN_55 : idxs_30;
  assign GEN_263 = r_btb_update_valid ? GEN_56 : idxs_31;
  assign GEN_264 = r_btb_update_valid ? GEN_57 : idxs_32;
  assign GEN_265 = r_btb_update_valid ? GEN_58 : idxs_33;
  assign GEN_266 = r_btb_update_valid ? GEN_59 : idxs_34;
  assign GEN_267 = r_btb_update_valid ? GEN_60 : idxs_35;
  assign GEN_268 = r_btb_update_valid ? GEN_61 : idxs_36;
  assign GEN_269 = r_btb_update_valid ? GEN_62 : idxs_37;
  assign GEN_270 = r_btb_update_valid ? GEN_63 : idxs_38;
  assign GEN_271 = r_btb_update_valid ? GEN_64 : idxs_39;
  assign GEN_273 = r_btb_update_valid ? GEN_65 : tgts_0;
  assign GEN_274 = r_btb_update_valid ? GEN_66 : tgts_1;
  assign GEN_275 = r_btb_update_valid ? GEN_67 : tgts_2;
  assign GEN_276 = r_btb_update_valid ? GEN_68 : tgts_3;
  assign GEN_277 = r_btb_update_valid ? GEN_69 : tgts_4;
  assign GEN_278 = r_btb_update_valid ? GEN_70 : tgts_5;
  assign GEN_279 = r_btb_update_valid ? GEN_71 : tgts_6;
  assign GEN_280 = r_btb_update_valid ? GEN_72 : tgts_7;
  assign GEN_281 = r_btb_update_valid ? GEN_73 : tgts_8;
  assign GEN_282 = r_btb_update_valid ? GEN_74 : tgts_9;
  assign GEN_283 = r_btb_update_valid ? GEN_75 : tgts_10;
  assign GEN_284 = r_btb_update_valid ? GEN_76 : tgts_11;
  assign GEN_285 = r_btb_update_valid ? GEN_77 : tgts_12;
  assign GEN_286 = r_btb_update_valid ? GEN_78 : tgts_13;
  assign GEN_287 = r_btb_update_valid ? GEN_79 : tgts_14;
  assign GEN_288 = r_btb_update_valid ? GEN_80 : tgts_15;
  assign GEN_289 = r_btb_update_valid ? GEN_81 : tgts_16;
  assign GEN_290 = r_btb_update_valid ? GEN_82 : tgts_17;
  assign GEN_291 = r_btb_update_valid ? GEN_83 : tgts_18;
  assign GEN_292 = r_btb_update_valid ? GEN_84 : tgts_19;
  assign GEN_293 = r_btb_update_valid ? GEN_85 : tgts_20;
  assign GEN_294 = r_btb_update_valid ? GEN_86 : tgts_21;
  assign GEN_295 = r_btb_update_valid ? GEN_87 : tgts_22;
  assign GEN_296 = r_btb_update_valid ? GEN_88 : tgts_23;
  assign GEN_297 = r_btb_update_valid ? GEN_89 : tgts_24;
  assign GEN_298 = r_btb_update_valid ? GEN_90 : tgts_25;
  assign GEN_299 = r_btb_update_valid ? GEN_91 : tgts_26;
  assign GEN_300 = r_btb_update_valid ? GEN_92 : tgts_27;
  assign GEN_301 = r_btb_update_valid ? GEN_93 : tgts_28;
  assign GEN_302 = r_btb_update_valid ? GEN_94 : tgts_29;
  assign GEN_303 = r_btb_update_valid ? GEN_95 : tgts_30;
  assign GEN_304 = r_btb_update_valid ? GEN_96 : tgts_31;
  assign GEN_305 = r_btb_update_valid ? GEN_97 : tgts_32;
  assign GEN_306 = r_btb_update_valid ? GEN_98 : tgts_33;
  assign GEN_307 = r_btb_update_valid ? GEN_99 : tgts_34;
  assign GEN_308 = r_btb_update_valid ? GEN_100 : tgts_35;
  assign GEN_309 = r_btb_update_valid ? GEN_101 : tgts_36;
  assign GEN_310 = r_btb_update_valid ? GEN_102 : tgts_37;
  assign GEN_311 = r_btb_update_valid ? GEN_103 : tgts_38;
  assign GEN_312 = r_btb_update_valid ? GEN_104 : tgts_39;
  assign GEN_314 = r_btb_update_valid ? GEN_105 : idxPages_0;
  assign GEN_315 = r_btb_update_valid ? GEN_106 : idxPages_1;
  assign GEN_316 = r_btb_update_valid ? GEN_107 : idxPages_2;
  assign GEN_317 = r_btb_update_valid ? GEN_108 : idxPages_3;
  assign GEN_318 = r_btb_update_valid ? GEN_109 : idxPages_4;
  assign GEN_319 = r_btb_update_valid ? GEN_110 : idxPages_5;
  assign GEN_320 = r_btb_update_valid ? GEN_111 : idxPages_6;
  assign GEN_321 = r_btb_update_valid ? GEN_112 : idxPages_7;
  assign GEN_322 = r_btb_update_valid ? GEN_113 : idxPages_8;
  assign GEN_323 = r_btb_update_valid ? GEN_114 : idxPages_9;
  assign GEN_324 = r_btb_update_valid ? GEN_115 : idxPages_10;
  assign GEN_325 = r_btb_update_valid ? GEN_116 : idxPages_11;
  assign GEN_326 = r_btb_update_valid ? GEN_117 : idxPages_12;
  assign GEN_327 = r_btb_update_valid ? GEN_118 : idxPages_13;
  assign GEN_328 = r_btb_update_valid ? GEN_119 : idxPages_14;
  assign GEN_329 = r_btb_update_valid ? GEN_120 : idxPages_15;
  assign GEN_330 = r_btb_update_valid ? GEN_121 : idxPages_16;
  assign GEN_331 = r_btb_update_valid ? GEN_122 : idxPages_17;
  assign GEN_332 = r_btb_update_valid ? GEN_123 : idxPages_18;
  assign GEN_333 = r_btb_update_valid ? GEN_124 : idxPages_19;
  assign GEN_334 = r_btb_update_valid ? GEN_125 : idxPages_20;
  assign GEN_335 = r_btb_update_valid ? GEN_126 : idxPages_21;
  assign GEN_336 = r_btb_update_valid ? GEN_127 : idxPages_22;
  assign GEN_337 = r_btb_update_valid ? GEN_128 : idxPages_23;
  assign GEN_338 = r_btb_update_valid ? GEN_129 : idxPages_24;
  assign GEN_339 = r_btb_update_valid ? GEN_130 : idxPages_25;
  assign GEN_340 = r_btb_update_valid ? GEN_131 : idxPages_26;
  assign GEN_341 = r_btb_update_valid ? GEN_132 : idxPages_27;
  assign GEN_342 = r_btb_update_valid ? GEN_133 : idxPages_28;
  assign GEN_343 = r_btb_update_valid ? GEN_134 : idxPages_29;
  assign GEN_344 = r_btb_update_valid ? GEN_135 : idxPages_30;
  assign GEN_345 = r_btb_update_valid ? GEN_136 : idxPages_31;
  assign GEN_346 = r_btb_update_valid ? GEN_137 : idxPages_32;
  assign GEN_347 = r_btb_update_valid ? GEN_138 : idxPages_33;
  assign GEN_348 = r_btb_update_valid ? GEN_139 : idxPages_34;
  assign GEN_349 = r_btb_update_valid ? GEN_140 : idxPages_35;
  assign GEN_350 = r_btb_update_valid ? GEN_141 : idxPages_36;
  assign GEN_351 = r_btb_update_valid ? GEN_142 : idxPages_37;
  assign GEN_352 = r_btb_update_valid ? GEN_143 : idxPages_38;
  assign GEN_353 = r_btb_update_valid ? GEN_144 : idxPages_39;
  assign GEN_355 = r_btb_update_valid ? GEN_145 : tgtPages_0;
  assign GEN_356 = r_btb_update_valid ? GEN_146 : tgtPages_1;
  assign GEN_357 = r_btb_update_valid ? GEN_147 : tgtPages_2;
  assign GEN_358 = r_btb_update_valid ? GEN_148 : tgtPages_3;
  assign GEN_359 = r_btb_update_valid ? GEN_149 : tgtPages_4;
  assign GEN_360 = r_btb_update_valid ? GEN_150 : tgtPages_5;
  assign GEN_361 = r_btb_update_valid ? GEN_151 : tgtPages_6;
  assign GEN_362 = r_btb_update_valid ? GEN_152 : tgtPages_7;
  assign GEN_363 = r_btb_update_valid ? GEN_153 : tgtPages_8;
  assign GEN_364 = r_btb_update_valid ? GEN_154 : tgtPages_9;
  assign GEN_365 = r_btb_update_valid ? GEN_155 : tgtPages_10;
  assign GEN_366 = r_btb_update_valid ? GEN_156 : tgtPages_11;
  assign GEN_367 = r_btb_update_valid ? GEN_157 : tgtPages_12;
  assign GEN_368 = r_btb_update_valid ? GEN_158 : tgtPages_13;
  assign GEN_369 = r_btb_update_valid ? GEN_159 : tgtPages_14;
  assign GEN_370 = r_btb_update_valid ? GEN_160 : tgtPages_15;
  assign GEN_371 = r_btb_update_valid ? GEN_161 : tgtPages_16;
  assign GEN_372 = r_btb_update_valid ? GEN_162 : tgtPages_17;
  assign GEN_373 = r_btb_update_valid ? GEN_163 : tgtPages_18;
  assign GEN_374 = r_btb_update_valid ? GEN_164 : tgtPages_19;
  assign GEN_375 = r_btb_update_valid ? GEN_165 : tgtPages_20;
  assign GEN_376 = r_btb_update_valid ? GEN_166 : tgtPages_21;
  assign GEN_377 = r_btb_update_valid ? GEN_167 : tgtPages_22;
  assign GEN_378 = r_btb_update_valid ? GEN_168 : tgtPages_23;
  assign GEN_379 = r_btb_update_valid ? GEN_169 : tgtPages_24;
  assign GEN_380 = r_btb_update_valid ? GEN_170 : tgtPages_25;
  assign GEN_381 = r_btb_update_valid ? GEN_171 : tgtPages_26;
  assign GEN_382 = r_btb_update_valid ? GEN_172 : tgtPages_27;
  assign GEN_383 = r_btb_update_valid ? GEN_173 : tgtPages_28;
  assign GEN_384 = r_btb_update_valid ? GEN_174 : tgtPages_29;
  assign GEN_385 = r_btb_update_valid ? GEN_175 : tgtPages_30;
  assign GEN_386 = r_btb_update_valid ? GEN_176 : tgtPages_31;
  assign GEN_387 = r_btb_update_valid ? GEN_177 : tgtPages_32;
  assign GEN_388 = r_btb_update_valid ? GEN_178 : tgtPages_33;
  assign GEN_389 = r_btb_update_valid ? GEN_179 : tgtPages_34;
  assign GEN_390 = r_btb_update_valid ? GEN_180 : tgtPages_35;
  assign GEN_391 = r_btb_update_valid ? GEN_181 : tgtPages_36;
  assign GEN_392 = r_btb_update_valid ? GEN_182 : tgtPages_37;
  assign GEN_393 = r_btb_update_valid ? GEN_183 : tgtPages_38;
  assign GEN_394 = r_btb_update_valid ? GEN_184 : tgtPages_39;
  assign GEN_395 = r_btb_update_valid ? T_1623 : {{24'd0}, isValid};
  assign GEN_396 = r_btb_update_valid ? T_1627 : {{24'd0}, isReturn};
  assign GEN_397 = r_btb_update_valid ? T_1631 : {{24'd0}, isJump};
  assign GEN_399 = r_btb_update_valid ? GEN_185 : brIdx_0;
  assign GEN_400 = r_btb_update_valid ? GEN_186 : brIdx_1;
  assign GEN_401 = r_btb_update_valid ? GEN_187 : brIdx_2;
  assign GEN_402 = r_btb_update_valid ? GEN_188 : brIdx_3;
  assign GEN_403 = r_btb_update_valid ? GEN_189 : brIdx_4;
  assign GEN_404 = r_btb_update_valid ? GEN_190 : brIdx_5;
  assign GEN_405 = r_btb_update_valid ? GEN_191 : brIdx_6;
  assign GEN_406 = r_btb_update_valid ? GEN_192 : brIdx_7;
  assign GEN_407 = r_btb_update_valid ? GEN_193 : brIdx_8;
  assign GEN_408 = r_btb_update_valid ? GEN_194 : brIdx_9;
  assign GEN_409 = r_btb_update_valid ? GEN_195 : brIdx_10;
  assign GEN_410 = r_btb_update_valid ? GEN_196 : brIdx_11;
  assign GEN_411 = r_btb_update_valid ? GEN_197 : brIdx_12;
  assign GEN_412 = r_btb_update_valid ? GEN_198 : brIdx_13;
  assign GEN_413 = r_btb_update_valid ? GEN_199 : brIdx_14;
  assign GEN_414 = r_btb_update_valid ? GEN_200 : brIdx_15;
  assign GEN_415 = r_btb_update_valid ? GEN_201 : brIdx_16;
  assign GEN_416 = r_btb_update_valid ? GEN_202 : brIdx_17;
  assign GEN_417 = r_btb_update_valid ? GEN_203 : brIdx_18;
  assign GEN_418 = r_btb_update_valid ? GEN_204 : brIdx_19;
  assign GEN_419 = r_btb_update_valid ? GEN_205 : brIdx_20;
  assign GEN_420 = r_btb_update_valid ? GEN_206 : brIdx_21;
  assign GEN_421 = r_btb_update_valid ? GEN_207 : brIdx_22;
  assign GEN_422 = r_btb_update_valid ? GEN_208 : brIdx_23;
  assign GEN_423 = r_btb_update_valid ? GEN_209 : brIdx_24;
  assign GEN_424 = r_btb_update_valid ? GEN_210 : brIdx_25;
  assign GEN_425 = r_btb_update_valid ? GEN_211 : brIdx_26;
  assign GEN_426 = r_btb_update_valid ? GEN_212 : brIdx_27;
  assign GEN_427 = r_btb_update_valid ? GEN_213 : brIdx_28;
  assign GEN_428 = r_btb_update_valid ? GEN_214 : brIdx_29;
  assign GEN_429 = r_btb_update_valid ? GEN_215 : brIdx_30;
  assign GEN_430 = r_btb_update_valid ? GEN_216 : brIdx_31;
  assign GEN_431 = r_btb_update_valid ? GEN_217 : brIdx_32;
  assign GEN_432 = r_btb_update_valid ? GEN_218 : brIdx_33;
  assign GEN_433 = r_btb_update_valid ? GEN_219 : brIdx_34;
  assign GEN_434 = r_btb_update_valid ? GEN_220 : brIdx_35;
  assign GEN_435 = r_btb_update_valid ? GEN_221 : brIdx_36;
  assign GEN_436 = r_btb_update_valid ? GEN_222 : brIdx_37;
  assign GEN_437 = r_btb_update_valid ? GEN_223 : brIdx_38;
  assign GEN_438 = r_btb_update_valid ? GEN_224 : brIdx_39;
  assign GEN_439 = r_btb_update_valid ? GEN_225 : pages_0;
  assign GEN_440 = r_btb_update_valid ? GEN_226 : pages_2;
  assign GEN_441 = r_btb_update_valid ? GEN_227 : pages_4;
  assign GEN_442 = r_btb_update_valid ? GEN_228 : pages_1;
  assign GEN_443 = r_btb_update_valid ? GEN_229 : pages_3;
  assign GEN_444 = r_btb_update_valid ? GEN_230 : pages_5;
  assign GEN_445 = r_btb_update_valid ? T_1651 : {{2'd0}, pageValid};
  assign T_1653 = hitsVec != 40'h0;
  assign T_1655 = hitsVec[0];
  assign T_1656 = hitsVec[1];
  assign T_1657 = hitsVec[2];
  assign T_1658 = hitsVec[3];
  assign T_1659 = hitsVec[4];
  assign T_1660 = hitsVec[5];
  assign T_1661 = hitsVec[6];
  assign T_1662 = hitsVec[7];
  assign T_1663 = hitsVec[8];
  assign T_1664 = hitsVec[9];
  assign T_1665 = hitsVec[10];
  assign T_1666 = hitsVec[11];
  assign T_1667 = hitsVec[12];
  assign T_1668 = hitsVec[13];
  assign T_1669 = hitsVec[14];
  assign T_1670 = hitsVec[15];
  assign T_1671 = hitsVec[16];
  assign T_1672 = hitsVec[17];
  assign T_1673 = hitsVec[18];
  assign T_1674 = hitsVec[19];
  assign T_1675 = hitsVec[20];
  assign T_1676 = hitsVec[21];
  assign T_1677 = hitsVec[22];
  assign T_1678 = hitsVec[23];
  assign T_1679 = hitsVec[24];
  assign T_1680 = hitsVec[25];
  assign T_1681 = hitsVec[26];
  assign T_1682 = hitsVec[27];
  assign T_1683 = hitsVec[28];
  assign T_1684 = hitsVec[29];
  assign T_1685 = hitsVec[30];
  assign T_1686 = hitsVec[31];
  assign T_1687 = hitsVec[32];
  assign T_1688 = hitsVec[33];
  assign T_1689 = hitsVec[34];
  assign T_1690 = hitsVec[35];
  assign T_1691 = hitsVec[36];
  assign T_1692 = hitsVec[37];
  assign T_1693 = hitsVec[38];
  assign T_1694 = hitsVec[39];
  assign T_1696 = T_1655 ? tgtPagesOH_0 : 6'h0;
  assign T_1698 = T_1656 ? tgtPagesOH_1 : 6'h0;
  assign T_1700 = T_1657 ? tgtPagesOH_2 : 6'h0;
  assign T_1702 = T_1658 ? tgtPagesOH_3 : 6'h0;
  assign T_1704 = T_1659 ? tgtPagesOH_4 : 6'h0;
  assign T_1706 = T_1660 ? tgtPagesOH_5 : 6'h0;
  assign T_1708 = T_1661 ? tgtPagesOH_6 : 6'h0;
  assign T_1710 = T_1662 ? tgtPagesOH_7 : 6'h0;
  assign T_1712 = T_1663 ? tgtPagesOH_8 : 6'h0;
  assign T_1714 = T_1664 ? tgtPagesOH_9 : 6'h0;
  assign T_1716 = T_1665 ? tgtPagesOH_10 : 6'h0;
  assign T_1718 = T_1666 ? tgtPagesOH_11 : 6'h0;
  assign T_1720 = T_1667 ? tgtPagesOH_12 : 6'h0;
  assign T_1722 = T_1668 ? tgtPagesOH_13 : 6'h0;
  assign T_1724 = T_1669 ? tgtPagesOH_14 : 6'h0;
  assign T_1726 = T_1670 ? tgtPagesOH_15 : 6'h0;
  assign T_1728 = T_1671 ? tgtPagesOH_16 : 6'h0;
  assign T_1730 = T_1672 ? tgtPagesOH_17 : 6'h0;
  assign T_1732 = T_1673 ? tgtPagesOH_18 : 6'h0;
  assign T_1734 = T_1674 ? tgtPagesOH_19 : 6'h0;
  assign T_1736 = T_1675 ? tgtPagesOH_20 : 6'h0;
  assign T_1738 = T_1676 ? tgtPagesOH_21 : 6'h0;
  assign T_1740 = T_1677 ? tgtPagesOH_22 : 6'h0;
  assign T_1742 = T_1678 ? tgtPagesOH_23 : 6'h0;
  assign T_1744 = T_1679 ? tgtPagesOH_24 : 6'h0;
  assign T_1746 = T_1680 ? tgtPagesOH_25 : 6'h0;
  assign T_1748 = T_1681 ? tgtPagesOH_26 : 6'h0;
  assign T_1750 = T_1682 ? tgtPagesOH_27 : 6'h0;
  assign T_1752 = T_1683 ? tgtPagesOH_28 : 6'h0;
  assign T_1754 = T_1684 ? tgtPagesOH_29 : 6'h0;
  assign T_1756 = T_1685 ? tgtPagesOH_30 : 6'h0;
  assign T_1758 = T_1686 ? tgtPagesOH_31 : 6'h0;
  assign T_1760 = T_1687 ? tgtPagesOH_32 : 6'h0;
  assign T_1762 = T_1688 ? tgtPagesOH_33 : 6'h0;
  assign T_1764 = T_1689 ? tgtPagesOH_34 : 6'h0;
  assign T_1766 = T_1690 ? tgtPagesOH_35 : 6'h0;
  assign T_1768 = T_1691 ? tgtPagesOH_36 : 6'h0;
  assign T_1770 = T_1692 ? tgtPagesOH_37 : 6'h0;
  assign T_1772 = T_1693 ? tgtPagesOH_38 : 6'h0;
  assign T_1774 = T_1694 ? tgtPagesOH_39 : 6'h0;
  assign T_1776 = T_1696 | T_1698;
  assign T_1777 = T_1776 | T_1700;
  assign T_1778 = T_1777 | T_1702;
  assign T_1779 = T_1778 | T_1704;
  assign T_1780 = T_1779 | T_1706;
  assign T_1781 = T_1780 | T_1708;
  assign T_1782 = T_1781 | T_1710;
  assign T_1783 = T_1782 | T_1712;
  assign T_1784 = T_1783 | T_1714;
  assign T_1785 = T_1784 | T_1716;
  assign T_1786 = T_1785 | T_1718;
  assign T_1787 = T_1786 | T_1720;
  assign T_1788 = T_1787 | T_1722;
  assign T_1789 = T_1788 | T_1724;
  assign T_1790 = T_1789 | T_1726;
  assign T_1791 = T_1790 | T_1728;
  assign T_1792 = T_1791 | T_1730;
  assign T_1793 = T_1792 | T_1732;
  assign T_1794 = T_1793 | T_1734;
  assign T_1795 = T_1794 | T_1736;
  assign T_1796 = T_1795 | T_1738;
  assign T_1797 = T_1796 | T_1740;
  assign T_1798 = T_1797 | T_1742;
  assign T_1799 = T_1798 | T_1744;
  assign T_1800 = T_1799 | T_1746;
  assign T_1801 = T_1800 | T_1748;
  assign T_1802 = T_1801 | T_1750;
  assign T_1803 = T_1802 | T_1752;
  assign T_1804 = T_1803 | T_1754;
  assign T_1805 = T_1804 | T_1756;
  assign T_1806 = T_1805 | T_1758;
  assign T_1807 = T_1806 | T_1760;
  assign T_1808 = T_1807 | T_1762;
  assign T_1809 = T_1808 | T_1764;
  assign T_1810 = T_1809 | T_1766;
  assign T_1811 = T_1810 | T_1768;
  assign T_1812 = T_1811 | T_1770;
  assign T_1813 = T_1812 | T_1772;
  assign T_1814 = T_1813 | T_1774;
  assign T_1815 = T_1814;
  assign T_1816 = T_1815[0];
  assign T_1817 = T_1815[1];
  assign T_1818 = T_1815[2];
  assign T_1819 = T_1815[3];
  assign T_1820 = T_1815[4];
  assign T_1821 = T_1815[5];
  assign T_1823 = T_1816 ? pages_0 : 27'h0;
  assign T_1825 = T_1817 ? pages_1 : 27'h0;
  assign T_1827 = T_1818 ? pages_2 : 27'h0;
  assign T_1829 = T_1819 ? pages_3 : 27'h0;
  assign T_1831 = T_1820 ? pages_4 : 27'h0;
  assign T_1833 = T_1821 ? pages_5 : 27'h0;
  assign T_1835 = T_1823 | T_1825;
  assign T_1836 = T_1835 | T_1827;
  assign T_1837 = T_1836 | T_1829;
  assign T_1838 = T_1837 | T_1831;
  assign T_1839 = T_1838 | T_1833;
  assign T_1840 = T_1839;
  assign T_1882 = T_1655 ? tgts_0 : 11'h0;
  assign T_1884 = T_1656 ? tgts_1 : 11'h0;
  assign T_1886 = T_1657 ? tgts_2 : 11'h0;
  assign T_1888 = T_1658 ? tgts_3 : 11'h0;
  assign T_1890 = T_1659 ? tgts_4 : 11'h0;
  assign T_1892 = T_1660 ? tgts_5 : 11'h0;
  assign T_1894 = T_1661 ? tgts_6 : 11'h0;
  assign T_1896 = T_1662 ? tgts_7 : 11'h0;
  assign T_1898 = T_1663 ? tgts_8 : 11'h0;
  assign T_1900 = T_1664 ? tgts_9 : 11'h0;
  assign T_1902 = T_1665 ? tgts_10 : 11'h0;
  assign T_1904 = T_1666 ? tgts_11 : 11'h0;
  assign T_1906 = T_1667 ? tgts_12 : 11'h0;
  assign T_1908 = T_1668 ? tgts_13 : 11'h0;
  assign T_1910 = T_1669 ? tgts_14 : 11'h0;
  assign T_1912 = T_1670 ? tgts_15 : 11'h0;
  assign T_1914 = T_1671 ? tgts_16 : 11'h0;
  assign T_1916 = T_1672 ? tgts_17 : 11'h0;
  assign T_1918 = T_1673 ? tgts_18 : 11'h0;
  assign T_1920 = T_1674 ? tgts_19 : 11'h0;
  assign T_1922 = T_1675 ? tgts_20 : 11'h0;
  assign T_1924 = T_1676 ? tgts_21 : 11'h0;
  assign T_1926 = T_1677 ? tgts_22 : 11'h0;
  assign T_1928 = T_1678 ? tgts_23 : 11'h0;
  assign T_1930 = T_1679 ? tgts_24 : 11'h0;
  assign T_1932 = T_1680 ? tgts_25 : 11'h0;
  assign T_1934 = T_1681 ? tgts_26 : 11'h0;
  assign T_1936 = T_1682 ? tgts_27 : 11'h0;
  assign T_1938 = T_1683 ? tgts_28 : 11'h0;
  assign T_1940 = T_1684 ? tgts_29 : 11'h0;
  assign T_1942 = T_1685 ? tgts_30 : 11'h0;
  assign T_1944 = T_1686 ? tgts_31 : 11'h0;
  assign T_1946 = T_1687 ? tgts_32 : 11'h0;
  assign T_1948 = T_1688 ? tgts_33 : 11'h0;
  assign T_1950 = T_1689 ? tgts_34 : 11'h0;
  assign T_1952 = T_1690 ? tgts_35 : 11'h0;
  assign T_1954 = T_1691 ? tgts_36 : 11'h0;
  assign T_1956 = T_1692 ? tgts_37 : 11'h0;
  assign T_1958 = T_1693 ? tgts_38 : 11'h0;
  assign T_1960 = T_1694 ? tgts_39 : 11'h0;
  assign T_1962 = T_1882 | T_1884;
  assign T_1963 = T_1962 | T_1886;
  assign T_1964 = T_1963 | T_1888;
  assign T_1965 = T_1964 | T_1890;
  assign T_1966 = T_1965 | T_1892;
  assign T_1967 = T_1966 | T_1894;
  assign T_1968 = T_1967 | T_1896;
  assign T_1969 = T_1968 | T_1898;
  assign T_1970 = T_1969 | T_1900;
  assign T_1971 = T_1970 | T_1902;
  assign T_1972 = T_1971 | T_1904;
  assign T_1973 = T_1972 | T_1906;
  assign T_1974 = T_1973 | T_1908;
  assign T_1975 = T_1974 | T_1910;
  assign T_1976 = T_1975 | T_1912;
  assign T_1977 = T_1976 | T_1914;
  assign T_1978 = T_1977 | T_1916;
  assign T_1979 = T_1978 | T_1918;
  assign T_1980 = T_1979 | T_1920;
  assign T_1981 = T_1980 | T_1922;
  assign T_1982 = T_1981 | T_1924;
  assign T_1983 = T_1982 | T_1926;
  assign T_1984 = T_1983 | T_1928;
  assign T_1985 = T_1984 | T_1930;
  assign T_1986 = T_1985 | T_1932;
  assign T_1987 = T_1986 | T_1934;
  assign T_1988 = T_1987 | T_1936;
  assign T_1989 = T_1988 | T_1938;
  assign T_1990 = T_1989 | T_1940;
  assign T_1991 = T_1990 | T_1942;
  assign T_1992 = T_1991 | T_1944;
  assign T_1993 = T_1992 | T_1946;
  assign T_1994 = T_1993 | T_1948;
  assign T_1995 = T_1994 | T_1950;
  assign T_1996 = T_1995 | T_1952;
  assign T_1997 = T_1996 | T_1954;
  assign T_1998 = T_1997 | T_1956;
  assign T_1999 = T_1998 | T_1958;
  assign T_2000 = T_1999 | T_1960;
  assign T_2001 = T_2000;
  assign GEN_486 = {{1'd0}, T_2001};
  assign T_2002 = GEN_486 << 1;
  assign T_2003 = {T_1840,T_2002};
  assign T_2004 = hitsVec[39:32];
  assign T_2005 = hitsVec[31:0];
  assign T_2007 = T_2004 != 8'h0;
  assign GEN_487 = {{24'd0}, T_2004};
  assign T_2008 = GEN_487 | T_2005;
  assign T_2009 = T_2008[31:16];
  assign T_2010 = T_2008[15:0];
  assign T_2012 = T_2009 != 16'h0;
  assign T_2013 = T_2009 | T_2010;
  assign T_2014 = T_2013[15:8];
  assign T_2015 = T_2013[7:0];
  assign T_2017 = T_2014 != 8'h0;
  assign T_2018 = T_2014 | T_2015;
  assign T_2019 = T_2018[7:4];
  assign T_2020 = T_2018[3:0];
  assign T_2022 = T_2019 != 4'h0;
  assign T_2023 = T_2019 | T_2020;
  assign T_2024 = T_2023[3:2];
  assign T_2025 = T_2023[1:0];
  assign T_2027 = T_2024 != 2'h0;
  assign T_2028 = T_2024 | T_2025;
  assign T_2029 = T_2028[1];
  assign T_2030 = {T_2027,T_2029};
  assign T_2031 = {T_2022,T_2030};
  assign T_2032 = {T_2017,T_2031};
  assign T_2033 = {T_2012,T_2032};
  assign T_2034 = {T_2007,T_2033};
  assign T_2076 = T_1655 ? brIdx_0 : 1'h0;
  assign T_2078 = T_1656 ? brIdx_1 : 1'h0;
  assign T_2080 = T_1657 ? brIdx_2 : 1'h0;
  assign T_2082 = T_1658 ? brIdx_3 : 1'h0;
  assign T_2084 = T_1659 ? brIdx_4 : 1'h0;
  assign T_2086 = T_1660 ? brIdx_5 : 1'h0;
  assign T_2088 = T_1661 ? brIdx_6 : 1'h0;
  assign T_2090 = T_1662 ? brIdx_7 : 1'h0;
  assign T_2092 = T_1663 ? brIdx_8 : 1'h0;
  assign T_2094 = T_1664 ? brIdx_9 : 1'h0;
  assign T_2096 = T_1665 ? brIdx_10 : 1'h0;
  assign T_2098 = T_1666 ? brIdx_11 : 1'h0;
  assign T_2100 = T_1667 ? brIdx_12 : 1'h0;
  assign T_2102 = T_1668 ? brIdx_13 : 1'h0;
  assign T_2104 = T_1669 ? brIdx_14 : 1'h0;
  assign T_2106 = T_1670 ? brIdx_15 : 1'h0;
  assign T_2108 = T_1671 ? brIdx_16 : 1'h0;
  assign T_2110 = T_1672 ? brIdx_17 : 1'h0;
  assign T_2112 = T_1673 ? brIdx_18 : 1'h0;
  assign T_2114 = T_1674 ? brIdx_19 : 1'h0;
  assign T_2116 = T_1675 ? brIdx_20 : 1'h0;
  assign T_2118 = T_1676 ? brIdx_21 : 1'h0;
  assign T_2120 = T_1677 ? brIdx_22 : 1'h0;
  assign T_2122 = T_1678 ? brIdx_23 : 1'h0;
  assign T_2124 = T_1679 ? brIdx_24 : 1'h0;
  assign T_2126 = T_1680 ? brIdx_25 : 1'h0;
  assign T_2128 = T_1681 ? brIdx_26 : 1'h0;
  assign T_2130 = T_1682 ? brIdx_27 : 1'h0;
  assign T_2132 = T_1683 ? brIdx_28 : 1'h0;
  assign T_2134 = T_1684 ? brIdx_29 : 1'h0;
  assign T_2136 = T_1685 ? brIdx_30 : 1'h0;
  assign T_2138 = T_1686 ? brIdx_31 : 1'h0;
  assign T_2140 = T_1687 ? brIdx_32 : 1'h0;
  assign T_2142 = T_1688 ? brIdx_33 : 1'h0;
  assign T_2144 = T_1689 ? brIdx_34 : 1'h0;
  assign T_2146 = T_1690 ? brIdx_35 : 1'h0;
  assign T_2148 = T_1691 ? brIdx_36 : 1'h0;
  assign T_2150 = T_1692 ? brIdx_37 : 1'h0;
  assign T_2152 = T_1693 ? brIdx_38 : 1'h0;
  assign T_2154 = T_1694 ? brIdx_39 : 1'h0;
  assign T_2156 = T_2076 | T_2078;
  assign T_2157 = T_2156 | T_2080;
  assign T_2158 = T_2157 | T_2082;
  assign T_2159 = T_2158 | T_2084;
  assign T_2160 = T_2159 | T_2086;
  assign T_2161 = T_2160 | T_2088;
  assign T_2162 = T_2161 | T_2090;
  assign T_2163 = T_2162 | T_2092;
  assign T_2164 = T_2163 | T_2094;
  assign T_2165 = T_2164 | T_2096;
  assign T_2166 = T_2165 | T_2098;
  assign T_2167 = T_2166 | T_2100;
  assign T_2168 = T_2167 | T_2102;
  assign T_2169 = T_2168 | T_2104;
  assign T_2170 = T_2169 | T_2106;
  assign T_2171 = T_2170 | T_2108;
  assign T_2172 = T_2171 | T_2110;
  assign T_2173 = T_2172 | T_2112;
  assign T_2174 = T_2173 | T_2114;
  assign T_2175 = T_2174 | T_2116;
  assign T_2176 = T_2175 | T_2118;
  assign T_2177 = T_2176 | T_2120;
  assign T_2178 = T_2177 | T_2122;
  assign T_2179 = T_2178 | T_2124;
  assign T_2180 = T_2179 | T_2126;
  assign T_2181 = T_2180 | T_2128;
  assign T_2182 = T_2181 | T_2130;
  assign T_2183 = T_2182 | T_2132;
  assign T_2184 = T_2183 | T_2134;
  assign T_2185 = T_2184 | T_2136;
  assign T_2186 = T_2185 | T_2138;
  assign T_2187 = T_2186 | T_2140;
  assign T_2188 = T_2187 | T_2142;
  assign T_2189 = T_2188 | T_2144;
  assign T_2190 = T_2189 | T_2146;
  assign T_2191 = T_2190 | T_2148;
  assign T_2192 = T_2191 | T_2150;
  assign T_2193 = T_2192 | T_2152;
  assign T_2194 = T_2193 | T_2154;
  assign T_2195 = T_2194;
  assign T_2197 = ~ io_resp_bits_bridx;
  assign T_2199 = io_resp_bits_taken ? T_2197 : 1'h0;
  assign T_2200 = ~ T_2199;
  assign T_2201 = 2'h1 << T_2200;
  assign T_2203 = T_2201 - 2'h1;
  assign T_2204 = T_2203[1:0];
  assign T_2206 = {T_2204,1'h1};
  assign T_2209_T_2227_addr = T_2226[6:0];
  assign T_2209_T_2227_en = 1'h1;
  assign T_2209_T_2227_data = T_2209[T_2209_T_2227_addr];
  assign T_2209_T_2234_data = T_2243;
  assign T_2209_T_2234_addr = T_2233[6:0];
  assign T_2209_T_2234_mask = T_2231;
  assign T_2209_T_2234_en = T_2231;
  assign T_2212 = hitsVec & isJump;
  assign T_2214 = T_2212 != 40'h0;
  assign T_2216 = T_2214 == 1'h0;
  assign T_2217 = io_req_valid & io_resp_valid;
  assign T_2218 = T_2217 & T_2216;
  assign T_2222_history = T_2211;
  assign T_2222_value = T_2209_T_2227_data;
  assign T_2225 = io_req_bits_addr[8:1];
  assign GEN_488 = {{1'd0}, T_2211};
  assign T_2226 = T_2225 ^ GEN_488;
  assign T_2228 = T_2222_value[0];
  assign T_2229 = T_2211[6:1];
  assign T_2230 = {T_2228,T_2229};
  assign GEN_446 = T_2218 ? T_2230 : T_2211;
  assign T_2231 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T_2232 = io_bht_update_bits_pc[8:1];
  assign GEN_489 = {{1'd0}, io_bht_update_bits_prediction_bits_bht_history};
  assign T_2233 = T_2232 ^ GEN_489;
  assign T_2235 = io_bht_update_bits_prediction_bits_bht_value[1];
  assign T_2236 = io_bht_update_bits_prediction_bits_bht_value[0];
  assign T_2237 = T_2235 & T_2236;
  assign T_2240 = T_2235 | T_2236;
  assign T_2241 = T_2240 & io_bht_update_bits_taken;
  assign T_2242 = T_2237 | T_2241;
  assign T_2243 = {io_bht_update_bits_taken,T_2242};
  assign T_2244 = io_bht_update_bits_prediction_bits_bht_history[6:1];
  assign T_2245 = {io_bht_update_bits_taken,T_2244};
  assign GEN_447 = io_bht_update_bits_mispredict ? T_2245 : GEN_446;
  assign GEN_453 = T_2231 ? GEN_447 : GEN_446;
  assign T_2248 = T_2228 == 1'h0;
  assign T_2249 = T_2248 & T_2216;
  assign GEN_454 = T_2249 ? 1'h0 : 1'h1;
  assign T_2263 = hitsVec & isReturn;
  assign T_2265 = T_2263 != 40'h0;
  assign T_2267 = T_2252 == 2'h0;
  assign T_2269 = T_2267 == 1'h0;
  assign T_2270 = T_2269 & T_2265;
  assign GEN_5 = GEN_455;
  assign GEN_455 = T_2254 ? T_2261_1 : T_2261_0;
  assign GEN_457 = T_2270 ? GEN_5 : T_2003;
  assign T_2272 = T_2252 < 2'h2;
  assign T_2274 = T_2252 + 2'h1;
  assign T_2275 = T_2274[1:0];
  assign GEN_458 = T_2272 ? T_2275 : T_2252;
  assign T_2281 = T_2254 + 1'h1;
  assign T_2282 = T_2281[0:0];
  assign GEN_6 = io_ras_update_bits_returnAddr;
  assign GEN_459 = 1'h0 == T_2282 ? GEN_6 : T_2261_0;
  assign GEN_460 = T_2282 ? GEN_6 : T_2261_1;
  assign GEN_461 = T_2265 ? io_ras_update_bits_returnAddr : GEN_457;
  assign GEN_462 = io_ras_update_bits_isCall ? GEN_458 : T_2252;
  assign GEN_464 = io_ras_update_bits_isCall ? GEN_459 : T_2261_0;
  assign GEN_465 = io_ras_update_bits_isCall ? GEN_460 : T_2261_1;
  assign GEN_466 = io_ras_update_bits_isCall ? T_2282 : T_2254;
  assign GEN_467 = io_ras_update_bits_isCall ? GEN_461 : GEN_457;
  assign T_2285 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T_2287 = io_ras_update_bits_isCall == 1'h0;
  assign T_2288 = T_2287 & T_2285;
  assign T_2294 = T_2252 - 2'h1;
  assign T_2295 = T_2294[1:0];
  assign T_2301 = T_2254 - 1'h1;
  assign T_2302 = T_2301[0:0];
  assign GEN_468 = T_2269 ? T_2295 : GEN_462;
  assign GEN_469 = T_2269 ? T_2302 : GEN_466;
  assign GEN_470 = T_2288 ? GEN_468 : GEN_462;
  assign GEN_471 = T_2288 ? GEN_469 : GEN_466;
  assign GEN_472 = io_ras_update_valid ? GEN_470 : T_2252;
  assign GEN_474 = io_ras_update_valid ? GEN_464 : T_2261_0;
  assign GEN_475 = io_ras_update_valid ? GEN_465 : T_2261_1;
  assign GEN_476 = io_ras_update_valid ? GEN_471 : T_2254;
  assign GEN_477 = io_ras_update_valid ? GEN_467 : GEN_457;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_231 = {1{$random}};
  idxs_0 = GEN_231[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_272 = {1{$random}};
  idxs_1 = GEN_272[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_313 = {1{$random}};
  idxs_2 = GEN_313[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_354 = {1{$random}};
  idxs_3 = GEN_354[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_398 = {1{$random}};
  idxs_4 = GEN_398[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_448 = {1{$random}};
  idxs_5 = GEN_448[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_449 = {1{$random}};
  idxs_6 = GEN_449[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_450 = {1{$random}};
  idxs_7 = GEN_450[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_451 = {1{$random}};
  idxs_8 = GEN_451[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_452 = {1{$random}};
  idxs_9 = GEN_452[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_456 = {1{$random}};
  idxs_10 = GEN_456[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_463 = {1{$random}};
  idxs_11 = GEN_463[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_473 = {1{$random}};
  idxs_12 = GEN_473[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_480 = {1{$random}};
  idxs_13 = GEN_480[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_482 = {1{$random}};
  idxs_14 = GEN_482[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_484 = {1{$random}};
  idxs_15 = GEN_484[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_490 = {1{$random}};
  idxs_16 = GEN_490[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_491 = {1{$random}};
  idxs_17 = GEN_491[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_492 = {1{$random}};
  idxs_18 = GEN_492[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_493 = {1{$random}};
  idxs_19 = GEN_493[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_494 = {1{$random}};
  idxs_20 = GEN_494[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_495 = {1{$random}};
  idxs_21 = GEN_495[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_496 = {1{$random}};
  idxs_22 = GEN_496[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_497 = {1{$random}};
  idxs_23 = GEN_497[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_498 = {1{$random}};
  idxs_24 = GEN_498[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_499 = {1{$random}};
  idxs_25 = GEN_499[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_500 = {1{$random}};
  idxs_26 = GEN_500[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_501 = {1{$random}};
  idxs_27 = GEN_501[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_502 = {1{$random}};
  idxs_28 = GEN_502[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_503 = {1{$random}};
  idxs_29 = GEN_503[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_504 = {1{$random}};
  idxs_30 = GEN_504[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_505 = {1{$random}};
  idxs_31 = GEN_505[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_506 = {1{$random}};
  idxs_32 = GEN_506[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_507 = {1{$random}};
  idxs_33 = GEN_507[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_508 = {1{$random}};
  idxs_34 = GEN_508[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_509 = {1{$random}};
  idxs_35 = GEN_509[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_510 = {1{$random}};
  idxs_36 = GEN_510[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_511 = {1{$random}};
  idxs_37 = GEN_511[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_512 = {1{$random}};
  idxs_38 = GEN_512[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_513 = {1{$random}};
  idxs_39 = GEN_513[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_514 = {1{$random}};
  idxPages_0 = GEN_514[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_515 = {1{$random}};
  idxPages_1 = GEN_515[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_516 = {1{$random}};
  idxPages_2 = GEN_516[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_517 = {1{$random}};
  idxPages_3 = GEN_517[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_518 = {1{$random}};
  idxPages_4 = GEN_518[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_519 = {1{$random}};
  idxPages_5 = GEN_519[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_520 = {1{$random}};
  idxPages_6 = GEN_520[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_521 = {1{$random}};
  idxPages_7 = GEN_521[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_522 = {1{$random}};
  idxPages_8 = GEN_522[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_523 = {1{$random}};
  idxPages_9 = GEN_523[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_524 = {1{$random}};
  idxPages_10 = GEN_524[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_525 = {1{$random}};
  idxPages_11 = GEN_525[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_526 = {1{$random}};
  idxPages_12 = GEN_526[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_527 = {1{$random}};
  idxPages_13 = GEN_527[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_528 = {1{$random}};
  idxPages_14 = GEN_528[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_529 = {1{$random}};
  idxPages_15 = GEN_529[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_530 = {1{$random}};
  idxPages_16 = GEN_530[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_531 = {1{$random}};
  idxPages_17 = GEN_531[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_532 = {1{$random}};
  idxPages_18 = GEN_532[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_533 = {1{$random}};
  idxPages_19 = GEN_533[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_534 = {1{$random}};
  idxPages_20 = GEN_534[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_535 = {1{$random}};
  idxPages_21 = GEN_535[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_536 = {1{$random}};
  idxPages_22 = GEN_536[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_537 = {1{$random}};
  idxPages_23 = GEN_537[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_538 = {1{$random}};
  idxPages_24 = GEN_538[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_539 = {1{$random}};
  idxPages_25 = GEN_539[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_540 = {1{$random}};
  idxPages_26 = GEN_540[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_541 = {1{$random}};
  idxPages_27 = GEN_541[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_542 = {1{$random}};
  idxPages_28 = GEN_542[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_543 = {1{$random}};
  idxPages_29 = GEN_543[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_544 = {1{$random}};
  idxPages_30 = GEN_544[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_545 = {1{$random}};
  idxPages_31 = GEN_545[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_546 = {1{$random}};
  idxPages_32 = GEN_546[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_547 = {1{$random}};
  idxPages_33 = GEN_547[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_548 = {1{$random}};
  idxPages_34 = GEN_548[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_549 = {1{$random}};
  idxPages_35 = GEN_549[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_550 = {1{$random}};
  idxPages_36 = GEN_550[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_551 = {1{$random}};
  idxPages_37 = GEN_551[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_552 = {1{$random}};
  idxPages_38 = GEN_552[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_553 = {1{$random}};
  idxPages_39 = GEN_553[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_554 = {1{$random}};
  tgts_0 = GEN_554[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_555 = {1{$random}};
  tgts_1 = GEN_555[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_556 = {1{$random}};
  tgts_2 = GEN_556[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_557 = {1{$random}};
  tgts_3 = GEN_557[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_558 = {1{$random}};
  tgts_4 = GEN_558[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_559 = {1{$random}};
  tgts_5 = GEN_559[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_560 = {1{$random}};
  tgts_6 = GEN_560[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_561 = {1{$random}};
  tgts_7 = GEN_561[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_562 = {1{$random}};
  tgts_8 = GEN_562[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_563 = {1{$random}};
  tgts_9 = GEN_563[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_564 = {1{$random}};
  tgts_10 = GEN_564[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_565 = {1{$random}};
  tgts_11 = GEN_565[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_566 = {1{$random}};
  tgts_12 = GEN_566[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_567 = {1{$random}};
  tgts_13 = GEN_567[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_568 = {1{$random}};
  tgts_14 = GEN_568[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_569 = {1{$random}};
  tgts_15 = GEN_569[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_570 = {1{$random}};
  tgts_16 = GEN_570[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_571 = {1{$random}};
  tgts_17 = GEN_571[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_572 = {1{$random}};
  tgts_18 = GEN_572[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_573 = {1{$random}};
  tgts_19 = GEN_573[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_574 = {1{$random}};
  tgts_20 = GEN_574[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_575 = {1{$random}};
  tgts_21 = GEN_575[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_576 = {1{$random}};
  tgts_22 = GEN_576[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_577 = {1{$random}};
  tgts_23 = GEN_577[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_578 = {1{$random}};
  tgts_24 = GEN_578[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_579 = {1{$random}};
  tgts_25 = GEN_579[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_580 = {1{$random}};
  tgts_26 = GEN_580[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_581 = {1{$random}};
  tgts_27 = GEN_581[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_582 = {1{$random}};
  tgts_28 = GEN_582[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_583 = {1{$random}};
  tgts_29 = GEN_583[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_584 = {1{$random}};
  tgts_30 = GEN_584[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_585 = {1{$random}};
  tgts_31 = GEN_585[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_586 = {1{$random}};
  tgts_32 = GEN_586[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_587 = {1{$random}};
  tgts_33 = GEN_587[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_588 = {1{$random}};
  tgts_34 = GEN_588[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_589 = {1{$random}};
  tgts_35 = GEN_589[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_590 = {1{$random}};
  tgts_36 = GEN_590[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_591 = {1{$random}};
  tgts_37 = GEN_591[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_592 = {1{$random}};
  tgts_38 = GEN_592[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_593 = {1{$random}};
  tgts_39 = GEN_593[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_594 = {1{$random}};
  tgtPages_0 = GEN_594[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_595 = {1{$random}};
  tgtPages_1 = GEN_595[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_596 = {1{$random}};
  tgtPages_2 = GEN_596[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_597 = {1{$random}};
  tgtPages_3 = GEN_597[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_598 = {1{$random}};
  tgtPages_4 = GEN_598[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_599 = {1{$random}};
  tgtPages_5 = GEN_599[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_600 = {1{$random}};
  tgtPages_6 = GEN_600[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_601 = {1{$random}};
  tgtPages_7 = GEN_601[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_602 = {1{$random}};
  tgtPages_8 = GEN_602[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_603 = {1{$random}};
  tgtPages_9 = GEN_603[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_604 = {1{$random}};
  tgtPages_10 = GEN_604[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_605 = {1{$random}};
  tgtPages_11 = GEN_605[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_606 = {1{$random}};
  tgtPages_12 = GEN_606[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_607 = {1{$random}};
  tgtPages_13 = GEN_607[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_608 = {1{$random}};
  tgtPages_14 = GEN_608[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_609 = {1{$random}};
  tgtPages_15 = GEN_609[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_610 = {1{$random}};
  tgtPages_16 = GEN_610[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_611 = {1{$random}};
  tgtPages_17 = GEN_611[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_612 = {1{$random}};
  tgtPages_18 = GEN_612[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_613 = {1{$random}};
  tgtPages_19 = GEN_613[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_614 = {1{$random}};
  tgtPages_20 = GEN_614[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_615 = {1{$random}};
  tgtPages_21 = GEN_615[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_616 = {1{$random}};
  tgtPages_22 = GEN_616[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_617 = {1{$random}};
  tgtPages_23 = GEN_617[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_618 = {1{$random}};
  tgtPages_24 = GEN_618[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_619 = {1{$random}};
  tgtPages_25 = GEN_619[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_620 = {1{$random}};
  tgtPages_26 = GEN_620[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_621 = {1{$random}};
  tgtPages_27 = GEN_621[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_622 = {1{$random}};
  tgtPages_28 = GEN_622[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_623 = {1{$random}};
  tgtPages_29 = GEN_623[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_624 = {1{$random}};
  tgtPages_30 = GEN_624[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_625 = {1{$random}};
  tgtPages_31 = GEN_625[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_626 = {1{$random}};
  tgtPages_32 = GEN_626[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_627 = {1{$random}};
  tgtPages_33 = GEN_627[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_628 = {1{$random}};
  tgtPages_34 = GEN_628[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_629 = {1{$random}};
  tgtPages_35 = GEN_629[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_630 = {1{$random}};
  tgtPages_36 = GEN_630[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_631 = {1{$random}};
  tgtPages_37 = GEN_631[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_632 = {1{$random}};
  tgtPages_38 = GEN_632[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_633 = {1{$random}};
  tgtPages_39 = GEN_633[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_634 = {1{$random}};
  pages_0 = GEN_634[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_635 = {1{$random}};
  pages_1 = GEN_635[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_636 = {1{$random}};
  pages_2 = GEN_636[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_637 = {1{$random}};
  pages_3 = GEN_637[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_638 = {1{$random}};
  pages_4 = GEN_638[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_639 = {1{$random}};
  pages_5 = GEN_639[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_640 = {1{$random}};
  pageValid = GEN_640[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_641 = {2{$random}};
  isValid = GEN_641[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_642 = {2{$random}};
  isReturn = GEN_642[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_643 = {2{$random}};
  isJump = GEN_643[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_644 = {1{$random}};
  brIdx_0 = GEN_644[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_645 = {1{$random}};
  brIdx_1 = GEN_645[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_646 = {1{$random}};
  brIdx_2 = GEN_646[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_647 = {1{$random}};
  brIdx_3 = GEN_647[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_648 = {1{$random}};
  brIdx_4 = GEN_648[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_649 = {1{$random}};
  brIdx_5 = GEN_649[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_650 = {1{$random}};
  brIdx_6 = GEN_650[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_651 = {1{$random}};
  brIdx_7 = GEN_651[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_652 = {1{$random}};
  brIdx_8 = GEN_652[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_653 = {1{$random}};
  brIdx_9 = GEN_653[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_654 = {1{$random}};
  brIdx_10 = GEN_654[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_655 = {1{$random}};
  brIdx_11 = GEN_655[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_656 = {1{$random}};
  brIdx_12 = GEN_656[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_657 = {1{$random}};
  brIdx_13 = GEN_657[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_658 = {1{$random}};
  brIdx_14 = GEN_658[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_659 = {1{$random}};
  brIdx_15 = GEN_659[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_660 = {1{$random}};
  brIdx_16 = GEN_660[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_661 = {1{$random}};
  brIdx_17 = GEN_661[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_662 = {1{$random}};
  brIdx_18 = GEN_662[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_663 = {1{$random}};
  brIdx_19 = GEN_663[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_664 = {1{$random}};
  brIdx_20 = GEN_664[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_665 = {1{$random}};
  brIdx_21 = GEN_665[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_666 = {1{$random}};
  brIdx_22 = GEN_666[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_667 = {1{$random}};
  brIdx_23 = GEN_667[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_668 = {1{$random}};
  brIdx_24 = GEN_668[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_669 = {1{$random}};
  brIdx_25 = GEN_669[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_670 = {1{$random}};
  brIdx_26 = GEN_670[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_671 = {1{$random}};
  brIdx_27 = GEN_671[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_672 = {1{$random}};
  brIdx_28 = GEN_672[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_673 = {1{$random}};
  brIdx_29 = GEN_673[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_674 = {1{$random}};
  brIdx_30 = GEN_674[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_675 = {1{$random}};
  brIdx_31 = GEN_675[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_676 = {1{$random}};
  brIdx_32 = GEN_676[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_677 = {1{$random}};
  brIdx_33 = GEN_677[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_678 = {1{$random}};
  brIdx_34 = GEN_678[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_679 = {1{$random}};
  brIdx_35 = GEN_679[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_680 = {1{$random}};
  brIdx_36 = GEN_680[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_681 = {1{$random}};
  brIdx_37 = GEN_681[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_682 = {1{$random}};
  brIdx_38 = GEN_682[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_683 = {1{$random}};
  brIdx_39 = GEN_683[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_684 = {1{$random}};
  T_777 = GEN_684[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_685 = {1{$random}};
  T_778_prediction_valid = GEN_685[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_686 = {1{$random}};
  T_778_prediction_bits_taken = GEN_686[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_687 = {1{$random}};
  T_778_prediction_bits_mask = GEN_687[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_688 = {1{$random}};
  T_778_prediction_bits_bridx = GEN_688[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_689 = {2{$random}};
  T_778_prediction_bits_target = GEN_689[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_690 = {1{$random}};
  T_778_prediction_bits_entry = GEN_690[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_691 = {1{$random}};
  T_778_prediction_bits_bht_history = GEN_691[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_692 = {1{$random}};
  T_778_prediction_bits_bht_value = GEN_692[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_693 = {2{$random}};
  T_778_pc = GEN_693[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_694 = {2{$random}};
  T_778_target = GEN_694[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_695 = {1{$random}};
  T_778_taken = GEN_695[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_696 = {1{$random}};
  T_778_isValid = GEN_696[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_697 = {1{$random}};
  T_778_isJump = GEN_697[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_698 = {1{$random}};
  T_778_isReturn = GEN_698[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_699 = {2{$random}};
  T_778_br_pc = GEN_699[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_700 = {1{$random}};
  nextRepl = GEN_700[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_701 = {1{$random}};
  nextPageRepl = GEN_701[2:0];
  `endif
  GEN_702 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    T_2209[initvar] = GEN_702[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_703 = {1{$random}};
  T_2211 = GEN_703[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_704 = {1{$random}};
  T_2252 = GEN_704[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_705 = {1{$random}};
  T_2254 = GEN_705[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_706 = {2{$random}};
  T_2261_0 = GEN_706[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_707 = {2{$random}};
  T_2261_1 = GEN_707[38:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h0 == T_1615) begin
          idxs_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1 == T_1615) begin
          idxs_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2 == T_1615) begin
          idxs_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3 == T_1615) begin
          idxs_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h4 == T_1615) begin
          idxs_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h5 == T_1615) begin
          idxs_5 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h6 == T_1615) begin
          idxs_6 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h7 == T_1615) begin
          idxs_7 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h8 == T_1615) begin
          idxs_8 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h9 == T_1615) begin
          idxs_9 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'ha == T_1615) begin
          idxs_10 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hb == T_1615) begin
          idxs_11 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hc == T_1615) begin
          idxs_12 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hd == T_1615) begin
          idxs_13 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'he == T_1615) begin
          idxs_14 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hf == T_1615) begin
          idxs_15 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h10 == T_1615) begin
          idxs_16 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h11 == T_1615) begin
          idxs_17 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h12 == T_1615) begin
          idxs_18 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h13 == T_1615) begin
          idxs_19 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h14 == T_1615) begin
          idxs_20 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h15 == T_1615) begin
          idxs_21 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h16 == T_1615) begin
          idxs_22 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h17 == T_1615) begin
          idxs_23 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h18 == T_1615) begin
          idxs_24 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h19 == T_1615) begin
          idxs_25 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1a == T_1615) begin
          idxs_26 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1b == T_1615) begin
          idxs_27 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1c == T_1615) begin
          idxs_28 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1d == T_1615) begin
          idxs_29 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1e == T_1615) begin
          idxs_30 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1f == T_1615) begin
          idxs_31 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_1615) begin
          idxs_32 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_1615) begin
          idxs_33 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_1615) begin
          idxs_34 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_1615) begin
          idxs_35 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_1615) begin
          idxs_36 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_1615) begin
          idxs_37 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_1615) begin
          idxs_38 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_1615) begin
          idxs_39 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h0 == T_1615) begin
          idxPages_0 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1 == T_1615) begin
          idxPages_1 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2 == T_1615) begin
          idxPages_2 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3 == T_1615) begin
          idxPages_3 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h4 == T_1615) begin
          idxPages_4 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h5 == T_1615) begin
          idxPages_5 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h6 == T_1615) begin
          idxPages_6 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h7 == T_1615) begin
          idxPages_7 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h8 == T_1615) begin
          idxPages_8 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h9 == T_1615) begin
          idxPages_9 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'ha == T_1615) begin
          idxPages_10 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hb == T_1615) begin
          idxPages_11 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hc == T_1615) begin
          idxPages_12 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hd == T_1615) begin
          idxPages_13 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'he == T_1615) begin
          idxPages_14 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hf == T_1615) begin
          idxPages_15 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h10 == T_1615) begin
          idxPages_16 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h11 == T_1615) begin
          idxPages_17 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h12 == T_1615) begin
          idxPages_18 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h13 == T_1615) begin
          idxPages_19 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h14 == T_1615) begin
          idxPages_20 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h15 == T_1615) begin
          idxPages_21 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h16 == T_1615) begin
          idxPages_22 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h17 == T_1615) begin
          idxPages_23 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h18 == T_1615) begin
          idxPages_24 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h19 == T_1615) begin
          idxPages_25 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1a == T_1615) begin
          idxPages_26 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1b == T_1615) begin
          idxPages_27 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1c == T_1615) begin
          idxPages_28 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1d == T_1615) begin
          idxPages_29 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1e == T_1615) begin
          idxPages_30 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1f == T_1615) begin
          idxPages_31 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_1615) begin
          idxPages_32 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_1615) begin
          idxPages_33 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_1615) begin
          idxPages_34 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_1615) begin
          idxPages_35 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_1615) begin
          idxPages_36 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_1615) begin
          idxPages_37 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_1615) begin
          idxPages_38 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_1615) begin
          idxPages_39 <= GEN_2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h0 == T_1615) begin
          tgts_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1 == T_1615) begin
          tgts_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2 == T_1615) begin
          tgts_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3 == T_1615) begin
          tgts_3 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h4 == T_1615) begin
          tgts_4 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h5 == T_1615) begin
          tgts_5 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h6 == T_1615) begin
          tgts_6 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h7 == T_1615) begin
          tgts_7 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h8 == T_1615) begin
          tgts_8 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h9 == T_1615) begin
          tgts_9 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'ha == T_1615) begin
          tgts_10 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hb == T_1615) begin
          tgts_11 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hc == T_1615) begin
          tgts_12 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hd == T_1615) begin
          tgts_13 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'he == T_1615) begin
          tgts_14 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hf == T_1615) begin
          tgts_15 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h10 == T_1615) begin
          tgts_16 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h11 == T_1615) begin
          tgts_17 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h12 == T_1615) begin
          tgts_18 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h13 == T_1615) begin
          tgts_19 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h14 == T_1615) begin
          tgts_20 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h15 == T_1615) begin
          tgts_21 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h16 == T_1615) begin
          tgts_22 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h17 == T_1615) begin
          tgts_23 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h18 == T_1615) begin
          tgts_24 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h19 == T_1615) begin
          tgts_25 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1a == T_1615) begin
          tgts_26 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1b == T_1615) begin
          tgts_27 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1c == T_1615) begin
          tgts_28 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1d == T_1615) begin
          tgts_29 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1e == T_1615) begin
          tgts_30 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1f == T_1615) begin
          tgts_31 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_1615) begin
          tgts_32 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_1615) begin
          tgts_33 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_1615) begin
          tgts_34 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_1615) begin
          tgts_35 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_1615) begin
          tgts_36 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_1615) begin
          tgts_37 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_1615) begin
          tgts_38 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_1615) begin
          tgts_39 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h0 == T_1615) begin
          tgtPages_0 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1 == T_1615) begin
          tgtPages_1 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2 == T_1615) begin
          tgtPages_2 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3 == T_1615) begin
          tgtPages_3 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h4 == T_1615) begin
          tgtPages_4 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h5 == T_1615) begin
          tgtPages_5 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h6 == T_1615) begin
          tgtPages_6 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h7 == T_1615) begin
          tgtPages_7 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h8 == T_1615) begin
          tgtPages_8 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h9 == T_1615) begin
          tgtPages_9 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'ha == T_1615) begin
          tgtPages_10 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hb == T_1615) begin
          tgtPages_11 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hc == T_1615) begin
          tgtPages_12 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hd == T_1615) begin
          tgtPages_13 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'he == T_1615) begin
          tgtPages_14 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hf == T_1615) begin
          tgtPages_15 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h10 == T_1615) begin
          tgtPages_16 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h11 == T_1615) begin
          tgtPages_17 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h12 == T_1615) begin
          tgtPages_18 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h13 == T_1615) begin
          tgtPages_19 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h14 == T_1615) begin
          tgtPages_20 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h15 == T_1615) begin
          tgtPages_21 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h16 == T_1615) begin
          tgtPages_22 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h17 == T_1615) begin
          tgtPages_23 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h18 == T_1615) begin
          tgtPages_24 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h19 == T_1615) begin
          tgtPages_25 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1a == T_1615) begin
          tgtPages_26 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1b == T_1615) begin
          tgtPages_27 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1c == T_1615) begin
          tgtPages_28 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1d == T_1615) begin
          tgtPages_29 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1e == T_1615) begin
          tgtPages_30 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1f == T_1615) begin
          tgtPages_31 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_1615) begin
          tgtPages_32 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_1615) begin
          tgtPages_33 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_1615) begin
          tgtPages_34 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_1615) begin
          tgtPages_35 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_1615) begin
          tgtPages_36 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_1615) begin
          tgtPages_37 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_1615) begin
          tgtPages_38 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_1615) begin
          tgtPages_39 <= GEN_3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1640) begin
          if(T_1635) begin
            pages_0 <= T_1255;
          end else begin
            pages_0 <= T_964;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1647) begin
          if(T_1635) begin
            pages_1 <= T_964;
          end else begin
            pages_1 <= T_1255;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1641) begin
          if(T_1635) begin
            pages_2 <= T_1255;
          end else begin
            pages_2 <= T_964;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1648) begin
          if(T_1635) begin
            pages_3 <= T_964;
          end else begin
            pages_3 <= T_1255;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1642) begin
          if(T_1635) begin
            pages_4 <= T_1255;
          end else begin
            pages_4 <= T_964;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(T_1649) begin
          if(T_1635) begin
            pages_5 <= T_964;
          end else begin
            pages_5 <= T_1255;
          end
        end
      end
    end
    if(reset) begin
      pageValid <= 6'h0;
    end else begin
      pageValid <= GEN_445[5:0];
    end
    if(reset) begin
      isValid <= 40'h0;
    end else begin
      isValid <= GEN_395[39:0];
    end
    if(1'h0) begin
    end else begin
      isReturn <= GEN_396[39:0];
    end
    if(1'h0) begin
    end else begin
      isJump <= GEN_397[39:0];
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h0 == T_1615) begin
          brIdx_0 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1 == T_1615) begin
          brIdx_1 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h2 == T_1615) begin
          brIdx_2 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h3 == T_1615) begin
          brIdx_3 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h4 == T_1615) begin
          brIdx_4 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h5 == T_1615) begin
          brIdx_5 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h6 == T_1615) begin
          brIdx_6 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h7 == T_1615) begin
          brIdx_7 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h8 == T_1615) begin
          brIdx_8 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h9 == T_1615) begin
          brIdx_9 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'ha == T_1615) begin
          brIdx_10 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hb == T_1615) begin
          brIdx_11 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hc == T_1615) begin
          brIdx_12 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hd == T_1615) begin
          brIdx_13 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'he == T_1615) begin
          brIdx_14 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'hf == T_1615) begin
          brIdx_15 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h10 == T_1615) begin
          brIdx_16 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h11 == T_1615) begin
          brIdx_17 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h12 == T_1615) begin
          brIdx_18 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h13 == T_1615) begin
          brIdx_19 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h14 == T_1615) begin
          brIdx_20 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h15 == T_1615) begin
          brIdx_21 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h16 == T_1615) begin
          brIdx_22 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h17 == T_1615) begin
          brIdx_23 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h18 == T_1615) begin
          brIdx_24 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h19 == T_1615) begin
          brIdx_25 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1a == T_1615) begin
          brIdx_26 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1b == T_1615) begin
          brIdx_27 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1c == T_1615) begin
          brIdx_28 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1d == T_1615) begin
          brIdx_29 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1e == T_1615) begin
          brIdx_30 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h1f == T_1615) begin
          brIdx_31 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h20 == T_1615) begin
          brIdx_32 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h21 == T_1615) begin
          brIdx_33 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h22 == T_1615) begin
          brIdx_34 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h23 == T_1615) begin
          brIdx_35 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h24 == T_1615) begin
          brIdx_36 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h25 == T_1615) begin
          brIdx_37 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h26 == T_1615) begin
          brIdx_38 <= GEN_4;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(r_btb_update_valid) begin
        if(6'h27 == T_1615) begin
          brIdx_39 <= GEN_4;
        end
      end
    end
    if(reset) begin
      T_777 <= 1'h0;
    end else begin
      T_777 <= io_btb_update_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_valid <= io_btb_update_bits_prediction_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_taken <= io_btb_update_bits_prediction_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_mask <= io_btb_update_bits_prediction_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_bridx <= io_btb_update_bits_prediction_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_target <= io_btb_update_bits_prediction_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_entry <= io_btb_update_bits_prediction_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_bht_history <= io_btb_update_bits_prediction_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_prediction_bits_bht_value <= io_btb_update_bits_prediction_bits_bht_value;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_pc <= io_btb_update_bits_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_target <= io_btb_update_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_taken <= io_btb_update_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_isValid <= io_btb_update_bits_isValid;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_isJump <= io_btb_update_bits_isJump;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_isReturn <= io_btb_update_bits_isReturn;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_btb_update_valid) begin
        T_778_br_pc <= io_btb_update_bits_br_pc;
      end
    end
    if(reset) begin
      nextRepl <= 6'h0;
    end else begin
      if(T_1548) begin
        if(T_1551) begin
          nextRepl <= 6'h0;
        end else begin
          nextRepl <= T_1554;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1603) begin
        if(T_1611) begin
          nextPageRepl <= {{2'd0}, T_1612};
        end else begin
          nextPageRepl <= T_1609;
        end
      end
    end
    if(T_2209_T_2234_en & T_2209_T_2234_mask) begin
      T_2209[T_2209_T_2234_addr] <= T_2209_T_2234_data;
    end
    if(1'h0) begin
    end else begin
      if(T_2231) begin
        if(io_bht_update_bits_mispredict) begin
          T_2211 <= T_2245;
        end else begin
          if(T_2218) begin
            T_2211 <= T_2230;
          end
        end
      end else begin
        if(T_2218) begin
          T_2211 <= T_2230;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(T_2288) begin
          if(T_2269) begin
            T_2252 <= T_2295;
          end else begin
            if(io_ras_update_bits_isCall) begin
              if(T_2272) begin
                T_2252 <= T_2275;
              end
            end
          end
        end else begin
          if(io_ras_update_bits_isCall) begin
            if(T_2272) begin
              T_2252 <= T_2275;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(T_2288) begin
          if(T_2269) begin
            T_2254 <= T_2302;
          end else begin
            if(io_ras_update_bits_isCall) begin
              T_2254 <= T_2282;
            end
          end
        end else begin
          if(io_ras_update_bits_isCall) begin
            T_2254 <= T_2282;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(io_ras_update_bits_isCall) begin
          if(1'h0 == T_2282) begin
            T_2261_0 <= GEN_6;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ras_update_valid) begin
        if(io_ras_update_bits_isCall) begin
          if(T_2282) begin
            T_2261_1 <= GEN_6;
          end
        end
      end
    end
  end
endmodule
module Frontend(
  input   clk,
  input   reset,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input   io_cpu_req_bits_speculative,
  input   io_cpu_resp_ready,
  output  io_cpu_resp_valid,
  output  io_cpu_resp_bits_btb_valid,
  output  io_cpu_resp_bits_btb_bits_taken,
  output [1:0] io_cpu_resp_bits_btb_bits_mask,
  output  io_cpu_resp_bits_btb_bits_bridx,
  output [38:0] io_cpu_resp_bits_btb_bits_target,
  output [5:0] io_cpu_resp_bits_btb_bits_entry,
  output [6:0] io_cpu_resp_bits_btb_bits_bht_history,
  output [1:0] io_cpu_resp_bits_btb_bits_bht_value,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output [1:0] io_cpu_resp_bits_mask,
  output  io_cpu_resp_bits_xcpt_if,
  output  io_cpu_resp_bits_replay,
  input   io_cpu_btb_update_valid,
  input   io_cpu_btb_update_bits_prediction_valid,
  input   io_cpu_btb_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_mask,
  input   io_cpu_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_btb_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input  [38:0] io_cpu_btb_update_bits_target,
  input   io_cpu_btb_update_bits_taken,
  input   io_cpu_btb_update_bits_isValid,
  input   io_cpu_btb_update_bits_isJump,
  input   io_cpu_btb_update_bits_isReturn,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input   io_cpu_bht_update_valid,
  input   io_cpu_bht_update_bits_prediction_valid,
  input   io_cpu_bht_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_mask,
  input   io_cpu_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_bht_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input   io_cpu_bht_update_bits_taken,
  input   io_cpu_bht_update_bits_mispredict,
  input   io_cpu_ras_update_valid,
  input   io_cpu_ras_update_bits_isCall,
  input   io_cpu_ras_update_bits_isReturn,
  input  [38:0] io_cpu_ras_update_bits_returnAddr,
  input   io_cpu_ras_update_bits_prediction_valid,
  input   io_cpu_ras_update_bits_prediction_bits_taken,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_mask,
  input   io_cpu_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_ras_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
  input   io_cpu_flush_icache,
  input   io_cpu_flush_tlb,
  output [39:0] io_cpu_npc,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_req_valid;
  wire [38:0] icache_io_req_bits_addr;
  wire [19:0] icache_io_s1_ppn;
  wire  icache_io_s1_kill;
  wire  icache_io_s2_kill;
  wire  icache_io_resp_ready;
  wire  icache_io_resp_valid;
  wire [15:0] icache_io_resp_bits_data;
  wire [63:0] icache_io_resp_bits_datablock;
  wire  icache_io_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [10:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [27:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_pum;
  wire  tlb_io_ptw_req_bits_mxr;
  wire [26:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [15:0] tlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [37:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [3:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  reg [39:0] s1_pc_;
  reg [63:0] GEN_16;
  wire [39:0] T_1483;
  wire [39:0] T_1485;
  wire [39:0] s1_pc;
  reg  s1_speculative;
  reg [31:0] GEN_26;
  reg  s1_same_block;
  reg [31:0] GEN_28;
  reg  s2_valid;
  reg [31:0] GEN_29;
  reg [39:0] s2_pc;
  reg [63:0] GEN_30;
  reg  s2_btb_resp_valid;
  reg [31:0] GEN_31;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] GEN_32;
  reg [1:0] s2_btb_resp_bits_mask;
  reg [31:0] GEN_33;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] GEN_34;
  reg [38:0] s2_btb_resp_bits_target;
  reg [63:0] GEN_35;
  reg [5:0] s2_btb_resp_bits_entry;
  reg [31:0] GEN_36;
  reg [6:0] s2_btb_resp_bits_bht_history;
  reg [31:0] GEN_37;
  reg [1:0] s2_btb_resp_bits_bht_value;
  reg [31:0] GEN_38;
  reg  s2_xcpt_if;
  reg [31:0] GEN_39;
  reg  s2_speculative;
  reg [31:0] GEN_40;
  reg  s2_cacheable;
  reg [31:0] GEN_41;
  wire [39:0] T_1511;
  wire [39:0] T_1513;
  wire [39:0] T_1514;
  wire [40:0] T_1516;
  wire [39:0] ntpc;
  wire [39:0] T_1518;
  wire [39:0] T_1520;
  wire  ntpc_same_block;
  wire [39:0] predicted_npc;
  wire  predicted_taken;
  wire  T_1523;
  wire  icmiss;
  wire [39:0] npc;
  wire  T_1525;
  wire  T_1527;
  wire  T_1528;
  wire  T_1530;
  wire  T_1531;
  wire  s0_same_block;
  wire  T_1533;
  wire  stall;
  wire  T_1535;
  wire  T_1537;
  wire  T_1538;
  wire  T_1540;
  wire  T_1541;
  wire  T_1542;
  wire  T_1543;
  wire  T_1544;
  wire [39:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [39:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [39:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [39:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  BTB_1_clk;
  wire  BTB_1_reset;
  wire  BTB_1_io_req_valid;
  wire [38:0] BTB_1_io_req_bits_addr;
  wire  BTB_1_io_resp_valid;
  wire  BTB_1_io_resp_bits_taken;
  wire [1:0] BTB_1_io_resp_bits_mask;
  wire  BTB_1_io_resp_bits_bridx;
  wire [38:0] BTB_1_io_resp_bits_target;
  wire [5:0] BTB_1_io_resp_bits_entry;
  wire [6:0] BTB_1_io_resp_bits_bht_history;
  wire [1:0] BTB_1_io_resp_bits_bht_value;
  wire  BTB_1_io_btb_update_valid;
  wire  BTB_1_io_btb_update_bits_prediction_valid;
  wire  BTB_1_io_btb_update_bits_prediction_bits_taken;
  wire [1:0] BTB_1_io_btb_update_bits_prediction_bits_mask;
  wire  BTB_1_io_btb_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_btb_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_btb_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1_io_btb_update_bits_pc;
  wire [38:0] BTB_1_io_btb_update_bits_target;
  wire  BTB_1_io_btb_update_bits_taken;
  wire  BTB_1_io_btb_update_bits_isValid;
  wire  BTB_1_io_btb_update_bits_isJump;
  wire  BTB_1_io_btb_update_bits_isReturn;
  wire [38:0] BTB_1_io_btb_update_bits_br_pc;
  wire  BTB_1_io_bht_update_valid;
  wire  BTB_1_io_bht_update_bits_prediction_valid;
  wire  BTB_1_io_bht_update_bits_prediction_bits_taken;
  wire [1:0] BTB_1_io_bht_update_bits_prediction_bits_mask;
  wire  BTB_1_io_bht_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_bht_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_bht_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1_io_bht_update_bits_pc;
  wire  BTB_1_io_bht_update_bits_taken;
  wire  BTB_1_io_bht_update_bits_mispredict;
  wire  BTB_1_io_ras_update_valid;
  wire  BTB_1_io_ras_update_bits_isCall;
  wire  BTB_1_io_ras_update_bits_isReturn;
  wire [38:0] BTB_1_io_ras_update_bits_returnAddr;
  wire  BTB_1_io_ras_update_bits_prediction_valid;
  wire  BTB_1_io_ras_update_bits_prediction_bits_taken;
  wire [1:0] BTB_1_io_ras_update_bits_prediction_bits_mask;
  wire  BTB_1_io_ras_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1_io_ras_update_bits_prediction_bits_target;
  wire [5:0] BTB_1_io_ras_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1_io_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1_io_ras_update_bits_prediction_bits_bht_value;
  wire  T_1556;
  wire  GEN_17;
  wire  GEN_18;
  wire [1:0] GEN_19;
  wire  GEN_20;
  wire [38:0] GEN_21;
  wire [5:0] GEN_22;
  wire [6:0] GEN_23;
  wire [1:0] GEN_24;
  wire  T_1558;
  wire  T_1559;
  wire [39:0] T_1560;
  wire [39:0] GEN_25;
  wire [27:0] T_1567;
  wire  T_1574;
  wire  T_1575;
  wire  T_1576;
  wire  T_1577;
  wire  T_1578;
  wire  T_1579;
  wire  T_1581;
  wire  T_1582;
  wire  T_1586;
  wire  T_1587;
  wire  T_1588;
  wire  T_1589;
  wire  T_1590;
  wire [39:0] T_1591;
  wire  T_1592;
  wire [5:0] GEN_27;
  wire [5:0] T_1593;
  wire [63:0] T_1594;
  wire  T_1596;
  wire [2:0] T_1597;
  wire  T_1600;
  wire  T_1602;
  wire  T_1603;
  ICache icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_ppn(icache_io_s1_ppn),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_ready(icache_io_resp_ready),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_datablock(icache_io_resp_bits_datablock),
    .io_invalidate(icache_io_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(tlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(tlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(tlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  BTB BTB_1 (
    .clk(BTB_1_clk),
    .reset(BTB_1_reset),
    .io_req_valid(BTB_1_io_req_valid),
    .io_req_bits_addr(BTB_1_io_req_bits_addr),
    .io_resp_valid(BTB_1_io_resp_valid),
    .io_resp_bits_taken(BTB_1_io_resp_bits_taken),
    .io_resp_bits_mask(BTB_1_io_resp_bits_mask),
    .io_resp_bits_bridx(BTB_1_io_resp_bits_bridx),
    .io_resp_bits_target(BTB_1_io_resp_bits_target),
    .io_resp_bits_entry(BTB_1_io_resp_bits_entry),
    .io_resp_bits_bht_history(BTB_1_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(BTB_1_io_resp_bits_bht_value),
    .io_btb_update_valid(BTB_1_io_btb_update_valid),
    .io_btb_update_bits_prediction_valid(BTB_1_io_btb_update_bits_prediction_valid),
    .io_btb_update_bits_prediction_bits_taken(BTB_1_io_btb_update_bits_prediction_bits_taken),
    .io_btb_update_bits_prediction_bits_mask(BTB_1_io_btb_update_bits_prediction_bits_mask),
    .io_btb_update_bits_prediction_bits_bridx(BTB_1_io_btb_update_bits_prediction_bits_bridx),
    .io_btb_update_bits_prediction_bits_target(BTB_1_io_btb_update_bits_prediction_bits_target),
    .io_btb_update_bits_prediction_bits_entry(BTB_1_io_btb_update_bits_prediction_bits_entry),
    .io_btb_update_bits_prediction_bits_bht_history(BTB_1_io_btb_update_bits_prediction_bits_bht_history),
    .io_btb_update_bits_prediction_bits_bht_value(BTB_1_io_btb_update_bits_prediction_bits_bht_value),
    .io_btb_update_bits_pc(BTB_1_io_btb_update_bits_pc),
    .io_btb_update_bits_target(BTB_1_io_btb_update_bits_target),
    .io_btb_update_bits_taken(BTB_1_io_btb_update_bits_taken),
    .io_btb_update_bits_isValid(BTB_1_io_btb_update_bits_isValid),
    .io_btb_update_bits_isJump(BTB_1_io_btb_update_bits_isJump),
    .io_btb_update_bits_isReturn(BTB_1_io_btb_update_bits_isReturn),
    .io_btb_update_bits_br_pc(BTB_1_io_btb_update_bits_br_pc),
    .io_bht_update_valid(BTB_1_io_bht_update_valid),
    .io_bht_update_bits_prediction_valid(BTB_1_io_bht_update_bits_prediction_valid),
    .io_bht_update_bits_prediction_bits_taken(BTB_1_io_bht_update_bits_prediction_bits_taken),
    .io_bht_update_bits_prediction_bits_mask(BTB_1_io_bht_update_bits_prediction_bits_mask),
    .io_bht_update_bits_prediction_bits_bridx(BTB_1_io_bht_update_bits_prediction_bits_bridx),
    .io_bht_update_bits_prediction_bits_target(BTB_1_io_bht_update_bits_prediction_bits_target),
    .io_bht_update_bits_prediction_bits_entry(BTB_1_io_bht_update_bits_prediction_bits_entry),
    .io_bht_update_bits_prediction_bits_bht_history(BTB_1_io_bht_update_bits_prediction_bits_bht_history),
    .io_bht_update_bits_prediction_bits_bht_value(BTB_1_io_bht_update_bits_prediction_bits_bht_value),
    .io_bht_update_bits_pc(BTB_1_io_bht_update_bits_pc),
    .io_bht_update_bits_taken(BTB_1_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(BTB_1_io_bht_update_bits_mispredict),
    .io_ras_update_valid(BTB_1_io_ras_update_valid),
    .io_ras_update_bits_isCall(BTB_1_io_ras_update_bits_isCall),
    .io_ras_update_bits_isReturn(BTB_1_io_ras_update_bits_isReturn),
    .io_ras_update_bits_returnAddr(BTB_1_io_ras_update_bits_returnAddr),
    .io_ras_update_bits_prediction_valid(BTB_1_io_ras_update_bits_prediction_valid),
    .io_ras_update_bits_prediction_bits_taken(BTB_1_io_ras_update_bits_prediction_bits_taken),
    .io_ras_update_bits_prediction_bits_mask(BTB_1_io_ras_update_bits_prediction_bits_mask),
    .io_ras_update_bits_prediction_bits_bridx(BTB_1_io_ras_update_bits_prediction_bits_bridx),
    .io_ras_update_bits_prediction_bits_target(BTB_1_io_ras_update_bits_prediction_bits_target),
    .io_ras_update_bits_prediction_bits_entry(BTB_1_io_ras_update_bits_prediction_bits_entry),
    .io_ras_update_bits_prediction_bits_bht_history(BTB_1_io_ras_update_bits_prediction_bits_bht_history),
    .io_ras_update_bits_prediction_bits_bht_value(BTB_1_io_ras_update_bits_prediction_bits_bht_value)
  );
  assign io_cpu_resp_valid = T_1590;
  assign io_cpu_resp_bits_btb_valid = s2_btb_resp_valid;
  assign io_cpu_resp_bits_btb_bits_taken = s2_btb_resp_bits_taken;
  assign io_cpu_resp_bits_btb_bits_mask = s2_btb_resp_bits_mask;
  assign io_cpu_resp_bits_btb_bits_bridx = s2_btb_resp_bits_bridx;
  assign io_cpu_resp_bits_btb_bits_target = s2_btb_resp_bits_target;
  assign io_cpu_resp_bits_btb_bits_entry = s2_btb_resp_bits_entry;
  assign io_cpu_resp_bits_btb_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign io_cpu_resp_bits_btb_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_bits_data = T_1594[31:0];
  assign io_cpu_resp_bits_mask = T_1597[1:0];
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign io_cpu_resp_bits_replay = T_1603;
  assign io_cpu_npc = T_1591;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = tlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = tlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_req_valid = T_1575;
  assign icache_io_req_bits_addr = io_cpu_npc[38:0];
  assign icache_io_s1_ppn = tlb_io_resp_ppn;
  assign icache_io_s1_kill = T_1579;
  assign icache_io_s2_kill = T_1582;
  assign icache_io_resp_ready = T_1587;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_mem_acquire_ready = io_mem_acquire_ready;
  assign icache_io_mem_grant_valid = io_mem_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_1556;
  assign tlb_io_req_bits_vpn = T_1567;
  assign tlb_io_req_bits_passthrough = 1'h0;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_store = 1'h0;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_1483 = ~ s1_pc_;
  assign T_1485 = T_1483 | 40'h1;
  assign s1_pc = ~ T_1485;
  assign T_1511 = ~ s1_pc;
  assign T_1513 = T_1511 | 40'h3;
  assign T_1514 = ~ T_1513;
  assign T_1516 = T_1514 + 40'h4;
  assign ntpc = T_1516[39:0];
  assign T_1518 = ntpc & 40'h8;
  assign T_1520 = s1_pc & 40'h8;
  assign ntpc_same_block = T_1518 == T_1520;
  assign predicted_npc = GEN_25;
  assign predicted_taken = T_1558;
  assign T_1523 = icache_io_resp_valid == 1'h0;
  assign icmiss = s2_valid & T_1523;
  assign npc = icmiss ? s2_pc : predicted_npc;
  assign T_1525 = predicted_taken == 1'h0;
  assign T_1527 = icmiss == 1'h0;
  assign T_1528 = T_1525 & T_1527;
  assign T_1530 = io_cpu_req_valid == 1'h0;
  assign T_1531 = T_1528 & T_1530;
  assign s0_same_block = T_1531 & ntpc_same_block;
  assign T_1533 = io_cpu_resp_ready == 1'h0;
  assign stall = io_cpu_resp_valid & T_1533;
  assign T_1535 = stall == 1'h0;
  assign T_1537 = tlb_io_resp_miss == 1'h0;
  assign T_1538 = s0_same_block & T_1537;
  assign T_1540 = s2_speculative == 1'h0;
  assign T_1541 = s2_valid & T_1540;
  assign T_1542 = s1_speculative | T_1541;
  assign T_1543 = T_1542 | predicted_taken;
  assign T_1544 = icmiss ? s2_speculative : T_1543;
  assign GEN_0 = T_1527 ? s1_pc : s2_pc;
  assign GEN_1 = T_1527 ? s1_speculative : s2_speculative;
  assign GEN_2 = T_1527 ? tlb_io_resp_cacheable : s2_cacheable;
  assign GEN_3 = T_1527 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign GEN_4 = T_1535 ? T_1538 : s1_same_block;
  assign GEN_5 = T_1535 ? io_cpu_npc : s1_pc_;
  assign GEN_6 = T_1535 ? T_1544 : s1_speculative;
  assign GEN_7 = T_1535 ? T_1527 : s2_valid;
  assign GEN_8 = T_1535 ? GEN_0 : s2_pc;
  assign GEN_9 = T_1535 ? GEN_1 : s2_speculative;
  assign GEN_10 = T_1535 ? GEN_2 : s2_cacheable;
  assign GEN_11 = T_1535 ? GEN_3 : s2_xcpt_if;
  assign GEN_12 = io_cpu_req_valid ? 1'h0 : GEN_4;
  assign GEN_13 = io_cpu_req_valid ? io_cpu_npc : GEN_5;
  assign GEN_14 = io_cpu_req_valid ? io_cpu_req_bits_speculative : GEN_6;
  assign GEN_15 = io_cpu_req_valid ? 1'h0 : GEN_7;
  assign BTB_1_clk = clk;
  assign BTB_1_reset = reset;
  assign BTB_1_io_req_valid = T_1556;
  assign BTB_1_io_req_bits_addr = s1_pc_[38:0];
  assign BTB_1_io_btb_update_valid = io_cpu_btb_update_valid;
  assign BTB_1_io_btb_update_bits_prediction_valid = io_cpu_btb_update_bits_prediction_valid;
  assign BTB_1_io_btb_update_bits_prediction_bits_taken = io_cpu_btb_update_bits_prediction_bits_taken;
  assign BTB_1_io_btb_update_bits_prediction_bits_mask = io_cpu_btb_update_bits_prediction_bits_mask;
  assign BTB_1_io_btb_update_bits_prediction_bits_bridx = io_cpu_btb_update_bits_prediction_bits_bridx;
  assign BTB_1_io_btb_update_bits_prediction_bits_target = io_cpu_btb_update_bits_prediction_bits_target;
  assign BTB_1_io_btb_update_bits_prediction_bits_entry = io_cpu_btb_update_bits_prediction_bits_entry;
  assign BTB_1_io_btb_update_bits_prediction_bits_bht_history = io_cpu_btb_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_btb_update_bits_prediction_bits_bht_value = io_cpu_btb_update_bits_prediction_bits_bht_value;
  assign BTB_1_io_btb_update_bits_pc = io_cpu_btb_update_bits_pc;
  assign BTB_1_io_btb_update_bits_target = io_cpu_btb_update_bits_target;
  assign BTB_1_io_btb_update_bits_taken = io_cpu_btb_update_bits_taken;
  assign BTB_1_io_btb_update_bits_isValid = io_cpu_btb_update_bits_isValid;
  assign BTB_1_io_btb_update_bits_isJump = io_cpu_btb_update_bits_isJump;
  assign BTB_1_io_btb_update_bits_isReturn = io_cpu_btb_update_bits_isReturn;
  assign BTB_1_io_btb_update_bits_br_pc = io_cpu_btb_update_bits_br_pc;
  assign BTB_1_io_bht_update_valid = io_cpu_bht_update_valid;
  assign BTB_1_io_bht_update_bits_prediction_valid = io_cpu_bht_update_bits_prediction_valid;
  assign BTB_1_io_bht_update_bits_prediction_bits_taken = io_cpu_bht_update_bits_prediction_bits_taken;
  assign BTB_1_io_bht_update_bits_prediction_bits_mask = io_cpu_bht_update_bits_prediction_bits_mask;
  assign BTB_1_io_bht_update_bits_prediction_bits_bridx = io_cpu_bht_update_bits_prediction_bits_bridx;
  assign BTB_1_io_bht_update_bits_prediction_bits_target = io_cpu_bht_update_bits_prediction_bits_target;
  assign BTB_1_io_bht_update_bits_prediction_bits_entry = io_cpu_bht_update_bits_prediction_bits_entry;
  assign BTB_1_io_bht_update_bits_prediction_bits_bht_history = io_cpu_bht_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_bht_update_bits_prediction_bits_bht_value = io_cpu_bht_update_bits_prediction_bits_bht_value;
  assign BTB_1_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc;
  assign BTB_1_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken;
  assign BTB_1_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict;
  assign BTB_1_io_ras_update_valid = io_cpu_ras_update_valid;
  assign BTB_1_io_ras_update_bits_isCall = io_cpu_ras_update_bits_isCall;
  assign BTB_1_io_ras_update_bits_isReturn = io_cpu_ras_update_bits_isReturn;
  assign BTB_1_io_ras_update_bits_returnAddr = io_cpu_ras_update_bits_returnAddr;
  assign BTB_1_io_ras_update_bits_prediction_valid = io_cpu_ras_update_bits_prediction_valid;
  assign BTB_1_io_ras_update_bits_prediction_bits_taken = io_cpu_ras_update_bits_prediction_bits_taken;
  assign BTB_1_io_ras_update_bits_prediction_bits_mask = io_cpu_ras_update_bits_prediction_bits_mask;
  assign BTB_1_io_ras_update_bits_prediction_bits_bridx = io_cpu_ras_update_bits_prediction_bits_bridx;
  assign BTB_1_io_ras_update_bits_prediction_bits_target = io_cpu_ras_update_bits_prediction_bits_target;
  assign BTB_1_io_ras_update_bits_prediction_bits_entry = io_cpu_ras_update_bits_prediction_bits_entry;
  assign BTB_1_io_ras_update_bits_prediction_bits_bht_history = io_cpu_ras_update_bits_prediction_bits_bht_history;
  assign BTB_1_io_ras_update_bits_prediction_bits_bht_value = io_cpu_ras_update_bits_prediction_bits_bht_value;
  assign T_1556 = T_1535 & T_1527;
  assign GEN_17 = T_1556 ? BTB_1_io_resp_valid : s2_btb_resp_valid;
  assign GEN_18 = T_1556 ? BTB_1_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign GEN_19 = T_1556 ? BTB_1_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign GEN_20 = T_1556 ? BTB_1_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign GEN_21 = T_1556 ? BTB_1_io_resp_bits_target : s2_btb_resp_bits_target;
  assign GEN_22 = T_1556 ? BTB_1_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign GEN_23 = T_1556 ? BTB_1_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign GEN_24 = T_1556 ? BTB_1_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T_1558 = BTB_1_io_resp_valid & BTB_1_io_resp_bits_taken;
  assign T_1559 = BTB_1_io_resp_bits_target[38];
  assign T_1560 = {T_1559,BTB_1_io_resp_bits_target};
  assign GEN_25 = T_1558 ? T_1560 : ntpc;
  assign T_1567 = s1_pc[39:12];
  assign T_1574 = s0_same_block == 1'h0;
  assign T_1575 = T_1535 & T_1574;
  assign T_1576 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T_1577 = T_1576 | tlb_io_resp_xcpt_if;
  assign T_1578 = T_1577 | icmiss;
  assign T_1579 = T_1578 | io_cpu_flush_tlb;
  assign T_1581 = s2_cacheable == 1'h0;
  assign T_1582 = s2_speculative & T_1581;
  assign T_1586 = s1_same_block == 1'h0;
  assign T_1587 = T_1535 & T_1586;
  assign T_1588 = icache_io_resp_valid | icache_io_s2_kill;
  assign T_1589 = T_1588 | s2_xcpt_if;
  assign T_1590 = s2_valid & T_1589;
  assign T_1591 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T_1592 = s2_pc[2];
  assign GEN_27 = {{5'd0}, T_1592};
  assign T_1593 = GEN_27 << 5;
  assign T_1594 = icache_io_resp_bits_datablock >> T_1593;
  assign T_1596 = s2_pc[1];
  assign T_1597 = 3'h3 << T_1596;
  assign T_1600 = icache_io_s2_kill & T_1523;
  assign T_1602 = s2_xcpt_if == 1'h0;
  assign T_1603 = T_1600 & T_1602;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {2{$random}};
  s1_pc_ = GEN_16[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  s1_speculative = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  s1_same_block = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  s2_valid = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {2{$random}};
  s2_pc = GEN_30[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  s2_btb_resp_valid = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  s2_btb_resp_bits_taken = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  s2_btb_resp_bits_mask = GEN_33[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  s2_btb_resp_bits_bridx = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {2{$random}};
  s2_btb_resp_bits_target = GEN_35[38:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  s2_btb_resp_bits_entry = GEN_36[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  s2_btb_resp_bits_bht_history = GEN_37[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  s2_btb_resp_bits_bht_value = GEN_38[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  s2_xcpt_if = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  s2_speculative = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  s2_cacheable = GEN_41[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_pc_ <= io_cpu_npc;
      end else begin
        if(T_1535) begin
          s1_pc_ <= io_cpu_npc;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_speculative <= io_cpu_req_bits_speculative;
      end else begin
        if(T_1535) begin
          if(icmiss) begin
            s1_speculative <= s2_speculative;
          end else begin
            s1_speculative <= T_1543;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_same_block <= 1'h0;
      end else begin
        if(T_1535) begin
          s1_same_block <= T_1538;
        end
      end
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else begin
      if(io_cpu_req_valid) begin
        s2_valid <= 1'h0;
      end else begin
        if(T_1535) begin
          s2_valid <= T_1527;
        end
      end
    end
    if(reset) begin
      s2_pc <= 40'h1000;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_pc <= s1_pc;
        end
      end
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else begin
      if(T_1556) begin
        s2_btb_resp_valid <= BTB_1_io_resp_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_taken <= BTB_1_io_resp_bits_taken;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_mask <= BTB_1_io_resp_bits_mask;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_bridx <= BTB_1_io_resp_bits_bridx;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_target <= BTB_1_io_resp_bits_target;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_entry <= BTB_1_io_resp_bits_entry;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_bht_history <= BTB_1_io_resp_bits_bht_history;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1556) begin
        s2_btb_resp_bits_bht_value <= BTB_1_io_resp_bits_bht_value;
      end
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_xcpt_if <= tlb_io_resp_xcpt_if;
        end
      end
    end
    if(reset) begin
      s2_speculative <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_speculative <= s1_speculative;
        end
      end
    end
    if(reset) begin
      s2_cacheable <= 1'h0;
    end else begin
      if(T_1535) begin
        if(T_1527) begin
          s2_cacheable <= tlb_io_resp_cacheable;
        end
      end
    end
  end
endmodule
module WritebackUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [2:0] io_req_bits_addr_beat,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_req_bits_voluntary,
  input  [2:0] io_req_bits_r_type,
  input  [63:0] io_req_bits_data,
  input  [3:0] io_req_bits_way_en,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_data_req_ready,
  output  io_data_req_valid,
  output [3:0] io_data_req_bits_way_en,
  output [11:0] io_data_req_bits_addr,
  input  [63:0] io_data_resp,
  input   io_release_ready,
  output  io_release_valid,
  output [2:0] io_release_bits_addr_beat,
  output [25:0] io_release_bits_addr_block,
  output [1:0] io_release_bits_client_xact_id,
  output  io_release_bits_voluntary,
  output [2:0] io_release_bits_r_type,
  output [63:0] io_release_bits_data
);
  reg  active;
  reg [31:0] GEN_6;
  reg  r1_data_req_fired;
  reg [31:0] GEN_7;
  reg  r2_data_req_fired;
  reg [31:0] GEN_8;
  reg [3:0] data_req_cnt;
  reg [31:0] GEN_10;
  wire  T_664;
  reg [2:0] beat_cnt;
  reg [31:0] GEN_31;
  wire [3:0] T_669;
  wire [2:0] T_670;
  wire [2:0] GEN_0;
  reg [2:0] req_addr_beat;
  reg [31:0] GEN_32;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_33;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_34;
  reg  req_voluntary;
  reg [31:0] GEN_35;
  reg [2:0] req_r_type;
  reg [31:0] GEN_36;
  reg [63:0] req_data;
  reg [63:0] GEN_37;
  reg [3:0] req_way_en;
  reg [31:0] GEN_38;
  wire  T_768;
  wire  T_769;
  wire  T_770;
  wire [4:0] T_773;
  wire [3:0] T_774;
  wire [3:0] GEN_2;
  wire  T_776;
  wire [1:0] T_783;
  wire [3:0] GEN_29;
  wire [4:0] T_784;
  wire [3:0] T_785;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire  T_789;
  wire  T_791;
  wire  T_794;
  wire  GEN_9;
  wire  GEN_11;
  wire  GEN_12;
  wire [3:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [3:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  T_795;
  wire  GEN_20;
  wire [3:0] GEN_21;
  wire [2:0] GEN_22;
  wire [25:0] GEN_23;
  wire [1:0] GEN_24;
  wire  GEN_25;
  wire [2:0] GEN_26;
  wire [63:0] GEN_27;
  wire [3:0] GEN_28;
  wire  T_799;
  wire [5:0] req_idx;
  wire  fire;
  wire [19:0] T_802;
  wire [2:0] T_803;
  wire [8:0] T_804;
  wire [11:0] GEN_30;
  wire [11:0] T_805;
  wire [3:0] GEN_1;
  reg [31:0] GEN_39;
  assign io_req_ready = T_799;
  assign io_meta_read_valid = fire;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_1;
  assign io_meta_read_bits_tag = T_802;
  assign io_data_req_valid = fire;
  assign io_data_req_bits_way_en = req_way_en;
  assign io_data_req_bits_addr = T_805;
  assign io_release_valid = GEN_18;
  assign io_release_bits_addr_beat = beat_cnt;
  assign io_release_bits_addr_block = req_addr_block;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign io_release_bits_voluntary = req_voluntary;
  assign io_release_bits_r_type = req_r_type;
  assign io_release_bits_data = io_data_resp;
  assign T_664 = io_release_ready & io_release_valid;
  assign T_669 = beat_cnt + 3'h1;
  assign T_670 = T_669[2:0];
  assign GEN_0 = T_664 ? T_670 : beat_cnt;
  assign T_768 = io_data_req_ready & io_data_req_valid;
  assign T_769 = io_meta_read_ready & io_meta_read_valid;
  assign T_770 = T_768 & T_769;
  assign T_773 = data_req_cnt + 4'h1;
  assign T_774 = T_773[3:0];
  assign GEN_2 = T_770 ? T_774 : data_req_cnt;
  assign T_776 = io_release_ready == 1'h0;
  assign T_783 = r1_data_req_fired ? 2'h2 : 2'h1;
  assign GEN_29 = {{2'd0}, T_783};
  assign T_784 = data_req_cnt - GEN_29;
  assign T_785 = T_784[3:0];
  assign GEN_3 = T_776 ? 1'h0 : T_770;
  assign GEN_4 = T_776 ? 1'h0 : r1_data_req_fired;
  assign GEN_5 = T_776 ? T_785 : GEN_2;
  assign T_789 = r1_data_req_fired == 1'h0;
  assign T_791 = data_req_cnt < 4'h8;
  assign T_794 = T_791 | T_776;
  assign GEN_9 = T_789 ? T_794 : active;
  assign GEN_11 = r2_data_req_fired ? GEN_3 : T_770;
  assign GEN_12 = r2_data_req_fired ? GEN_4 : r1_data_req_fired;
  assign GEN_13 = r2_data_req_fired ? GEN_5 : GEN_2;
  assign GEN_14 = r2_data_req_fired ? GEN_9 : active;
  assign GEN_15 = active ? GEN_11 : r1_data_req_fired;
  assign GEN_16 = active ? GEN_12 : r2_data_req_fired;
  assign GEN_17 = active ? GEN_13 : data_req_cnt;
  assign GEN_18 = active ? r2_data_req_fired : 1'h0;
  assign GEN_19 = active ? GEN_14 : active;
  assign T_795 = io_req_ready & io_req_valid;
  assign GEN_20 = T_795 ? 1'h1 : GEN_19;
  assign GEN_21 = T_795 ? 4'h0 : GEN_17;
  assign GEN_22 = T_795 ? io_req_bits_addr_beat : req_addr_beat;
  assign GEN_23 = T_795 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_24 = T_795 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign GEN_25 = T_795 ? io_req_bits_voluntary : req_voluntary;
  assign GEN_26 = T_795 ? io_req_bits_r_type : req_r_type;
  assign GEN_27 = T_795 ? io_req_bits_data : req_data;
  assign GEN_28 = T_795 ? io_req_bits_way_en : req_way_en;
  assign T_799 = active == 1'h0;
  assign req_idx = req_addr_block[5:0];
  assign fire = active & T_791;
  assign T_802 = req_addr_block[25:6];
  assign T_803 = data_req_cnt[2:0];
  assign T_804 = {req_idx,T_803};
  assign GEN_30 = {{3'd0}, T_804};
  assign T_805 = GEN_30 << 3;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_39[3:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  active = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  r1_data_req_fired = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  r2_data_req_fired = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  data_req_cnt = GEN_10[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  beat_cnt = GEN_31[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  req_addr_beat = GEN_32[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  req_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  req_client_xact_id = GEN_34[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  req_voluntary = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  req_r_type = GEN_36[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {2{$random}};
  req_data = GEN_37[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  req_way_en = GEN_38[3:0];
  `endif
  GEN_39 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else begin
      if(T_795) begin
        active <= 1'h1;
      end else begin
        if(active) begin
          if(r2_data_req_fired) begin
            if(T_789) begin
              active <= T_794;
            end
          end
        end
      end
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else begin
      if(active) begin
        if(r2_data_req_fired) begin
          if(T_776) begin
            r1_data_req_fired <= 1'h0;
          end else begin
            r1_data_req_fired <= T_770;
          end
        end else begin
          r1_data_req_fired <= T_770;
        end
      end
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else begin
      if(active) begin
        if(r2_data_req_fired) begin
          if(T_776) begin
            r2_data_req_fired <= 1'h0;
          end else begin
            r2_data_req_fired <= r1_data_req_fired;
          end
        end else begin
          r2_data_req_fired <= r1_data_req_fired;
        end
      end
    end
    if(reset) begin
      data_req_cnt <= 4'h0;
    end else begin
      if(T_795) begin
        data_req_cnt <= 4'h0;
      end else begin
        if(active) begin
          if(r2_data_req_fired) begin
            if(T_776) begin
              data_req_cnt <= T_785;
            end else begin
              if(T_770) begin
                data_req_cnt <= T_774;
              end
            end
          end else begin
            if(T_770) begin
              data_req_cnt <= T_774;
            end
          end
        end
      end
    end
    if(reset) begin
      beat_cnt <= 3'h0;
    end else begin
      if(T_664) begin
        beat_cnt <= T_670;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_addr_beat <= io_req_bits_addr_beat;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_addr_block <= io_req_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_client_xact_id <= io_req_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_voluntary <= io_req_bits_voluntary;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_r_type <= io_req_bits_r_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_data <= io_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_795) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
  end
endmodule
module ProbeUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_p_type,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_rep_ready,
  output  io_rep_valid,
  output [2:0] io_rep_bits_addr_beat,
  output [25:0] io_rep_bits_addr_block,
  output [1:0] io_rep_bits_client_xact_id,
  output  io_rep_bits_voluntary,
  output [2:0] io_rep_bits_r_type,
  output [63:0] io_rep_bits_data,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  input  [3:0] io_way_en,
  input   io_mshr_rdy,
  input  [1:0] io_block_state_state
);
  reg [3:0] state;
  reg [31:0] GEN_16;
  reg [1:0] old_coh_state;
  reg [31:0] GEN_17;
  reg [3:0] way_en;
  reg [31:0] GEN_18;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_19;
  reg [1:0] req_p_type;
  reg [31:0] GEN_20;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_21;
  wire  tag_matches;
  wire [1:0] miss_coh_state;
  wire [1:0] reply_coh_state;
  wire  T_1107;
  wire [2:0] T_1108;
  wire  T_1137;
  wire [2:0] T_1138;
  wire  T_1139;
  wire [2:0] T_1140;
  wire  T_1141;
  wire [2:0] T_1142;
  wire [2:0] reply_addr_beat;
  wire [25:0] reply_addr_block;
  wire [1:0] reply_client_xact_id;
  wire  reply_voluntary;
  wire [2:0] reply_r_type;
  wire [63:0] reply_data;
  wire  T_1197;
  wire  T_1198;
  wire  T_1200;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1204;
  wire  T_1205;
  wire  T_1207;
  wire  T_1208;
  wire  T_1209;
  wire  T_1211;
  wire  T_1212;
  wire [19:0] T_1213;
  wire  T_1214;
  wire [1:0] T_1217;
  wire [1:0] T_1219;
  wire [1:0] T_1221;
  wire [1:0] T_1244_state;
  wire  T_1266;
  wire  T_1267;
  wire [3:0] GEN_0;
  wire [25:0] GEN_1;
  wire [1:0] GEN_2;
  wire [1:0] GEN_3;
  wire  T_1268;
  wire [3:0] GEN_4;
  wire  T_1269;
  wire [3:0] GEN_5;
  wire  T_1270;
  wire  T_1272;
  wire [3:0] GEN_6;
  wire [3:0] GEN_7;
  wire [1:0] GEN_8;
  wire [3:0] GEN_9;
  wire  T_1273;
  wire  T_1274;
  wire  T_1275;
  wire [3:0] T_1276;
  wire [3:0] GEN_10;
  wire  T_1278;
  wire [3:0] T_1279;
  wire [3:0] GEN_11;
  wire  T_1280;
  wire [3:0] GEN_12;
  wire  T_1281;
  wire  T_1282;
  wire [3:0] GEN_13;
  wire  T_1283;
  wire [3:0] GEN_14;
  wire [3:0] GEN_15;
  reg [31:0] GEN_22;
  assign io_req_ready = T_1197;
  assign io_rep_valid = T_1198;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_data = reply_data;
  assign io_meta_read_valid = T_1212;
  assign io_meta_read_bits_idx = req_addr_block[5:0];
  assign io_meta_read_bits_way_en = GEN_15;
  assign io_meta_read_bits_tag = T_1213;
  assign io_meta_write_valid = T_1214;
  assign io_meta_write_bits_idx = req_addr_block[5:0];
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_data_tag = T_1213;
  assign io_meta_write_bits_data_coh_state = T_1244_state;
  assign io_wb_req_valid = T_1266;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign io_wb_req_bits_data = reply_data;
  assign io_wb_req_bits_way_en = way_en;
  assign tag_matches = way_en != 4'h0;
  assign miss_coh_state = 2'h0;
  assign reply_coh_state = tag_matches ? old_coh_state : miss_coh_state;
  assign T_1107 = reply_coh_state == 2'h2;
  assign T_1108 = T_1107 ? 3'h0 : 3'h3;
  assign T_1137 = 2'h2 == req_p_type;
  assign T_1138 = T_1137 ? T_1108 : 3'h3;
  assign T_1139 = 2'h1 == req_p_type;
  assign T_1140 = T_1139 ? T_1108 : T_1138;
  assign T_1141 = 2'h0 == req_p_type;
  assign T_1142 = T_1141 ? T_1108 : T_1140;
  assign reply_addr_beat = 3'h0;
  assign reply_addr_block = req_addr_block;
  assign reply_client_xact_id = 2'h0;
  assign reply_voluntary = 1'h0;
  assign reply_r_type = T_1142;
  assign reply_data = 64'h0;
  assign T_1197 = state == 4'h0;
  assign T_1198 = state == 4'h5;
  assign T_1200 = io_rep_valid == 1'h0;
  assign T_1201 = io_rep_bits_r_type == 3'h0;
  assign T_1202 = io_rep_bits_r_type == 3'h1;
  assign T_1203 = io_rep_bits_r_type == 3'h2;
  assign T_1204 = T_1201 | T_1202;
  assign T_1205 = T_1204 | T_1203;
  assign T_1207 = T_1205 == 1'h0;
  assign T_1208 = T_1200 | T_1207;
  assign T_1209 = T_1208 | reset;
  assign T_1211 = T_1209 == 1'h0;
  assign T_1212 = state == 4'h1;
  assign T_1213 = req_addr_block[25:6];
  assign T_1214 = state == 4'h8;
  assign T_1217 = T_1137 ? 2'h0 : old_coh_state;
  assign T_1219 = T_1139 ? 2'h0 : T_1217;
  assign T_1221 = T_1141 ? 2'h0 : T_1219;
  assign T_1244_state = T_1221;
  assign T_1266 = state == 4'h6;
  assign T_1267 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1267 ? 4'h1 : state;
  assign GEN_1 = T_1267 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_2 = T_1267 ? io_req_bits_p_type : req_p_type;
  assign GEN_3 = T_1267 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign T_1268 = io_meta_read_ready & io_meta_read_valid;
  assign GEN_4 = T_1268 ? 4'h2 : GEN_0;
  assign T_1269 = state == 4'h2;
  assign GEN_5 = T_1269 ? 4'h3 : GEN_4;
  assign T_1270 = state == 4'h3;
  assign T_1272 = io_mshr_rdy == 1'h0;
  assign GEN_6 = T_1272 ? 4'h1 : 4'h4;
  assign GEN_7 = T_1270 ? GEN_6 : GEN_5;
  assign GEN_8 = T_1270 ? io_block_state_state : old_coh_state;
  assign GEN_9 = T_1270 ? io_way_en : way_en;
  assign T_1273 = state == 4'h4;
  assign T_1274 = old_coh_state == 2'h2;
  assign T_1275 = tag_matches & T_1274;
  assign T_1276 = T_1275 ? 4'h6 : 4'h5;
  assign GEN_10 = T_1273 ? T_1276 : GEN_7;
  assign T_1278 = T_1198 & io_rep_ready;
  assign T_1279 = tag_matches ? 4'h8 : 4'h0;
  assign GEN_11 = T_1278 ? T_1279 : GEN_10;
  assign T_1280 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_12 = T_1280 ? 4'h7 : GEN_11;
  assign T_1281 = state == 4'h7;
  assign T_1282 = T_1281 & io_wb_req_ready;
  assign GEN_13 = T_1282 ? 4'h8 : GEN_12;
  assign T_1283 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_14 = T_1283 ? 4'h0 : GEN_13;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_22[3:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  state = GEN_16[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  old_coh_state = GEN_17[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  way_en = GEN_18[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {1{$random}};
  req_addr_block = GEN_19[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  req_p_type = GEN_20[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_21 = {1{$random}};
  req_client_xact_id = GEN_21[1:0];
  `endif
  GEN_22 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_1283) begin
        state <= 4'h0;
      end else begin
        if(T_1282) begin
          state <= 4'h8;
        end else begin
          if(T_1280) begin
            state <= 4'h7;
          end else begin
            if(T_1278) begin
              if(tag_matches) begin
                state <= 4'h8;
              end else begin
                state <= 4'h0;
              end
            end else begin
              if(T_1273) begin
                if(T_1275) begin
                  state <= 4'h6;
                end else begin
                  state <= 4'h5;
                end
              end else begin
                if(T_1270) begin
                  if(T_1272) begin
                    state <= 4'h1;
                  end else begin
                    state <= 4'h4;
                  end
                end else begin
                  if(T_1269) begin
                    state <= 4'h3;
                  end else begin
                    if(T_1268) begin
                      state <= 4'h2;
                    end else begin
                      if(T_1267) begin
                        state <= 4'h1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1270) begin
        old_coh_state <= io_block_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1270) begin
        way_en <= io_way_en;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1267) begin
        req_addr_block <= io_req_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1267) begin
        req_p_type <= io_req_bits_p_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1267) begin
        req_client_xact_id <= io_req_bits_client_xact_id;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1211) begin
          $fwrite(32'h80000002,"Assertion failed: ProbeUnit should not send releases with data\n    at nbdcache.scala:677 assert(!io.rep.valid || !io.rep.bits.hasData(),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Arbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_tag,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_tag,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_tag,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire  grant_1;
  wire  T_564;
  wire  T_566;
  wire  T_567;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_564;
  assign io_out_valid = T_567;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_tag = GEN_3;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_564 = grant_1 & io_out_ready;
  assign T_566 = grant_1 == 1'h0;
  assign T_567 = T_566 | io_in_1_valid;
endmodule
module Arbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_data_tag,
  input  [1:0] io_in_0_bits_data_coh_state,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_data_tag,
  input  [1:0] io_in_1_bits_data_coh_state,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_data_tag,
  output [1:0] io_out_bits_data_coh_state,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire [1:0] GEN_4;
  wire  grant_1;
  wire  T_2390;
  wire  T_2392;
  wire  T_2393;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2390;
  assign io_out_valid = T_2393;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_data_tag = GEN_3;
  assign io_out_bits_data_coh_state = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data_coh_state : io_in_1_bits_data_coh_state;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_2390 = grant_1 & io_out_ready;
  assign T_2392 = grant_1 == 1'h0;
  assign T_2393 = T_2392 | io_in_1_valid;
endmodule
module LockingArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [10:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [10:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [10:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [10:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_is_builtin_type;
  wire [2:0] GEN_0_bits_a_type;
  wire [10:0] GEN_0_bits_union;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_10;
  wire [1:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire [10:0] GEN_15;
  wire [63:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [25:0] GEN_19;
  wire [1:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [2:0] GEN_23;
  wire [10:0] GEN_24;
  wire [63:0] GEN_25;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_is_builtin_type;
  wire [2:0] GEN_1_bits_a_type;
  wire [10:0] GEN_1_bits_union;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_is_builtin_type;
  wire [2:0] GEN_2_bits_a_type;
  wire [10:0] GEN_2_bits_union;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_is_builtin_type;
  wire [2:0] GEN_3_bits_a_type;
  wire [10:0] GEN_3_bits_union;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [25:0] GEN_4_bits_addr_block;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_is_builtin_type;
  wire [2:0] GEN_4_bits_a_type;
  wire [10:0] GEN_4_bits_union;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [25:0] GEN_5_bits_addr_block;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_is_builtin_type;
  wire [2:0] GEN_5_bits_a_type;
  wire [10:0] GEN_5_bits_union;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [25:0] GEN_6_bits_addr_block;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_is_builtin_type;
  wire [2:0] GEN_6_bits_a_type;
  wire [10:0] GEN_6_bits_union;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [25:0] GEN_7_bits_addr_block;
  wire [1:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_is_builtin_type;
  wire [2:0] GEN_7_bits_a_type;
  wire [10:0] GEN_7_bits_union;
  wire [63:0] GEN_7_bits_data;
  reg [2:0] T_882;
  reg [31:0] GEN_0;
  reg [1:0] T_884;
  reg [31:0] GEN_1;
  wire  T_886;
  wire [2:0] T_895_0;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire  T_900;
  wire [3:0] T_904;
  wire [2:0] T_905;
  wire [1:0] GEN_152;
  wire [2:0] GEN_153;
  wire [1:0] GEN_154;
  wire  T_907;
  wire  T_909;
  wire  T_911;
  wire  T_913;
  wire  T_914;
  wire  T_915;
  wire  T_917;
  wire  T_918;
  wire  T_919;
  wire  T_921;
  wire  T_922;
  wire  T_923;
  wire [1:0] GEN_155;
  wire [1:0] GEN_156;
  assign io_in_0_ready = T_915;
  assign io_in_1_ready = T_919;
  assign io_in_2_ready = T_923;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_addr_beat = GEN_3_bits_addr_beat;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_a_type = GEN_5_bits_a_type;
  assign io_out_bits_union = GEN_6_bits_union;
  assign io_out_bits_data = GEN_7_bits_data;
  assign io_chosen = GEN_154;
  assign choice = GEN_156;
  assign GEN_0_ready = GEN_17;
  assign GEN_0_valid = GEN_18;
  assign GEN_0_bits_addr_block = GEN_19;
  assign GEN_0_bits_client_xact_id = GEN_20;
  assign GEN_0_bits_addr_beat = GEN_21;
  assign GEN_0_bits_is_builtin_type = GEN_22;
  assign GEN_0_bits_a_type = GEN_23;
  assign GEN_0_bits_union = GEN_24;
  assign GEN_0_bits_data = GEN_25;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_ready : GEN_8;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_12;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_13;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_a_type : GEN_14;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_union : GEN_15;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_16;
  assign GEN_1_ready = GEN_17;
  assign GEN_1_valid = GEN_18;
  assign GEN_1_bits_addr_block = GEN_19;
  assign GEN_1_bits_client_xact_id = GEN_20;
  assign GEN_1_bits_addr_beat = GEN_21;
  assign GEN_1_bits_is_builtin_type = GEN_22;
  assign GEN_1_bits_a_type = GEN_23;
  assign GEN_1_bits_union = GEN_24;
  assign GEN_1_bits_data = GEN_25;
  assign GEN_2_ready = GEN_17;
  assign GEN_2_valid = GEN_18;
  assign GEN_2_bits_addr_block = GEN_19;
  assign GEN_2_bits_client_xact_id = GEN_20;
  assign GEN_2_bits_addr_beat = GEN_21;
  assign GEN_2_bits_is_builtin_type = GEN_22;
  assign GEN_2_bits_a_type = GEN_23;
  assign GEN_2_bits_union = GEN_24;
  assign GEN_2_bits_data = GEN_25;
  assign GEN_3_ready = GEN_17;
  assign GEN_3_valid = GEN_18;
  assign GEN_3_bits_addr_block = GEN_19;
  assign GEN_3_bits_client_xact_id = GEN_20;
  assign GEN_3_bits_addr_beat = GEN_21;
  assign GEN_3_bits_is_builtin_type = GEN_22;
  assign GEN_3_bits_a_type = GEN_23;
  assign GEN_3_bits_union = GEN_24;
  assign GEN_3_bits_data = GEN_25;
  assign GEN_4_ready = GEN_17;
  assign GEN_4_valid = GEN_18;
  assign GEN_4_bits_addr_block = GEN_19;
  assign GEN_4_bits_client_xact_id = GEN_20;
  assign GEN_4_bits_addr_beat = GEN_21;
  assign GEN_4_bits_is_builtin_type = GEN_22;
  assign GEN_4_bits_a_type = GEN_23;
  assign GEN_4_bits_union = GEN_24;
  assign GEN_4_bits_data = GEN_25;
  assign GEN_5_ready = GEN_17;
  assign GEN_5_valid = GEN_18;
  assign GEN_5_bits_addr_block = GEN_19;
  assign GEN_5_bits_client_xact_id = GEN_20;
  assign GEN_5_bits_addr_beat = GEN_21;
  assign GEN_5_bits_is_builtin_type = GEN_22;
  assign GEN_5_bits_a_type = GEN_23;
  assign GEN_5_bits_union = GEN_24;
  assign GEN_5_bits_data = GEN_25;
  assign GEN_6_ready = GEN_17;
  assign GEN_6_valid = GEN_18;
  assign GEN_6_bits_addr_block = GEN_19;
  assign GEN_6_bits_client_xact_id = GEN_20;
  assign GEN_6_bits_addr_beat = GEN_21;
  assign GEN_6_bits_is_builtin_type = GEN_22;
  assign GEN_6_bits_a_type = GEN_23;
  assign GEN_6_bits_union = GEN_24;
  assign GEN_6_bits_data = GEN_25;
  assign GEN_7_ready = GEN_17;
  assign GEN_7_valid = GEN_18;
  assign GEN_7_bits_addr_block = GEN_19;
  assign GEN_7_bits_client_xact_id = GEN_20;
  assign GEN_7_bits_addr_beat = GEN_21;
  assign GEN_7_bits_is_builtin_type = GEN_22;
  assign GEN_7_bits_a_type = GEN_23;
  assign GEN_7_bits_union = GEN_24;
  assign GEN_7_bits_data = GEN_25;
  assign T_886 = T_882 != 3'h0;
  assign T_895_0 = 3'h3;
  assign T_897 = io_out_bits_a_type == T_895_0;
  assign T_898 = io_out_bits_is_builtin_type & T_897;
  assign T_899 = io_out_ready & io_out_valid;
  assign T_900 = T_899 & T_898;
  assign T_904 = T_882 + 3'h1;
  assign T_905 = T_904[2:0];
  assign GEN_152 = T_900 ? io_chosen : T_884;
  assign GEN_153 = T_900 ? T_905 : T_882;
  assign GEN_154 = T_886 ? T_884 : choice;
  assign T_907 = io_in_0_valid | io_in_1_valid;
  assign T_909 = io_in_0_valid == 1'h0;
  assign T_911 = T_907 == 1'h0;
  assign T_913 = T_884 == 2'h0;
  assign T_914 = T_886 ? T_913 : 1'h1;
  assign T_915 = T_914 & io_out_ready;
  assign T_917 = T_884 == 2'h1;
  assign T_918 = T_886 ? T_917 : T_909;
  assign T_919 = T_918 & io_out_ready;
  assign T_921 = T_884 == 2'h2;
  assign T_922 = T_886 ? T_921 : T_911;
  assign T_923 = T_922 & io_out_ready;
  assign GEN_155 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_156 = io_in_0_valid ? 2'h0 : GEN_155;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_882 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_884 = GEN_1[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_882 <= 3'h0;
    end else begin
      if(T_900) begin
        T_882 <= T_905;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_900) begin
        T_884 <= io_chosen;
      end
    end
  end
endmodule
module Arbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_manager_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_manager_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_manager_id,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [2:0] GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire  T_637;
  wire  grant_1;
  wire  grant_2;
  wire  T_641;
  wire  T_642;
  wire  T_644;
  wire  T_645;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_641;
  assign io_in_2_ready = T_642;
  assign io_out_valid = T_645;
  assign io_out_bits_manager_xact_id = GEN_4;
  assign io_out_bits_manager_id = GEN_5;
  assign io_chosen = GEN_3;
  assign GEN_0 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_manager_id : io_in_2_bits_manager_id;
  assign GEN_3 = io_in_0_valid ? 2'h0 : GEN_0;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_manager_xact_id : GEN_1;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_manager_id : GEN_2;
  assign T_637 = io_in_0_valid | io_in_1_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_637 == 1'h0;
  assign T_641 = grant_1 & io_out_ready;
  assign T_642 = grant_2 & io_out_ready;
  assign T_644 = grant_2 == 1'h0;
  assign T_645 = T_644 | io_in_2_valid;
endmodule
module Arbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input  [3:0] io_in_1_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [3:0] io_out_bits_way_en,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [25:0] GEN_2;
  wire [1:0] GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_5;
  wire [63:0] GEN_6;
  wire [3:0] GEN_7;
  wire  grant_1;
  wire  T_1092;
  wire  T_1094;
  wire  T_1095;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1092;
  assign io_out_valid = T_1095;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_way_en = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr_block : io_in_1_bits_addr_block;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_voluntary : io_in_1_bits_voluntary;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_r_type : io_in_1_bits_r_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_1092 = grant_1 & io_out_ready;
  assign T_1094 = grant_1 == 1'h0;
  assign T_1095 = T_1094 | io_in_1_valid;
endmodule
module Arbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [6:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input   io_in_0_bits_phys,
  input  [4:0] io_in_0_bits_sdq_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [39:0] io_in_1_bits_addr,
  input  [6:0] io_in_1_bits_tag,
  input  [4:0] io_in_1_bits_cmd,
  input  [2:0] io_in_1_bits_typ,
  input   io_in_1_bits_phys,
  input  [4:0] io_in_1_bits_sdq_id,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [6:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output  io_out_bits_phys,
  output [4:0] io_out_bits_sdq_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [39:0] GEN_1;
  wire [6:0] GEN_2;
  wire [4:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire [4:0] GEN_6;
  wire  grant_1;
  wire  T_1510;
  wire  T_1512;
  wire  T_1513;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1510;
  assign io_out_valid = T_1513;
  assign io_out_bits_addr = GEN_1;
  assign io_out_bits_tag = GEN_2;
  assign io_out_bits_cmd = GEN_3;
  assign io_out_bits_typ = GEN_4;
  assign io_out_bits_phys = GEN_5;
  assign io_out_bits_sdq_id = GEN_6;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_typ : io_in_1_bits_typ;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_phys : io_in_1_bits_phys;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_sdq_id : io_in_1_bits_sdq_id;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_1510 = grant_1 & io_out_ready;
  assign T_1512 = grant_1 == 1'h0;
  assign T_1513 = T_1512 | io_in_1_valid;
endmodule
module Arbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_in_1_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  wire  GEN_0;
  wire  GEN_1;
  wire  grant_1;
  wire  T_58;
  wire  T_60;
  wire  T_61;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_58;
  assign io_out_valid = T_61;
  assign io_out_bits = GEN_1;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits : io_in_1_bits;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_58 = grant_1 & io_out_ready;
  assign T_60 = grant_1 == 1'h0;
  assign T_61 = T_60 | io_in_1_valid;
endmodule
module Queue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [39:0] io_enq_bits_addr,
  input  [6:0] io_enq_bits_tag,
  input  [4:0] io_enq_bits_cmd,
  input  [2:0] io_enq_bits_typ,
  input   io_enq_bits_phys,
  input  [4:0] io_enq_bits_sdq_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [39:0] io_deq_bits_addr,
  output [6:0] io_deq_bits_tag,
  output [4:0] io_deq_bits_cmd,
  output [2:0] io_deq_bits_typ,
  output  io_deq_bits_phys,
  output [4:0] io_deq_bits_sdq_id,
  output [4:0] io_count
);
  reg [39:0] ram_addr [0:15];
  reg [63:0] GEN_0;
  wire [39:0] ram_addr_T_704_data;
  wire [3:0] ram_addr_T_704_addr;
  wire  ram_addr_T_704_en;
  wire [39:0] ram_addr_T_622_data;
  wire [3:0] ram_addr_T_622_addr;
  wire  ram_addr_T_622_mask;
  wire  ram_addr_T_622_en;
  reg [6:0] ram_tag [0:15];
  reg [31:0] GEN_1;
  wire [6:0] ram_tag_T_704_data;
  wire [3:0] ram_tag_T_704_addr;
  wire  ram_tag_T_704_en;
  wire [6:0] ram_tag_T_622_data;
  wire [3:0] ram_tag_T_622_addr;
  wire  ram_tag_T_622_mask;
  wire  ram_tag_T_622_en;
  reg [4:0] ram_cmd [0:15];
  reg [31:0] GEN_2;
  wire [4:0] ram_cmd_T_704_data;
  wire [3:0] ram_cmd_T_704_addr;
  wire  ram_cmd_T_704_en;
  wire [4:0] ram_cmd_T_622_data;
  wire [3:0] ram_cmd_T_622_addr;
  wire  ram_cmd_T_622_mask;
  wire  ram_cmd_T_622_en;
  reg [2:0] ram_typ [0:15];
  reg [31:0] GEN_3;
  wire [2:0] ram_typ_T_704_data;
  wire [3:0] ram_typ_T_704_addr;
  wire  ram_typ_T_704_en;
  wire [2:0] ram_typ_T_622_data;
  wire [3:0] ram_typ_T_622_addr;
  wire  ram_typ_T_622_mask;
  wire  ram_typ_T_622_en;
  reg  ram_phys [0:15];
  reg [31:0] GEN_4;
  wire  ram_phys_T_704_data;
  wire [3:0] ram_phys_T_704_addr;
  wire  ram_phys_T_704_en;
  wire  ram_phys_T_622_data;
  wire [3:0] ram_phys_T_622_addr;
  wire  ram_phys_T_622_mask;
  wire  ram_phys_T_622_en;
  reg [4:0] ram_sdq_id [0:15];
  reg [31:0] GEN_5;
  wire [4:0] ram_sdq_id_T_704_data;
  wire [3:0] ram_sdq_id_T_704_addr;
  wire  ram_sdq_id_T_704_en;
  wire [4:0] ram_sdq_id_T_622_data;
  wire [3:0] ram_sdq_id_T_622_addr;
  wire  ram_sdq_id_T_622_mask;
  wire  ram_sdq_id_T_622_en;
  reg [3:0] T_614;
  reg [31:0] GEN_6;
  reg [3:0] T_616;
  reg [31:0] GEN_7;
  reg  maybe_full;
  reg [31:0] GEN_8;
  wire  ptr_match;
  wire  T_619;
  wire  empty;
  wire  full;
  wire  T_620;
  wire  do_enq;
  wire  T_621;
  wire  do_deq;
  wire [4:0] T_692;
  wire [3:0] T_693;
  wire [3:0] GEN_15;
  wire [4:0] T_697;
  wire [3:0] T_698;
  wire [3:0] GEN_16;
  wire  T_699;
  wire  GEN_17;
  wire  T_701;
  wire  T_703;
  wire [4:0] T_771;
  wire [3:0] ptr_diff;
  wire  T_772;
  wire [4:0] T_773;
  assign io_enq_ready = T_703;
  assign io_deq_valid = T_701;
  assign io_deq_bits_addr = ram_addr_T_704_data;
  assign io_deq_bits_tag = ram_tag_T_704_data;
  assign io_deq_bits_cmd = ram_cmd_T_704_data;
  assign io_deq_bits_typ = ram_typ_T_704_data;
  assign io_deq_bits_phys = ram_phys_T_704_data;
  assign io_deq_bits_sdq_id = ram_sdq_id_T_704_data;
  assign io_count = T_773;
  assign ram_addr_T_704_addr = T_616;
  assign ram_addr_T_704_en = 1'h1;
  assign ram_addr_T_704_data = ram_addr[ram_addr_T_704_addr];
  assign ram_addr_T_622_data = io_enq_bits_addr;
  assign ram_addr_T_622_addr = T_614;
  assign ram_addr_T_622_mask = do_enq;
  assign ram_addr_T_622_en = do_enq;
  assign ram_tag_T_704_addr = T_616;
  assign ram_tag_T_704_en = 1'h1;
  assign ram_tag_T_704_data = ram_tag[ram_tag_T_704_addr];
  assign ram_tag_T_622_data = io_enq_bits_tag;
  assign ram_tag_T_622_addr = T_614;
  assign ram_tag_T_622_mask = do_enq;
  assign ram_tag_T_622_en = do_enq;
  assign ram_cmd_T_704_addr = T_616;
  assign ram_cmd_T_704_en = 1'h1;
  assign ram_cmd_T_704_data = ram_cmd[ram_cmd_T_704_addr];
  assign ram_cmd_T_622_data = io_enq_bits_cmd;
  assign ram_cmd_T_622_addr = T_614;
  assign ram_cmd_T_622_mask = do_enq;
  assign ram_cmd_T_622_en = do_enq;
  assign ram_typ_T_704_addr = T_616;
  assign ram_typ_T_704_en = 1'h1;
  assign ram_typ_T_704_data = ram_typ[ram_typ_T_704_addr];
  assign ram_typ_T_622_data = io_enq_bits_typ;
  assign ram_typ_T_622_addr = T_614;
  assign ram_typ_T_622_mask = do_enq;
  assign ram_typ_T_622_en = do_enq;
  assign ram_phys_T_704_addr = T_616;
  assign ram_phys_T_704_en = 1'h1;
  assign ram_phys_T_704_data = ram_phys[ram_phys_T_704_addr];
  assign ram_phys_T_622_data = io_enq_bits_phys;
  assign ram_phys_T_622_addr = T_614;
  assign ram_phys_T_622_mask = do_enq;
  assign ram_phys_T_622_en = do_enq;
  assign ram_sdq_id_T_704_addr = T_616;
  assign ram_sdq_id_T_704_en = 1'h1;
  assign ram_sdq_id_T_704_data = ram_sdq_id[ram_sdq_id_T_704_addr];
  assign ram_sdq_id_T_622_data = io_enq_bits_sdq_id;
  assign ram_sdq_id_T_622_addr = T_614;
  assign ram_sdq_id_T_622_mask = do_enq;
  assign ram_sdq_id_T_622_en = do_enq;
  assign ptr_match = T_614 == T_616;
  assign T_619 = maybe_full == 1'h0;
  assign empty = ptr_match & T_619;
  assign full = ptr_match & maybe_full;
  assign T_620 = io_enq_ready & io_enq_valid;
  assign do_enq = T_620;
  assign T_621 = io_deq_ready & io_deq_valid;
  assign do_deq = T_621;
  assign T_692 = T_614 + 4'h1;
  assign T_693 = T_692[3:0];
  assign GEN_15 = do_enq ? T_693 : T_614;
  assign T_697 = T_616 + 4'h1;
  assign T_698 = T_697[3:0];
  assign GEN_16 = do_deq ? T_698 : T_616;
  assign T_699 = do_enq != do_deq;
  assign GEN_17 = T_699 ? do_enq : maybe_full;
  assign T_701 = empty == 1'h0;
  assign T_703 = full == 1'h0;
  assign T_771 = T_614 - T_616;
  assign ptr_diff = T_771[3:0];
  assign T_772 = maybe_full & ptr_match;
  assign T_773 = {T_772,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[39:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_tag[initvar] = GEN_1[6:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_cmd[initvar] = GEN_2[4:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_typ[initvar] = GEN_3[2:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_phys[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_sdq_id[initvar] = GEN_5[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_614 = GEN_6[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  T_616 = GEN_7[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  maybe_full = GEN_8[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_622_en & ram_addr_T_622_mask) begin
      ram_addr[ram_addr_T_622_addr] <= ram_addr_T_622_data;
    end
    if(ram_tag_T_622_en & ram_tag_T_622_mask) begin
      ram_tag[ram_tag_T_622_addr] <= ram_tag_T_622_data;
    end
    if(ram_cmd_T_622_en & ram_cmd_T_622_mask) begin
      ram_cmd[ram_cmd_T_622_addr] <= ram_cmd_T_622_data;
    end
    if(ram_typ_T_622_en & ram_typ_T_622_mask) begin
      ram_typ[ram_typ_T_622_addr] <= ram_typ_T_622_data;
    end
    if(ram_phys_T_622_en & ram_phys_T_622_mask) begin
      ram_phys[ram_phys_T_622_addr] <= ram_phys_T_622_data;
    end
    if(ram_sdq_id_T_622_en & ram_sdq_id_T_622_mask) begin
      ram_sdq_id[ram_sdq_id_T_622_addr] <= ram_sdq_id_T_622_data;
    end
    if(reset) begin
      T_614 <= 4'h0;
    end else begin
      if(do_enq) begin
        T_614 <= T_693;
      end
    end
    if(reset) begin
      T_616 <= 4'h0;
    end else begin
      if(do_deq) begin
        T_616 <= T_698;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_699) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module FinishQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output  io_count
);
  reg [2:0] ram_manager_xact_id [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_manager_xact_id_T_254_data;
  wire  ram_manager_xact_id_T_254_addr;
  wire  ram_manager_xact_id_T_254_en;
  wire [2:0] ram_manager_xact_id_T_224_data;
  wire  ram_manager_xact_id_T_224_addr;
  wire  ram_manager_xact_id_T_224_mask;
  wire  ram_manager_xact_id_T_224_en;
  reg  ram_manager_id [0:0];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_254_data;
  wire  ram_manager_id_T_254_addr;
  wire  ram_manager_id_T_254_en;
  wire  ram_manager_id_T_224_data;
  wire  ram_manager_id_T_224_addr;
  wire  ram_manager_id_T_224_mask;
  wire  ram_manager_id_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_2;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_7;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_254_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_254_data;
  assign io_count = T_279[0];
  assign ram_manager_xact_id_T_254_addr = 1'h0;
  assign ram_manager_xact_id_T_254_en = 1'h1;
  assign ram_manager_xact_id_T_254_data = ram_manager_xact_id[ram_manager_xact_id_T_254_addr];
  assign ram_manager_xact_id_T_224_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_224_addr = 1'h0;
  assign ram_manager_xact_id_T_224_mask = do_enq;
  assign ram_manager_xact_id_T_224_en = do_enq;
  assign ram_manager_id_T_254_addr = 1'h0;
  assign ram_manager_id_T_254_en = 1'h1;
  assign ram_manager_id_T_254_data = ram_manager_id[ram_manager_id_T_254_addr];
  assign ram_manager_id_T_224_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_224_addr = 1'h0;
  assign ram_manager_id_T_224_mask = do_enq;
  assign ram_manager_id_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_7 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[2:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  maybe_full = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_224_en & ram_manager_xact_id_T_224_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_224_addr] <= ram_manager_xact_id_T_224_data;
    end
    if(ram_manager_id_T_224_en & ram_manager_id_T_224_mask) begin
      ram_manager_id[ram_manager_id_T_224_addr] <= ram_manager_id_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module MSHR(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [6:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [10:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [6:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_41;
  wire [1:0] T_1659_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_42;
  reg [39:0] req_addr;
  reg [63:0] GEN_43;
  reg [6:0] req_tag;
  reg [31:0] GEN_44;
  reg [4:0] req_cmd;
  reg [31:0] GEN_45;
  reg [2:0] req_typ;
  reg [31:0] GEN_46;
  reg  req_phys;
  reg [31:0] GEN_47;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_48;
  reg  req_tag_match;
  reg [31:0] GEN_49;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_50;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_51;
  reg [3:0] req_way_en;
  reg [31:0] GEN_52;
  wire [5:0] req_idx;
  wire [5:0] T_2007;
  wire  idx_match;
  wire  T_2008;
  wire  T_2009;
  wire  T_2010;
  wire  T_2011;
  wire  T_2012;
  wire  T_2013;
  wire  T_2014;
  wire  T_2015;
  wire  T_2016;
  wire  T_2017;
  wire  T_2018;
  wire  T_2019;
  wire  T_2020;
  wire  T_2021;
  wire  T_2022;
  wire  T_2023;
  wire  T_2024;
  wire  T_2025;
  wire  T_2026;
  wire  T_2027;
  wire  T_2028;
  wire  T_2029;
  wire  T_2031;
  wire  cmd_requires_second_acquire;
  reg  dirties_coh;
  reg [31:0] GEN_53;
  wire [2:0] T_2040_0;
  wire [3:0] GEN_36;
  wire  T_2042;
  wire  T_2043;
  wire  T_2044;
  wire  T_2045;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_54;
  wire  T_2048;
  wire [3:0] T_2050;
  wire [2:0] T_2051;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2053;
  wire  T_2054;
  wire  refill_done;
  wire  T_2055;
  wire  T_2056;
  wire  T_2057;
  wire  T_2058;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire  T_2064;
  wire  T_2065;
  wire  T_2067;
  wire  T_2068;
  wire  T_2069;
  wire  sec_rdy;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [6:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [6:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2137;
  wire  T_2138;
  wire  T_2139;
  wire  T_2140;
  wire  T_2142;
  wire  T_2144;
  wire  T_2145;
  wire  T_2146;
  wire  T_2147;
  wire  T_2148;
  wire  T_2149;
  wire [4:0] T_2150;
  wire  T_2151;
  wire  T_2152;
  wire  T_2153;
  wire  T_2154;
  wire  T_2155;
  wire  T_2156;
  wire  T_2157;
  wire [1:0] T_2158;
  wire [1:0] T_2159;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2210;
  wire [1:0] coh_on_hit_state;
  wire  T_2256;
  wire  T_2257;
  wire [3:0] GEN_1;
  wire  T_2258;
  wire [3:0] GEN_2;
  wire  T_2259;
  wire  T_2260;
  wire [3:0] GEN_3;
  wire  T_2262;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2263;
  wire [3:0] GEN_6;
  wire  T_2265;
  wire [3:0] GEN_7;
  wire  T_2267;
  wire [3:0] GEN_8;
  wire  T_2268;
  wire [3:0] GEN_9;
  wire  T_2273;
  wire [4:0] GEN_10;
  wire  T_2281;
  wire [4:0] GEN_11;
  wire  GEN_12;
  wire  T_2301;
  wire  T_2302;
  wire  T_2303;
  wire  T_2307;
  wire [3:0] GEN_13;
  wire [1:0] GEN_14;
  wire  T_2309;
  wire [3:0] GEN_15;
  wire [3:0] GEN_16;
  wire [1:0] GEN_17;
  wire  T_2311;
  wire [3:0] T_2313;
  wire [3:0] GEN_18;
  wire [39:0] GEN_19;
  wire [6:0] GEN_20;
  wire [4:0] GEN_21;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire [4:0] GEN_24;
  wire  GEN_25;
  wire [19:0] GEN_26;
  wire [1:0] GEN_27;
  wire [3:0] GEN_28;
  wire  GEN_29;
  wire [3:0] GEN_30;
  wire [1:0] GEN_31;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  can_finish;
  wire  T_2344;
  wire  T_2346;
  wire  T_2348;
  wire  T_2349;
  wire [2:0] T_2373_manager_xact_id;
  wire  T_2373_manager_id;
  wire  T_2396;
  wire  T_2397;
  wire  T_2398;
  wire  T_2399;
  wire [8:0] GEN_37;
  wire [8:0] T_2400;
  wire [8:0] GEN_38;
  wire [8:0] T_2401;
  wire [11:0] GEN_39;
  wire [11:0] T_2402;
  wire [27:0] T_2403;
  wire  T_2405;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_55;
  wire  T_2408;
  wire [2:0] T_2410;
  wire [1:0] T_2411;
  wire [1:0] GEN_32;
  wire  T_2412;
  wire [1:0] GEN_33;
  wire  T_2415;
  wire  T_2422;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2431;
  wire [1:0] T_2459_state;
  wire [1:0] T_2481_state;
  wire [25:0] T_2505;
  wire [2:0] T_2510;
  wire [2:0] T_2546_addr_beat;
  wire [25:0] T_2546_addr_block;
  wire [1:0] T_2546_client_xact_id;
  wire  T_2546_voluntary;
  wire [2:0] T_2546_r_type;
  wire [63:0] T_2546_data;
  wire  T_2574;
  wire [25:0] T_2575;
  wire [5:0] T_2591;
  wire [25:0] T_2622_addr_block;
  wire [1:0] T_2622_client_xact_id;
  wire [2:0] T_2622_addr_beat;
  wire  T_2622_is_builtin_type;
  wire [2:0] T_2622_a_type;
  wire [10:0] T_2622_union;
  wire [63:0] T_2622_data;
  wire  T_2652;
  wire [5:0] T_2654;
  wire [31:0] T_2656;
  wire  T_2658;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [3:0] GEN_40;
  reg [31:0] GEN_56;
  Queue rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2148;
  assign io_req_sec_rdy = T_2405;
  assign io_idx_match = T_2399;
  assign io_tag = T_2403[19:0];
  assign io_mem_req_valid = T_2574;
  assign io_mem_req_bits_addr_block = T_2622_addr_block;
  assign io_mem_req_bits_client_xact_id = T_2622_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_2622_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_2622_is_builtin_type;
  assign io_mem_req_bits_a_type = T_2622_a_type;
  assign io_mem_req_bits_union = T_2622_union;
  assign io_mem_req_bits_data = T_2622_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2402;
  assign io_meta_read_valid = T_2146;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_40;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2429;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2481_state;
  assign io_replay_valid = T_2652;
  assign io_replay_bits_addr = {{8'd0}, T_2656};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_35;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2396;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2055;
  assign io_wb_req_bits_addr_beat = T_2546_addr_beat;
  assign io_wb_req_bits_addr_block = T_2546_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2546_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2546_voluntary;
  assign io_wb_req_bits_r_type = T_2546_r_type;
  assign io_wb_req_bits_data = T_2546_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2426;
  assign T_1659_state = 2'h0;
  assign req_idx = req_addr[11:6];
  assign T_2007 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2007;
  assign T_2008 = io_req_bits_cmd == 5'h1;
  assign T_2009 = io_req_bits_cmd == 5'h7;
  assign T_2010 = T_2008 | T_2009;
  assign T_2011 = io_req_bits_cmd[3];
  assign T_2012 = io_req_bits_cmd == 5'h4;
  assign T_2013 = T_2011 | T_2012;
  assign T_2014 = T_2010 | T_2013;
  assign T_2015 = io_req_bits_cmd == 5'h3;
  assign T_2016 = T_2014 | T_2015;
  assign T_2017 = io_req_bits_cmd == 5'h6;
  assign T_2018 = T_2016 | T_2017;
  assign T_2019 = req_cmd == 5'h1;
  assign T_2020 = req_cmd == 5'h7;
  assign T_2021 = T_2019 | T_2020;
  assign T_2022 = req_cmd[3];
  assign T_2023 = req_cmd == 5'h4;
  assign T_2024 = T_2022 | T_2023;
  assign T_2025 = T_2021 | T_2024;
  assign T_2026 = req_cmd == 5'h3;
  assign T_2027 = T_2025 | T_2026;
  assign T_2028 = req_cmd == 5'h6;
  assign T_2029 = T_2027 | T_2028;
  assign T_2031 = T_2029 == 1'h0;
  assign cmd_requires_second_acquire = T_2018 & T_2031;
  assign T_2040_0 = 3'h5;
  assign GEN_36 = {{1'd0}, T_2040_0};
  assign T_2042 = io_mem_grant_bits_g_type == GEN_36;
  assign T_2043 = io_mem_grant_bits_g_type == 4'h0;
  assign T_2044 = io_mem_grant_bits_is_builtin_type ? T_2042 : T_2043;
  assign T_2045 = io_mem_grant_valid & T_2044;
  assign T_2048 = refill_cnt == 3'h7;
  assign T_2050 = refill_cnt + 3'h1;
  assign T_2051 = T_2050[2:0];
  assign GEN_0 = T_2045 ? T_2051 : refill_cnt;
  assign refill_count_done = T_2045 & T_2048;
  assign T_2053 = T_2044 == 1'h0;
  assign T_2054 = T_2053 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2054;
  assign T_2055 = state == 4'h1;
  assign T_2056 = state == 4'h2;
  assign T_2057 = state == 4'h3;
  assign T_2058 = T_2055 | T_2056;
  assign T_2059 = T_2058 | T_2057;
  assign T_2060 = state == 4'h4;
  assign T_2061 = state == 4'h5;
  assign T_2062 = T_2060 | T_2061;
  assign T_2064 = cmd_requires_second_acquire == 1'h0;
  assign T_2065 = T_2062 & T_2064;
  assign T_2067 = refill_done == 1'h0;
  assign T_2068 = T_2065 & T_2067;
  assign T_2069 = T_2059 | T_2068;
  assign sec_rdy = idx_match & T_2069;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2145;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_34;
  assign T_2137 = io_req_pri_val & io_req_pri_rdy;
  assign T_2138 = io_req_sec_val & sec_rdy;
  assign T_2139 = T_2137 | T_2138;
  assign T_2140 = io_req_bits_cmd == 5'h2;
  assign T_2142 = T_2140 | T_2015;
  assign T_2144 = T_2142 == 1'h0;
  assign T_2145 = T_2139 & T_2144;
  assign T_2146 = state == 4'h8;
  assign T_2147 = io_replay_ready & T_2146;
  assign T_2148 = state == 4'h0;
  assign T_2149 = T_2147 | T_2148;
  assign T_2150 = dirties_coh ? 5'h1 : req_cmd;
  assign T_2151 = T_2150 == 5'h1;
  assign T_2152 = T_2150 == 5'h7;
  assign T_2153 = T_2151 | T_2152;
  assign T_2154 = T_2150[3];
  assign T_2155 = T_2150 == 5'h4;
  assign T_2156 = T_2154 | T_2155;
  assign T_2157 = T_2153 | T_2156;
  assign T_2158 = T_2157 ? 2'h2 : 2'h1;
  assign T_2159 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2158;
  assign coh_on_grant_state = T_2159;
  assign T_2210 = T_2014 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2210;
  assign T_2256 = rpq_io_deq_valid == 1'h0;
  assign T_2257 = T_2146 & T_2256;
  assign GEN_1 = T_2257 ? 4'h0 : state;
  assign T_2258 = state == 4'h7;
  assign GEN_2 = T_2258 ? 4'h8 : GEN_1;
  assign T_2259 = state == 4'h6;
  assign T_2260 = T_2259 & io_meta_write_ready;
  assign GEN_3 = T_2260 ? 4'h7 : GEN_2;
  assign T_2262 = T_2061 & refill_done;
  assign GEN_4 = T_2262 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2262 ? coh_on_grant_state : new_coh_state_state;
  assign T_2263 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2263 ? 4'h5 : GEN_4;
  assign T_2265 = T_2057 & io_meta_write_ready;
  assign GEN_7 = T_2265 ? 4'h4 : GEN_6;
  assign T_2267 = T_2056 & io_mem_grant_valid;
  assign GEN_8 = T_2267 ? 4'h3 : GEN_7;
  assign T_2268 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2268 ? 4'h2 : GEN_8;
  assign T_2273 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign T_2281 = dirties_coh | T_2014;
  assign GEN_11 = T_2273 ? GEN_10 : req_cmd;
  assign GEN_12 = T_2273 ? T_2281 : dirties_coh;
  assign T_2301 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T_2302 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T_2303 = T_2301 | T_2302;
  assign T_2307 = T_2018 ? T_2303 : T_2303;
  assign GEN_13 = T_2307 ? 4'h6 : GEN_9;
  assign GEN_14 = T_2307 ? coh_on_hit_state : GEN_5;
  assign T_2309 = T_2307 == 1'h0;
  assign GEN_15 = T_2309 ? 4'h4 : GEN_13;
  assign GEN_16 = io_req_bits_tag_match ? GEN_15 : GEN_9;
  assign GEN_17 = io_req_bits_tag_match ? GEN_14 : GEN_5;
  assign T_2311 = io_req_bits_tag_match == 1'h0;
  assign T_2313 = T_2302 ? 4'h1 : 4'h3;
  assign GEN_18 = T_2311 ? T_2313 : GEN_16;
  assign GEN_19 = T_2137 ? io_req_bits_addr : req_addr;
  assign GEN_20 = T_2137 ? io_req_bits_tag : req_tag;
  assign GEN_21 = T_2137 ? io_req_bits_cmd : GEN_11;
  assign GEN_22 = T_2137 ? io_req_bits_typ : req_typ;
  assign GEN_23 = T_2137 ? io_req_bits_phys : req_phys;
  assign GEN_24 = T_2137 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_25 = T_2137 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_26 = T_2137 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_27 = T_2137 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_28 = T_2137 ? io_req_bits_way_en : req_way_en;
  assign GEN_29 = T_2137 ? T_2014 : GEN_12;
  assign GEN_30 = T_2137 ? GEN_18 : GEN_9;
  assign GEN_31 = T_2137 ? GEN_17 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2349;
  assign fq_io_enq_bits_manager_xact_id = T_2373_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2373_manager_id;
  assign fq_io_deq_ready = T_2397;
  assign can_finish = T_2148 | T_2060;
  assign T_2344 = io_mem_grant_bits_is_builtin_type & T_2043;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2348 = io_mem_grant_valid & T_2346;
  assign T_2349 = T_2348 & refill_done;
  assign T_2373_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2373_manager_id = io_mem_grant_bits_manager_id;
  assign T_2396 = fq_io_deq_valid & can_finish;
  assign T_2397 = io_mem_finish_ready & can_finish;
  assign T_2398 = state != 4'h0;
  assign T_2399 = T_2398 & idx_match;
  assign GEN_37 = {{3'd0}, req_idx};
  assign T_2400 = GEN_37 << 3;
  assign GEN_38 = {{6'd0}, refill_cnt};
  assign T_2401 = T_2400 | GEN_38;
  assign GEN_39 = {{3'd0}, T_2401};
  assign T_2402 = GEN_39 << 3;
  assign T_2403 = req_addr[39:12];
  assign T_2405 = sec_rdy & rpq_io_enq_ready;
  assign T_2408 = meta_hazard != 2'h0;
  assign T_2410 = meta_hazard + 2'h1;
  assign T_2411 = T_2410[1:0];
  assign GEN_32 = T_2408 ? T_2411 : meta_hazard;
  assign T_2412 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_33 = T_2412 ? 2'h1 : GEN_32;
  assign T_2415 = idx_match == 1'h0;
  assign T_2422 = T_2059 == 1'h0;
  assign T_2424 = meta_hazard == 2'h0;
  assign T_2425 = T_2422 & T_2424;
  assign T_2426 = T_2415 | T_2425;
  assign T_2429 = T_2259 | T_2057;
  assign T_2431 = req_old_meta_coh_state == 2'h2;
  assign T_2459_state = 2'h0;
  assign T_2481_state = T_2057 ? T_2459_state : new_coh_state_state;
  assign T_2505 = {req_old_meta_tag,req_idx};
  assign T_2510 = T_2431 ? 3'h0 : 3'h3;
  assign T_2546_addr_beat = 3'h0;
  assign T_2546_addr_block = T_2505;
  assign T_2546_client_xact_id = 2'h0;
  assign T_2546_voluntary = 1'h1;
  assign T_2546_r_type = T_2510;
  assign T_2546_data = 64'h0;
  assign T_2574 = T_2060 & fq_io_enq_ready;
  assign T_2575 = {io_tag,req_idx};
  assign T_2591 = {req_cmd,1'h1};
  assign T_2622_addr_block = T_2575;
  assign T_2622_client_xact_id = 2'h0;
  assign T_2622_addr_beat = 3'h0;
  assign T_2622_is_builtin_type = 1'h0;
  assign T_2622_a_type = {{2'd0}, T_2029};
  assign T_2622_union = {{5'd0}, T_2591};
  assign T_2622_data = 64'h0;
  assign T_2652 = T_2146 & rpq_io_deq_valid;
  assign T_2654 = rpq_io_deq_bits_addr[5:0];
  assign T_2656 = {T_2575,T_2654};
  assign T_2658 = io_meta_read_ready == 1'h0;
  assign GEN_34 = T_2658 ? 1'h0 : T_2149;
  assign GEN_35 = T_2658 ? 5'h5 : rpq_io_deq_bits_cmd;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_56[3:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  state = GEN_41[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  new_coh_state_state = GEN_42[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {2{$random}};
  req_addr = GEN_43[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  req_tag = GEN_44[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  req_cmd = GEN_45[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  req_typ = GEN_46[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  req_phys = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  req_sdq_id = GEN_48[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  req_tag_match = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  req_old_meta_tag = GEN_50[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  req_old_meta_coh_state = GEN_51[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  req_way_en = GEN_52[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  dirties_coh = GEN_53[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  refill_cnt = GEN_54[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  meta_hazard = GEN_55[1:0];
  `endif
  GEN_56 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2137) begin
        if(T_2311) begin
          if(T_2302) begin
            state <= 4'h1;
          end else begin
            state <= 4'h3;
          end
        end else begin
          if(io_req_bits_tag_match) begin
            if(T_2309) begin
              state <= 4'h4;
            end else begin
              if(T_2307) begin
                state <= 4'h6;
              end else begin
                if(T_2268) begin
                  state <= 4'h2;
                end else begin
                  if(T_2267) begin
                    state <= 4'h3;
                  end else begin
                    if(T_2265) begin
                      state <= 4'h4;
                    end else begin
                      if(T_2263) begin
                        state <= 4'h5;
                      end else begin
                        if(T_2262) begin
                          state <= 4'h6;
                        end else begin
                          if(T_2260) begin
                            state <= 4'h7;
                          end else begin
                            if(T_2258) begin
                              state <= 4'h8;
                            end else begin
                              if(T_2257) begin
                                state <= 4'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if(T_2268) begin
              state <= 4'h2;
            end else begin
              if(T_2267) begin
                state <= 4'h3;
              end else begin
                if(T_2265) begin
                  state <= 4'h4;
                end else begin
                  if(T_2263) begin
                    state <= 4'h5;
                  end else begin
                    if(T_2262) begin
                      state <= 4'h6;
                    end else begin
                      if(T_2260) begin
                        state <= 4'h7;
                      end else begin
                        if(T_2258) begin
                          state <= 4'h8;
                        end else begin
                          if(T_2257) begin
                            state <= 4'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if(T_2268) begin
          state <= 4'h2;
        end else begin
          if(T_2267) begin
            state <= 4'h3;
          end else begin
            if(T_2265) begin
              state <= 4'h4;
            end else begin
              if(T_2263) begin
                state <= 4'h5;
              end else begin
                if(T_2262) begin
                  state <= 4'h6;
                end else begin
                  if(T_2260) begin
                    state <= 4'h7;
                  end else begin
                    if(T_2258) begin
                      state <= 4'h8;
                    end else begin
                      if(T_2257) begin
                        state <= 4'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      new_coh_state_state <= T_1659_state;
    end else begin
      if(T_2137) begin
        if(io_req_bits_tag_match) begin
          if(T_2307) begin
            new_coh_state_state <= coh_on_hit_state;
          end else begin
            if(T_2262) begin
              new_coh_state_state <= coh_on_grant_state;
            end
          end
        end else begin
          if(T_2262) begin
            new_coh_state_state <= coh_on_grant_state;
          end
        end
      end else begin
        if(T_2262) begin
          new_coh_state_state <= coh_on_grant_state;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_cmd <= io_req_bits_cmd;
      end else begin
        if(T_2273) begin
          if(cmd_requires_second_acquire) begin
            req_cmd <= io_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_sdq_id <= io_req_bits_sdq_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_tag_match <= io_req_bits_tag_match;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_old_meta_tag <= io_req_bits_old_meta_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        dirties_coh <= T_2014;
      end else begin
        if(T_2273) begin
          dirties_coh <= T_2281;
        end
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_2045) begin
        refill_cnt <= T_2051;
      end
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      if(T_2412) begin
        meta_hazard <= 2'h1;
      end else begin
        if(T_2408) begin
          meta_hazard <= T_2411;
        end
      end
    end
  end
endmodule
module MSHR_1(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [6:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [10:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [6:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_41;
  wire [1:0] T_1659_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_42;
  reg [39:0] req_addr;
  reg [63:0] GEN_43;
  reg [6:0] req_tag;
  reg [31:0] GEN_44;
  reg [4:0] req_cmd;
  reg [31:0] GEN_45;
  reg [2:0] req_typ;
  reg [31:0] GEN_46;
  reg  req_phys;
  reg [31:0] GEN_47;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_48;
  reg  req_tag_match;
  reg [31:0] GEN_49;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_50;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_51;
  reg [3:0] req_way_en;
  reg [31:0] GEN_52;
  wire [5:0] req_idx;
  wire [5:0] T_2007;
  wire  idx_match;
  wire  T_2008;
  wire  T_2009;
  wire  T_2010;
  wire  T_2011;
  wire  T_2012;
  wire  T_2013;
  wire  T_2014;
  wire  T_2015;
  wire  T_2016;
  wire  T_2017;
  wire  T_2018;
  wire  T_2019;
  wire  T_2020;
  wire  T_2021;
  wire  T_2022;
  wire  T_2023;
  wire  T_2024;
  wire  T_2025;
  wire  T_2026;
  wire  T_2027;
  wire  T_2028;
  wire  T_2029;
  wire  T_2031;
  wire  cmd_requires_second_acquire;
  reg  dirties_coh;
  reg [31:0] GEN_53;
  wire [2:0] T_2040_0;
  wire [3:0] GEN_36;
  wire  T_2042;
  wire  T_2043;
  wire  T_2044;
  wire  T_2045;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_54;
  wire  T_2048;
  wire [3:0] T_2050;
  wire [2:0] T_2051;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2053;
  wire  T_2054;
  wire  refill_done;
  wire  T_2055;
  wire  T_2056;
  wire  T_2057;
  wire  T_2058;
  wire  T_2059;
  wire  T_2060;
  wire  T_2061;
  wire  T_2062;
  wire  T_2064;
  wire  T_2065;
  wire  T_2067;
  wire  T_2068;
  wire  T_2069;
  wire  sec_rdy;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [6:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [6:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2137;
  wire  T_2138;
  wire  T_2139;
  wire  T_2140;
  wire  T_2142;
  wire  T_2144;
  wire  T_2145;
  wire  T_2146;
  wire  T_2147;
  wire  T_2148;
  wire  T_2149;
  wire [4:0] T_2150;
  wire  T_2151;
  wire  T_2152;
  wire  T_2153;
  wire  T_2154;
  wire  T_2155;
  wire  T_2156;
  wire  T_2157;
  wire [1:0] T_2158;
  wire [1:0] T_2159;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2210;
  wire [1:0] coh_on_hit_state;
  wire  T_2256;
  wire  T_2257;
  wire [3:0] GEN_1;
  wire  T_2258;
  wire [3:0] GEN_2;
  wire  T_2259;
  wire  T_2260;
  wire [3:0] GEN_3;
  wire  T_2262;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2263;
  wire [3:0] GEN_6;
  wire  T_2265;
  wire [3:0] GEN_7;
  wire  T_2267;
  wire [3:0] GEN_8;
  wire  T_2268;
  wire [3:0] GEN_9;
  wire  T_2273;
  wire [4:0] GEN_10;
  wire  T_2281;
  wire [4:0] GEN_11;
  wire  GEN_12;
  wire  T_2301;
  wire  T_2302;
  wire  T_2303;
  wire  T_2307;
  wire [3:0] GEN_13;
  wire [1:0] GEN_14;
  wire  T_2309;
  wire [3:0] GEN_15;
  wire [3:0] GEN_16;
  wire [1:0] GEN_17;
  wire  T_2311;
  wire [3:0] T_2313;
  wire [3:0] GEN_18;
  wire [39:0] GEN_19;
  wire [6:0] GEN_20;
  wire [4:0] GEN_21;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire [4:0] GEN_24;
  wire  GEN_25;
  wire [19:0] GEN_26;
  wire [1:0] GEN_27;
  wire [3:0] GEN_28;
  wire  GEN_29;
  wire [3:0] GEN_30;
  wire [1:0] GEN_31;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  can_finish;
  wire  T_2344;
  wire  T_2346;
  wire  T_2348;
  wire  T_2349;
  wire [2:0] T_2373_manager_xact_id;
  wire  T_2373_manager_id;
  wire  T_2396;
  wire  T_2397;
  wire  T_2398;
  wire  T_2399;
  wire [8:0] GEN_37;
  wire [8:0] T_2400;
  wire [8:0] GEN_38;
  wire [8:0] T_2401;
  wire [11:0] GEN_39;
  wire [11:0] T_2402;
  wire [27:0] T_2403;
  wire  T_2405;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_55;
  wire  T_2408;
  wire [2:0] T_2410;
  wire [1:0] T_2411;
  wire [1:0] GEN_32;
  wire  T_2412;
  wire [1:0] GEN_33;
  wire  T_2415;
  wire  T_2422;
  wire  T_2424;
  wire  T_2425;
  wire  T_2426;
  wire  T_2429;
  wire  T_2431;
  wire [1:0] T_2459_state;
  wire [1:0] T_2481_state;
  wire [25:0] T_2505;
  wire [2:0] T_2510;
  wire [2:0] T_2546_addr_beat;
  wire [25:0] T_2546_addr_block;
  wire [1:0] T_2546_client_xact_id;
  wire  T_2546_voluntary;
  wire [2:0] T_2546_r_type;
  wire [63:0] T_2546_data;
  wire  T_2574;
  wire [25:0] T_2575;
  wire [5:0] T_2591;
  wire [25:0] T_2622_addr_block;
  wire [1:0] T_2622_client_xact_id;
  wire [2:0] T_2622_addr_beat;
  wire  T_2622_is_builtin_type;
  wire [2:0] T_2622_a_type;
  wire [10:0] T_2622_union;
  wire [63:0] T_2622_data;
  wire  T_2652;
  wire [5:0] T_2654;
  wire [31:0] T_2656;
  wire  T_2658;
  wire  GEN_34;
  wire [4:0] GEN_35;
  wire [3:0] GEN_40;
  reg [31:0] GEN_56;
  Queue rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2148;
  assign io_req_sec_rdy = T_2405;
  assign io_idx_match = T_2399;
  assign io_tag = T_2403[19:0];
  assign io_mem_req_valid = T_2574;
  assign io_mem_req_bits_addr_block = T_2622_addr_block;
  assign io_mem_req_bits_client_xact_id = T_2622_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_2622_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_2622_is_builtin_type;
  assign io_mem_req_bits_a_type = T_2622_a_type;
  assign io_mem_req_bits_union = T_2622_union;
  assign io_mem_req_bits_data = T_2622_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2402;
  assign io_meta_read_valid = T_2146;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_40;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2429;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2481_state;
  assign io_replay_valid = T_2652;
  assign io_replay_bits_addr = {{8'd0}, T_2656};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_35;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2396;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2055;
  assign io_wb_req_bits_addr_beat = T_2546_addr_beat;
  assign io_wb_req_bits_addr_block = T_2546_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2546_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2546_voluntary;
  assign io_wb_req_bits_r_type = T_2546_r_type;
  assign io_wb_req_bits_data = T_2546_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2426;
  assign T_1659_state = 2'h0;
  assign req_idx = req_addr[11:6];
  assign T_2007 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2007;
  assign T_2008 = io_req_bits_cmd == 5'h1;
  assign T_2009 = io_req_bits_cmd == 5'h7;
  assign T_2010 = T_2008 | T_2009;
  assign T_2011 = io_req_bits_cmd[3];
  assign T_2012 = io_req_bits_cmd == 5'h4;
  assign T_2013 = T_2011 | T_2012;
  assign T_2014 = T_2010 | T_2013;
  assign T_2015 = io_req_bits_cmd == 5'h3;
  assign T_2016 = T_2014 | T_2015;
  assign T_2017 = io_req_bits_cmd == 5'h6;
  assign T_2018 = T_2016 | T_2017;
  assign T_2019 = req_cmd == 5'h1;
  assign T_2020 = req_cmd == 5'h7;
  assign T_2021 = T_2019 | T_2020;
  assign T_2022 = req_cmd[3];
  assign T_2023 = req_cmd == 5'h4;
  assign T_2024 = T_2022 | T_2023;
  assign T_2025 = T_2021 | T_2024;
  assign T_2026 = req_cmd == 5'h3;
  assign T_2027 = T_2025 | T_2026;
  assign T_2028 = req_cmd == 5'h6;
  assign T_2029 = T_2027 | T_2028;
  assign T_2031 = T_2029 == 1'h0;
  assign cmd_requires_second_acquire = T_2018 & T_2031;
  assign T_2040_0 = 3'h5;
  assign GEN_36 = {{1'd0}, T_2040_0};
  assign T_2042 = io_mem_grant_bits_g_type == GEN_36;
  assign T_2043 = io_mem_grant_bits_g_type == 4'h0;
  assign T_2044 = io_mem_grant_bits_is_builtin_type ? T_2042 : T_2043;
  assign T_2045 = io_mem_grant_valid & T_2044;
  assign T_2048 = refill_cnt == 3'h7;
  assign T_2050 = refill_cnt + 3'h1;
  assign T_2051 = T_2050[2:0];
  assign GEN_0 = T_2045 ? T_2051 : refill_cnt;
  assign refill_count_done = T_2045 & T_2048;
  assign T_2053 = T_2044 == 1'h0;
  assign T_2054 = T_2053 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2054;
  assign T_2055 = state == 4'h1;
  assign T_2056 = state == 4'h2;
  assign T_2057 = state == 4'h3;
  assign T_2058 = T_2055 | T_2056;
  assign T_2059 = T_2058 | T_2057;
  assign T_2060 = state == 4'h4;
  assign T_2061 = state == 4'h5;
  assign T_2062 = T_2060 | T_2061;
  assign T_2064 = cmd_requires_second_acquire == 1'h0;
  assign T_2065 = T_2062 & T_2064;
  assign T_2067 = refill_done == 1'h0;
  assign T_2068 = T_2065 & T_2067;
  assign T_2069 = T_2059 | T_2068;
  assign sec_rdy = idx_match & T_2069;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2145;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_34;
  assign T_2137 = io_req_pri_val & io_req_pri_rdy;
  assign T_2138 = io_req_sec_val & sec_rdy;
  assign T_2139 = T_2137 | T_2138;
  assign T_2140 = io_req_bits_cmd == 5'h2;
  assign T_2142 = T_2140 | T_2015;
  assign T_2144 = T_2142 == 1'h0;
  assign T_2145 = T_2139 & T_2144;
  assign T_2146 = state == 4'h8;
  assign T_2147 = io_replay_ready & T_2146;
  assign T_2148 = state == 4'h0;
  assign T_2149 = T_2147 | T_2148;
  assign T_2150 = dirties_coh ? 5'h1 : req_cmd;
  assign T_2151 = T_2150 == 5'h1;
  assign T_2152 = T_2150 == 5'h7;
  assign T_2153 = T_2151 | T_2152;
  assign T_2154 = T_2150[3];
  assign T_2155 = T_2150 == 5'h4;
  assign T_2156 = T_2154 | T_2155;
  assign T_2157 = T_2153 | T_2156;
  assign T_2158 = T_2157 ? 2'h2 : 2'h1;
  assign T_2159 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2158;
  assign coh_on_grant_state = T_2159;
  assign T_2210 = T_2014 ? 2'h2 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2210;
  assign T_2256 = rpq_io_deq_valid == 1'h0;
  assign T_2257 = T_2146 & T_2256;
  assign GEN_1 = T_2257 ? 4'h0 : state;
  assign T_2258 = state == 4'h7;
  assign GEN_2 = T_2258 ? 4'h8 : GEN_1;
  assign T_2259 = state == 4'h6;
  assign T_2260 = T_2259 & io_meta_write_ready;
  assign GEN_3 = T_2260 ? 4'h7 : GEN_2;
  assign T_2262 = T_2061 & refill_done;
  assign GEN_4 = T_2262 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2262 ? coh_on_grant_state : new_coh_state_state;
  assign T_2263 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2263 ? 4'h5 : GEN_4;
  assign T_2265 = T_2057 & io_meta_write_ready;
  assign GEN_7 = T_2265 ? 4'h4 : GEN_6;
  assign T_2267 = T_2056 & io_mem_grant_valid;
  assign GEN_8 = T_2267 ? 4'h3 : GEN_7;
  assign T_2268 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2268 ? 4'h2 : GEN_8;
  assign T_2273 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign T_2281 = dirties_coh | T_2014;
  assign GEN_11 = T_2273 ? GEN_10 : req_cmd;
  assign GEN_12 = T_2273 ? T_2281 : dirties_coh;
  assign T_2301 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T_2302 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T_2303 = T_2301 | T_2302;
  assign T_2307 = T_2018 ? T_2303 : T_2303;
  assign GEN_13 = T_2307 ? 4'h6 : GEN_9;
  assign GEN_14 = T_2307 ? coh_on_hit_state : GEN_5;
  assign T_2309 = T_2307 == 1'h0;
  assign GEN_15 = T_2309 ? 4'h4 : GEN_13;
  assign GEN_16 = io_req_bits_tag_match ? GEN_15 : GEN_9;
  assign GEN_17 = io_req_bits_tag_match ? GEN_14 : GEN_5;
  assign T_2311 = io_req_bits_tag_match == 1'h0;
  assign T_2313 = T_2302 ? 4'h1 : 4'h3;
  assign GEN_18 = T_2311 ? T_2313 : GEN_16;
  assign GEN_19 = T_2137 ? io_req_bits_addr : req_addr;
  assign GEN_20 = T_2137 ? io_req_bits_tag : req_tag;
  assign GEN_21 = T_2137 ? io_req_bits_cmd : GEN_11;
  assign GEN_22 = T_2137 ? io_req_bits_typ : req_typ;
  assign GEN_23 = T_2137 ? io_req_bits_phys : req_phys;
  assign GEN_24 = T_2137 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_25 = T_2137 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_26 = T_2137 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_27 = T_2137 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_28 = T_2137 ? io_req_bits_way_en : req_way_en;
  assign GEN_29 = T_2137 ? T_2014 : GEN_12;
  assign GEN_30 = T_2137 ? GEN_18 : GEN_9;
  assign GEN_31 = T_2137 ? GEN_17 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2349;
  assign fq_io_enq_bits_manager_xact_id = T_2373_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2373_manager_id;
  assign fq_io_deq_ready = T_2397;
  assign can_finish = T_2148 | T_2060;
  assign T_2344 = io_mem_grant_bits_is_builtin_type & T_2043;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2348 = io_mem_grant_valid & T_2346;
  assign T_2349 = T_2348 & refill_done;
  assign T_2373_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2373_manager_id = io_mem_grant_bits_manager_id;
  assign T_2396 = fq_io_deq_valid & can_finish;
  assign T_2397 = io_mem_finish_ready & can_finish;
  assign T_2398 = state != 4'h0;
  assign T_2399 = T_2398 & idx_match;
  assign GEN_37 = {{3'd0}, req_idx};
  assign T_2400 = GEN_37 << 3;
  assign GEN_38 = {{6'd0}, refill_cnt};
  assign T_2401 = T_2400 | GEN_38;
  assign GEN_39 = {{3'd0}, T_2401};
  assign T_2402 = GEN_39 << 3;
  assign T_2403 = req_addr[39:12];
  assign T_2405 = sec_rdy & rpq_io_enq_ready;
  assign T_2408 = meta_hazard != 2'h0;
  assign T_2410 = meta_hazard + 2'h1;
  assign T_2411 = T_2410[1:0];
  assign GEN_32 = T_2408 ? T_2411 : meta_hazard;
  assign T_2412 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_33 = T_2412 ? 2'h1 : GEN_32;
  assign T_2415 = idx_match == 1'h0;
  assign T_2422 = T_2059 == 1'h0;
  assign T_2424 = meta_hazard == 2'h0;
  assign T_2425 = T_2422 & T_2424;
  assign T_2426 = T_2415 | T_2425;
  assign T_2429 = T_2259 | T_2057;
  assign T_2431 = req_old_meta_coh_state == 2'h2;
  assign T_2459_state = 2'h0;
  assign T_2481_state = T_2057 ? T_2459_state : new_coh_state_state;
  assign T_2505 = {req_old_meta_tag,req_idx};
  assign T_2510 = T_2431 ? 3'h0 : 3'h3;
  assign T_2546_addr_beat = 3'h0;
  assign T_2546_addr_block = T_2505;
  assign T_2546_client_xact_id = 2'h1;
  assign T_2546_voluntary = 1'h1;
  assign T_2546_r_type = T_2510;
  assign T_2546_data = 64'h0;
  assign T_2574 = T_2060 & fq_io_enq_ready;
  assign T_2575 = {io_tag,req_idx};
  assign T_2591 = {req_cmd,1'h1};
  assign T_2622_addr_block = T_2575;
  assign T_2622_client_xact_id = 2'h1;
  assign T_2622_addr_beat = 3'h0;
  assign T_2622_is_builtin_type = 1'h0;
  assign T_2622_a_type = {{2'd0}, T_2029};
  assign T_2622_union = {{5'd0}, T_2591};
  assign T_2622_data = 64'h0;
  assign T_2652 = T_2146 & rpq_io_deq_valid;
  assign T_2654 = rpq_io_deq_bits_addr[5:0];
  assign T_2656 = {T_2575,T_2654};
  assign T_2658 = io_meta_read_ready == 1'h0;
  assign GEN_34 = T_2658 ? 1'h0 : T_2149;
  assign GEN_35 = T_2658 ? 5'h5 : rpq_io_deq_bits_cmd;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_56[3:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  state = GEN_41[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  new_coh_state_state = GEN_42[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {2{$random}};
  req_addr = GEN_43[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  req_tag = GEN_44[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  req_cmd = GEN_45[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  req_typ = GEN_46[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  req_phys = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  req_sdq_id = GEN_48[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  req_tag_match = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  req_old_meta_tag = GEN_50[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  req_old_meta_coh_state = GEN_51[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  req_way_en = GEN_52[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  dirties_coh = GEN_53[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  refill_cnt = GEN_54[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  meta_hazard = GEN_55[1:0];
  `endif
  GEN_56 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2137) begin
        if(T_2311) begin
          if(T_2302) begin
            state <= 4'h1;
          end else begin
            state <= 4'h3;
          end
        end else begin
          if(io_req_bits_tag_match) begin
            if(T_2309) begin
              state <= 4'h4;
            end else begin
              if(T_2307) begin
                state <= 4'h6;
              end else begin
                if(T_2268) begin
                  state <= 4'h2;
                end else begin
                  if(T_2267) begin
                    state <= 4'h3;
                  end else begin
                    if(T_2265) begin
                      state <= 4'h4;
                    end else begin
                      if(T_2263) begin
                        state <= 4'h5;
                      end else begin
                        if(T_2262) begin
                          state <= 4'h6;
                        end else begin
                          if(T_2260) begin
                            state <= 4'h7;
                          end else begin
                            if(T_2258) begin
                              state <= 4'h8;
                            end else begin
                              if(T_2257) begin
                                state <= 4'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if(T_2268) begin
              state <= 4'h2;
            end else begin
              if(T_2267) begin
                state <= 4'h3;
              end else begin
                if(T_2265) begin
                  state <= 4'h4;
                end else begin
                  if(T_2263) begin
                    state <= 4'h5;
                  end else begin
                    if(T_2262) begin
                      state <= 4'h6;
                    end else begin
                      if(T_2260) begin
                        state <= 4'h7;
                      end else begin
                        if(T_2258) begin
                          state <= 4'h8;
                        end else begin
                          if(T_2257) begin
                            state <= 4'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if(T_2268) begin
          state <= 4'h2;
        end else begin
          if(T_2267) begin
            state <= 4'h3;
          end else begin
            if(T_2265) begin
              state <= 4'h4;
            end else begin
              if(T_2263) begin
                state <= 4'h5;
              end else begin
                if(T_2262) begin
                  state <= 4'h6;
                end else begin
                  if(T_2260) begin
                    state <= 4'h7;
                  end else begin
                    if(T_2258) begin
                      state <= 4'h8;
                    end else begin
                      if(T_2257) begin
                        state <= 4'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      new_coh_state_state <= T_1659_state;
    end else begin
      if(T_2137) begin
        if(io_req_bits_tag_match) begin
          if(T_2307) begin
            new_coh_state_state <= coh_on_hit_state;
          end else begin
            if(T_2262) begin
              new_coh_state_state <= coh_on_grant_state;
            end
          end
        end else begin
          if(T_2262) begin
            new_coh_state_state <= coh_on_grant_state;
          end
        end
      end else begin
        if(T_2262) begin
          new_coh_state_state <= coh_on_grant_state;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_cmd <= io_req_bits_cmd;
      end else begin
        if(T_2273) begin
          if(cmd_requires_second_acquire) begin
            req_cmd <= io_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_sdq_id <= io_req_bits_sdq_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_tag_match <= io_req_bits_tag_match;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_old_meta_tag <= io_req_bits_old_meta_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_old_meta_coh_state <= io_req_bits_old_meta_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        req_way_en <= io_req_bits_way_en;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2137) begin
        dirties_coh <= T_2014;
      end else begin
        if(T_2273) begin
          dirties_coh <= T_2281;
        end
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_2045) begin
        refill_cnt <= T_2051;
      end
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      if(T_2412) begin
        meta_hazard <= 2'h1;
      end else begin
        if(T_2408) begin
          meta_hazard <= T_2411;
        end
      end
    end
  end
endmodule
module Arbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits = io_in_0_bits;
  assign io_chosen = 1'h0;
endmodule
module Arbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [6:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_replay,
  input   io_in_0_bits_has_data,
  input  [63:0] io_in_0_bits_data_word_bypass,
  input  [63:0] io_in_0_bits_store_data,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [6:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output [63:0] io_out_bits_data,
  output  io_out_bits_replay,
  output  io_out_bits_has_data,
  output [63:0] io_out_bits_data_word_bypass,
  output [63:0] io_out_bits_store_data,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_chosen = 1'h0;
endmodule
module IOMSHR(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [6:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_acquire_ready,
  output  io_acquire_valid,
  output [25:0] io_acquire_bits_addr_block,
  output [1:0] io_acquire_bits_client_xact_id,
  output [2:0] io_acquire_bits_addr_beat,
  output  io_acquire_bits_is_builtin_type,
  output [2:0] io_acquire_bits_a_type,
  output [10:0] io_acquire_bits_union,
  output [63:0] io_acquire_bits_data,
  input   io_grant_valid,
  input  [2:0] io_grant_bits_addr_beat,
  input  [1:0] io_grant_bits_client_xact_id,
  input  [2:0] io_grant_bits_manager_xact_id,
  input   io_grant_bits_is_builtin_type,
  input  [3:0] io_grant_bits_g_type,
  input  [63:0] io_grant_bits_data,
  input   io_grant_bits_manager_id,
  input   io_finish_ready,
  output  io_finish_valid,
  output [2:0] io_finish_bits_manager_xact_id,
  output  io_finish_bits_manager_id,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [6:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_replay_next
);
  reg [39:0] req_addr;
  reg [63:0] GEN_16;
  reg [6:0] req_tag;
  reg [31:0] GEN_17;
  reg [4:0] req_cmd;
  reg [31:0] GEN_18;
  reg [2:0] req_typ;
  reg [31:0] GEN_19;
  reg  req_phys;
  reg [31:0] GEN_20;
  reg [63:0] req_data;
  reg [63:0] GEN_21;
  wire  req_cmd_sc;
  reg [63:0] grant_word;
  reg [63:0] GEN_22;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  reg [2:0] state;
  reg [31:0] GEN_23;
  wire  T_1076;
  wire  T_1081;
  wire  T_1082;
  wire  T_1084;
  wire  T_1086;
  wire [2:0] T_1110_manager_xact_id;
  wire  T_1110_manager_id;
  wire  T_1133;
  wire  T_1134;
  wire  T_1136;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  T_1140;
  wire  T_1143;
  wire  T_1147;
  wire  T_1151;
  wire  T_1154;
  wire [1:0] T_1155;
  wire  T_1156;
  wire [1:0] T_1158;
  wire  T_1160;
  wire [1:0] T_1163;
  wire [1:0] T_1164;
  wire [1:0] T_1167;
  wire [3:0] T_1168;
  wire  T_1169;
  wire [3:0] T_1171;
  wire  T_1173;
  wire [3:0] T_1176;
  wire [3:0] T_1177;
  wire [3:0] T_1180;
  wire [7:0] T_1181;
  wire [22:0] GEN_13;
  wire [22:0] beat_mask;
  wire  T_1186;
  wire [7:0] T_1187;
  wire [15:0] T_1188;
  wire [31:0] T_1189;
  wire [63:0] T_1190;
  wire  T_1192;
  wire [15:0] T_1193;
  wire [31:0] T_1194;
  wire [63:0] T_1195;
  wire  T_1197;
  wire [31:0] T_1198;
  wire [63:0] T_1199;
  wire [63:0] T_1200;
  wire [63:0] T_1201;
  wire [63:0] beat_data;
  wire [25:0] addr_block;
  wire [2:0] addr_beat;
  wire [2:0] addr_byte;
  wire [4:0] T_1243;
  wire [10:0] T_1244;
  wire [25:0] get_acquire_addr_block;
  wire [1:0] get_acquire_client_xact_id;
  wire [2:0] get_acquire_addr_beat;
  wire  get_acquire_is_builtin_type;
  wire [2:0] get_acquire_a_type;
  wire [10:0] get_acquire_union;
  wire [63:0] get_acquire_data;
  wire [7:0] T_1367;
  wire [8:0] T_1377;
  wire [10:0] T_1397;
  wire [25:0] put_acquire_addr_block;
  wire [1:0] put_acquire_client_xact_id;
  wire [2:0] put_acquire_addr_beat;
  wire  put_acquire_is_builtin_type;
  wire [2:0] put_acquire_a_type;
  wire [10:0] put_acquire_union;
  wire [63:0] put_acquire_data;
  wire [5:0] T_1496;
  wire [10:0] T_1498;
  wire [25:0] putAtomic_acquire_addr_block;
  wire [1:0] putAtomic_acquire_client_xact_id;
  wire [2:0] putAtomic_acquire_addr_beat;
  wire  putAtomic_acquire_is_builtin_type;
  wire [2:0] putAtomic_acquire_a_type;
  wire [10:0] putAtomic_acquire_union;
  wire [63:0] putAtomic_acquire_data;
  wire  T_1583;
  wire  T_1584;
  wire  T_1585;
  wire  T_1586;
  wire  T_1587;
  wire  T_1588;
  wire  T_1589;
  wire  T_1591;
  wire  T_1595;
  wire [25:0] T_1596_addr_block;
  wire [1:0] T_1596_client_xact_id;
  wire [2:0] T_1596_addr_beat;
  wire  T_1596_is_builtin_type;
  wire [2:0] T_1596_a_type;
  wire [10:0] T_1596_union;
  wire [63:0] T_1596_data;
  wire [25:0] T_1624_addr_block;
  wire [1:0] T_1624_client_xact_id;
  wire [2:0] T_1624_addr_beat;
  wire  T_1624_is_builtin_type;
  wire [2:0] T_1624_a_type;
  wire [10:0] T_1624_union;
  wire [63:0] T_1624_data;
  wire  T_1652;
  wire  T_1654;
  wire  T_1655;
  wire  T_1656;
  wire  T_1657;
  wire [31:0] T_1668;
  wire [31:0] T_1669;
  wire [31:0] T_1670;
  wire  T_1678;
  wire  T_1679;
  wire [31:0] T_1683;
  wire [31:0] T_1685;
  wire [63:0] T_1686;
  wire [15:0] T_1688;
  wire [15:0] T_1689;
  wire [15:0] T_1690;
  wire  T_1698;
  wire  T_1699;
  wire [47:0] T_1703;
  wire [47:0] T_1704;
  wire [47:0] T_1705;
  wire [63:0] T_1706;
  wire [7:0] T_1708;
  wire [7:0] T_1709;
  wire [7:0] T_1710;
  wire [7:0] T_1714;
  wire  T_1717;
  wire  T_1718;
  wire  T_1719;
  wire [55:0] T_1723;
  wire [55:0] T_1724;
  wire [55:0] T_1725;
  wire [63:0] T_1726;
  wire [63:0] GEN_14;
  wire [63:0] T_1727;
  wire  T_1729;
  wire [39:0] GEN_0;
  wire [6:0] GEN_1;
  wire [4:0] GEN_2;
  wire [2:0] GEN_3;
  wire  GEN_4;
  wire [63:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_1730;
  wire [2:0] GEN_7;
  wire  T_1732;
  wire [63:0] T_1745;
  wire [63:0] GEN_8;
  wire [2:0] GEN_9;
  wire [63:0] GEN_10;
  wire  T_1747;
  wire [2:0] GEN_11;
  wire  T_1748;
  wire [2:0] GEN_12;
  wire [63:0] GEN_15;
  reg [63:0] GEN_24;
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_ready = T_1076;
  assign io_acquire_valid = T_1583;
  assign io_acquire_bits_addr_block = T_1624_addr_block;
  assign io_acquire_bits_client_xact_id = T_1624_client_xact_id;
  assign io_acquire_bits_addr_beat = T_1624_addr_beat;
  assign io_acquire_bits_is_builtin_type = T_1624_is_builtin_type;
  assign io_acquire_bits_a_type = T_1624_a_type;
  assign io_acquire_bits_union = T_1624_union;
  assign io_acquire_bits_data = T_1624_data;
  assign io_finish_valid = T_1134;
  assign io_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_resp_valid = T_1657;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_bits_tag = req_tag;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_data = T_1727;
  assign io_resp_bits_replay = 1'h1;
  assign io_resp_bits_has_data = T_1595;
  assign io_resp_bits_data_word_bypass = GEN_15;
  assign io_resp_bits_store_data = req_data;
  assign io_replay_next = T_1656;
  assign req_cmd_sc = req_cmd == 5'h7;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_1086;
  assign fq_io_enq_bits_manager_xact_id = T_1110_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_1110_manager_id;
  assign fq_io_deq_ready = T_1136;
  assign T_1076 = state == 3'h0;
  assign T_1081 = io_grant_bits_g_type == 4'h0;
  assign T_1082 = io_grant_bits_is_builtin_type & T_1081;
  assign T_1084 = T_1082 == 1'h0;
  assign T_1086 = io_grant_valid & T_1084;
  assign T_1110_manager_xact_id = io_grant_bits_manager_xact_id;
  assign T_1110_manager_id = io_grant_bits_manager_id;
  assign T_1133 = state == 3'h4;
  assign T_1134 = fq_io_deq_valid & T_1133;
  assign T_1136 = io_finish_ready & T_1133;
  assign T_1137 = req_typ[1:0];
  assign T_1138 = req_typ[2];
  assign T_1140 = T_1138 == 1'h0;
  assign T_1143 = req_addr[0];
  assign T_1147 = T_1137 >= 2'h1;
  assign T_1151 = T_1143 | T_1147;
  assign T_1154 = T_1143 ? 1'h0 : 1'h1;
  assign T_1155 = {T_1151,T_1154};
  assign T_1156 = req_addr[1];
  assign T_1158 = T_1156 ? T_1155 : 2'h0;
  assign T_1160 = T_1137 >= 2'h2;
  assign T_1163 = T_1160 ? 2'h3 : 2'h0;
  assign T_1164 = T_1158 | T_1163;
  assign T_1167 = T_1156 ? 2'h0 : T_1155;
  assign T_1168 = {T_1164,T_1167};
  assign T_1169 = req_addr[2];
  assign T_1171 = T_1169 ? T_1168 : 4'h0;
  assign T_1173 = T_1137 >= 2'h3;
  assign T_1176 = T_1173 ? 4'hf : 4'h0;
  assign T_1177 = T_1171 | T_1176;
  assign T_1180 = T_1169 ? 4'h0 : T_1168;
  assign T_1181 = {T_1177,T_1180};
  assign GEN_13 = {{15'd0}, T_1181};
  assign beat_mask = GEN_13 << 4'h0;
  assign T_1186 = T_1137 == 2'h0;
  assign T_1187 = req_data[7:0];
  assign T_1188 = {T_1187,T_1187};
  assign T_1189 = {T_1188,T_1188};
  assign T_1190 = {T_1189,T_1189};
  assign T_1192 = T_1137 == 2'h1;
  assign T_1193 = req_data[15:0];
  assign T_1194 = {T_1193,T_1193};
  assign T_1195 = {T_1194,T_1194};
  assign T_1197 = T_1137 == 2'h2;
  assign T_1198 = req_data[31:0];
  assign T_1199 = {T_1198,T_1198};
  assign T_1200 = T_1197 ? T_1199 : req_data;
  assign T_1201 = T_1192 ? T_1195 : T_1200;
  assign beat_data = T_1186 ? T_1190 : T_1201;
  assign addr_block = req_addr[31:6];
  assign addr_beat = req_addr[5:3];
  assign addr_byte = req_addr[2:0];
  assign T_1243 = {addr_byte,T_1137};
  assign T_1244 = {T_1243,6'h0};
  assign get_acquire_addr_block = addr_block;
  assign get_acquire_client_xact_id = 2'h2;
  assign get_acquire_addr_beat = addr_beat;
  assign get_acquire_is_builtin_type = 1'h1;
  assign get_acquire_a_type = 3'h0;
  assign get_acquire_union = T_1244;
  assign get_acquire_data = 64'h0;
  assign T_1367 = beat_mask[7:0];
  assign T_1377 = {T_1367,1'h0};
  assign T_1397 = {{2'd0}, T_1377};
  assign put_acquire_addr_block = addr_block;
  assign put_acquire_client_xact_id = 2'h2;
  assign put_acquire_addr_beat = addr_beat;
  assign put_acquire_is_builtin_type = 1'h1;
  assign put_acquire_a_type = 3'h2;
  assign put_acquire_union = T_1397;
  assign put_acquire_data = beat_data;
  assign T_1496 = {req_cmd,1'h1};
  assign T_1498 = {T_1243,T_1496};
  assign putAtomic_acquire_addr_block = addr_block;
  assign putAtomic_acquire_client_xact_id = 2'h2;
  assign putAtomic_acquire_addr_beat = addr_beat;
  assign putAtomic_acquire_is_builtin_type = 1'h1;
  assign putAtomic_acquire_a_type = 3'h4;
  assign putAtomic_acquire_union = T_1498;
  assign putAtomic_acquire_data = beat_data;
  assign T_1583 = state == 3'h1;
  assign T_1584 = req_cmd[3];
  assign T_1585 = req_cmd == 5'h4;
  assign T_1586 = T_1584 | T_1585;
  assign T_1587 = req_cmd == 5'h0;
  assign T_1588 = req_cmd == 5'h6;
  assign T_1589 = T_1587 | T_1588;
  assign T_1591 = T_1589 | req_cmd_sc;
  assign T_1595 = T_1591 | T_1586;
  assign T_1596_addr_block = T_1595 ? get_acquire_addr_block : put_acquire_addr_block;
  assign T_1596_client_xact_id = T_1595 ? get_acquire_client_xact_id : put_acquire_client_xact_id;
  assign T_1596_addr_beat = T_1595 ? get_acquire_addr_beat : put_acquire_addr_beat;
  assign T_1596_is_builtin_type = T_1595 ? get_acquire_is_builtin_type : put_acquire_is_builtin_type;
  assign T_1596_a_type = T_1595 ? get_acquire_a_type : put_acquire_a_type;
  assign T_1596_union = T_1595 ? get_acquire_union : put_acquire_union;
  assign T_1596_data = T_1595 ? get_acquire_data : put_acquire_data;
  assign T_1624_addr_block = T_1586 ? putAtomic_acquire_addr_block : T_1596_addr_block;
  assign T_1624_client_xact_id = T_1586 ? putAtomic_acquire_client_xact_id : T_1596_client_xact_id;
  assign T_1624_addr_beat = T_1586 ? putAtomic_acquire_addr_beat : T_1596_addr_beat;
  assign T_1624_is_builtin_type = T_1586 ? putAtomic_acquire_is_builtin_type : T_1596_is_builtin_type;
  assign T_1624_a_type = T_1586 ? putAtomic_acquire_a_type : T_1596_a_type;
  assign T_1624_union = T_1586 ? putAtomic_acquire_union : T_1596_union;
  assign T_1624_data = T_1586 ? putAtomic_acquire_data : T_1596_data;
  assign T_1652 = state == 3'h2;
  assign T_1654 = io_resp_ready == 1'h0;
  assign T_1655 = io_resp_valid & T_1654;
  assign T_1656 = T_1652 | T_1655;
  assign T_1657 = state == 3'h3;
  assign T_1668 = grant_word[63:32];
  assign T_1669 = grant_word[31:0];
  assign T_1670 = T_1169 ? T_1668 : T_1669;
  assign T_1678 = T_1670[31];
  assign T_1679 = T_1140 & T_1678;
  assign T_1683 = T_1679 ? 32'hffffffff : 32'h0;
  assign T_1685 = T_1197 ? T_1683 : T_1668;
  assign T_1686 = {T_1685,T_1670};
  assign T_1688 = T_1686[31:16];
  assign T_1689 = T_1686[15:0];
  assign T_1690 = T_1156 ? T_1688 : T_1689;
  assign T_1698 = T_1690[15];
  assign T_1699 = T_1140 & T_1698;
  assign T_1703 = T_1699 ? 48'hffffffffffff : 48'h0;
  assign T_1704 = T_1686[63:16];
  assign T_1705 = T_1192 ? T_1703 : T_1704;
  assign T_1706 = {T_1705,T_1690};
  assign T_1708 = T_1706[15:8];
  assign T_1709 = T_1706[7:0];
  assign T_1710 = T_1143 ? T_1708 : T_1709;
  assign T_1714 = req_cmd_sc ? 8'h0 : T_1710;
  assign T_1717 = T_1186 | req_cmd_sc;
  assign T_1718 = T_1714[7];
  assign T_1719 = T_1140 & T_1718;
  assign T_1723 = T_1719 ? 56'hffffffffffffff : 56'h0;
  assign T_1724 = T_1706[63:8];
  assign T_1725 = T_1717 ? T_1723 : T_1724;
  assign T_1726 = {T_1725,T_1714};
  assign GEN_14 = {{63'd0}, req_cmd_sc};
  assign T_1727 = T_1726 | GEN_14;
  assign T_1729 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1729 ? io_req_bits_addr : req_addr;
  assign GEN_1 = T_1729 ? io_req_bits_tag : req_tag;
  assign GEN_2 = T_1729 ? io_req_bits_cmd : req_cmd;
  assign GEN_3 = T_1729 ? io_req_bits_typ : req_typ;
  assign GEN_4 = T_1729 ? io_req_bits_phys : req_phys;
  assign GEN_5 = T_1729 ? io_req_bits_data : req_data;
  assign GEN_6 = T_1729 ? 3'h1 : state;
  assign T_1730 = io_acquire_ready & io_acquire_valid;
  assign GEN_7 = T_1730 ? 3'h2 : GEN_6;
  assign T_1732 = T_1652 & io_grant_valid;
  assign T_1745 = io_grant_bits_data >> 7'h0;
  assign GEN_8 = T_1595 ? T_1745 : grant_word;
  assign GEN_9 = T_1732 ? 3'h3 : GEN_7;
  assign GEN_10 = T_1732 ? GEN_8 : grant_word;
  assign T_1747 = io_resp_ready & io_resp_valid;
  assign GEN_11 = T_1747 ? 3'h4 : GEN_9;
  assign T_1748 = io_finish_ready & io_finish_valid;
  assign GEN_12 = T_1748 ? 3'h0 : GEN_11;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_24[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {2{$random}};
  req_addr = GEN_16[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  req_tag = GEN_17[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  req_cmd = GEN_18[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_19 = {1{$random}};
  req_typ = GEN_19[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  req_phys = GEN_20[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_21 = {2{$random}};
  req_data = GEN_21[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_22 = {2{$random}};
  grant_word = GEN_22[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_23 = {1{$random}};
  state = GEN_23[2:0];
  `endif
  GEN_24 = {2{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_addr <= io_req_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_cmd <= io_req_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_typ <= io_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_phys <= io_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1729) begin
        req_data <= io_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1732) begin
        if(T_1595) begin
          grant_word <= T_1745;
        end
      end
    end
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_1748) begin
        state <= 3'h0;
      end else begin
        if(T_1747) begin
          state <= 3'h4;
        end else begin
          if(T_1732) begin
            state <= 3'h3;
          end else begin
            if(T_1730) begin
              state <= 3'h2;
            end else begin
              if(T_1729) begin
                state <= 3'h1;
              end
            end
          end
        end
      end
    end
  end
endmodule
module MSHRFile(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [6:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [6:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_secondary_miss,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [10:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [6:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [63:0] io_replay_bits_data,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy,
  output  io_fence_rdy,
  output  io_replay_next
);
  wire  T_2312;
  wire  T_2314;
  wire  T_2315;
  reg [16:0] sdq_val;
  reg [31:0] GEN_5;
  wire [16:0] T_2319;
  wire  T_2320;
  wire  T_2321;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire  T_2328;
  wire  T_2329;
  wire  T_2330;
  wire  T_2331;
  wire  T_2332;
  wire  T_2333;
  wire  T_2334;
  wire  T_2335;
  wire  T_2336;
  wire [4:0] T_2354;
  wire [4:0] T_2355;
  wire [4:0] T_2356;
  wire [4:0] T_2357;
  wire [4:0] T_2358;
  wire [4:0] T_2359;
  wire [4:0] T_2360;
  wire [4:0] T_2361;
  wire [4:0] T_2362;
  wire [4:0] T_2363;
  wire [4:0] T_2364;
  wire [4:0] T_2365;
  wire [4:0] T_2366;
  wire [4:0] T_2367;
  wire [4:0] T_2368;
  wire [4:0] sdq_alloc_id;
  wire  T_2371;
  wire  sdq_rdy;
  wire  T_2373;
  wire  T_2374;
  wire  T_2375;
  wire  T_2376;
  wire  T_2377;
  wire  T_2378;
  wire  T_2379;
  wire  T_2380;
  wire  T_2381;
  wire  sdq_enq;
  reg [63:0] sdq [0:16];
  reg [63:0] GEN_6;
  wire [63:0] sdq_T_3619_data;
  wire [4:0] sdq_T_3619_addr;
  wire  sdq_T_3619_en;
  reg [63:0] GEN_15;
  wire [63:0] sdq_T_2383_data;
  wire [4:0] sdq_T_2383_addr;
  wire  sdq_T_2383_mask;
  wire  sdq_T_2383_en;
  wire  idxMatch_0;
  wire  idxMatch_1;
  wire [19:0] tagList_0;
  wire [19:0] tagList_1;
  wire [19:0] T_2399;
  wire [19:0] T_2401;
  wire [19:0] T_2403;
  wire [19:0] T_2404;
  wire [27:0] T_2405;
  wire [27:0] GEN_0;
  wire  tag_match;
  wire [19:0] wbTagList_0;
  wire [19:0] wbTagList_1;
  wire [3:0] refillMux_0_way_en;
  wire [11:0] refillMux_0_addr;
  wire [3:0] refillMux_1_way_en;
  wire [11:0] refillMux_1_addr;
  wire  meta_read_arb_clk;
  wire  meta_read_arb_reset;
  wire  meta_read_arb_io_in_0_ready;
  wire  meta_read_arb_io_in_0_valid;
  wire [5:0] meta_read_arb_io_in_0_bits_idx;
  wire [3:0] meta_read_arb_io_in_0_bits_way_en;
  wire [19:0] meta_read_arb_io_in_0_bits_tag;
  wire  meta_read_arb_io_in_1_ready;
  wire  meta_read_arb_io_in_1_valid;
  wire [5:0] meta_read_arb_io_in_1_bits_idx;
  wire [3:0] meta_read_arb_io_in_1_bits_way_en;
  wire [19:0] meta_read_arb_io_in_1_bits_tag;
  wire  meta_read_arb_io_out_ready;
  wire  meta_read_arb_io_out_valid;
  wire [5:0] meta_read_arb_io_out_bits_idx;
  wire [3:0] meta_read_arb_io_out_bits_way_en;
  wire [19:0] meta_read_arb_io_out_bits_tag;
  wire  meta_read_arb_io_chosen;
  wire  meta_write_arb_clk;
  wire  meta_write_arb_reset;
  wire  meta_write_arb_io_in_0_ready;
  wire  meta_write_arb_io_in_0_valid;
  wire [5:0] meta_write_arb_io_in_0_bits_idx;
  wire [3:0] meta_write_arb_io_in_0_bits_way_en;
  wire [19:0] meta_write_arb_io_in_0_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_0_bits_data_coh_state;
  wire  meta_write_arb_io_in_1_ready;
  wire  meta_write_arb_io_in_1_valid;
  wire [5:0] meta_write_arb_io_in_1_bits_idx;
  wire [3:0] meta_write_arb_io_in_1_bits_way_en;
  wire [19:0] meta_write_arb_io_in_1_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_1_bits_data_coh_state;
  wire  meta_write_arb_io_out_ready;
  wire  meta_write_arb_io_out_valid;
  wire [5:0] meta_write_arb_io_out_bits_idx;
  wire [3:0] meta_write_arb_io_out_bits_way_en;
  wire [19:0] meta_write_arb_io_out_bits_data_tag;
  wire [1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire  meta_write_arb_io_chosen;
  wire  mem_req_arb_clk;
  wire  mem_req_arb_reset;
  wire  mem_req_arb_io_in_0_ready;
  wire  mem_req_arb_io_in_0_valid;
  wire [25:0] mem_req_arb_io_in_0_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_0_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_0_bits_addr_beat;
  wire  mem_req_arb_io_in_0_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_0_bits_a_type;
  wire [10:0] mem_req_arb_io_in_0_bits_union;
  wire [63:0] mem_req_arb_io_in_0_bits_data;
  wire  mem_req_arb_io_in_1_ready;
  wire  mem_req_arb_io_in_1_valid;
  wire [25:0] mem_req_arb_io_in_1_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_1_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_1_bits_addr_beat;
  wire  mem_req_arb_io_in_1_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_1_bits_a_type;
  wire [10:0] mem_req_arb_io_in_1_bits_union;
  wire [63:0] mem_req_arb_io_in_1_bits_data;
  wire  mem_req_arb_io_in_2_ready;
  wire  mem_req_arb_io_in_2_valid;
  wire [25:0] mem_req_arb_io_in_2_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_2_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_2_bits_addr_beat;
  wire  mem_req_arb_io_in_2_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_2_bits_a_type;
  wire [10:0] mem_req_arb_io_in_2_bits_union;
  wire [63:0] mem_req_arb_io_in_2_bits_data;
  wire  mem_req_arb_io_out_ready;
  wire  mem_req_arb_io_out_valid;
  wire [25:0] mem_req_arb_io_out_bits_addr_block;
  wire [1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_out_bits_addr_beat;
  wire  mem_req_arb_io_out_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_out_bits_a_type;
  wire [10:0] mem_req_arb_io_out_bits_union;
  wire [63:0] mem_req_arb_io_out_bits_data;
  wire [1:0] mem_req_arb_io_chosen;
  wire  mem_finish_arb_clk;
  wire  mem_finish_arb_reset;
  wire  mem_finish_arb_io_in_0_ready;
  wire  mem_finish_arb_io_in_0_valid;
  wire [2:0] mem_finish_arb_io_in_0_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_0_bits_manager_id;
  wire  mem_finish_arb_io_in_1_ready;
  wire  mem_finish_arb_io_in_1_valid;
  wire [2:0] mem_finish_arb_io_in_1_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_1_bits_manager_id;
  wire  mem_finish_arb_io_in_2_ready;
  wire  mem_finish_arb_io_in_2_valid;
  wire [2:0] mem_finish_arb_io_in_2_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_2_bits_manager_id;
  wire  mem_finish_arb_io_out_ready;
  wire  mem_finish_arb_io_out_valid;
  wire [2:0] mem_finish_arb_io_out_bits_manager_xact_id;
  wire  mem_finish_arb_io_out_bits_manager_id;
  wire [1:0] mem_finish_arb_io_chosen;
  wire  wb_req_arb_clk;
  wire  wb_req_arb_reset;
  wire  wb_req_arb_io_in_0_ready;
  wire  wb_req_arb_io_in_0_valid;
  wire [2:0] wb_req_arb_io_in_0_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_0_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_0_bits_client_xact_id;
  wire  wb_req_arb_io_in_0_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_0_bits_r_type;
  wire [63:0] wb_req_arb_io_in_0_bits_data;
  wire [3:0] wb_req_arb_io_in_0_bits_way_en;
  wire  wb_req_arb_io_in_1_ready;
  wire  wb_req_arb_io_in_1_valid;
  wire [2:0] wb_req_arb_io_in_1_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_1_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_1_bits_client_xact_id;
  wire  wb_req_arb_io_in_1_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_1_bits_r_type;
  wire [63:0] wb_req_arb_io_in_1_bits_data;
  wire [3:0] wb_req_arb_io_in_1_bits_way_en;
  wire  wb_req_arb_io_out_ready;
  wire  wb_req_arb_io_out_valid;
  wire [2:0] wb_req_arb_io_out_bits_addr_beat;
  wire [25:0] wb_req_arb_io_out_bits_addr_block;
  wire [1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire  wb_req_arb_io_out_bits_voluntary;
  wire [2:0] wb_req_arb_io_out_bits_r_type;
  wire [63:0] wb_req_arb_io_out_bits_data;
  wire [3:0] wb_req_arb_io_out_bits_way_en;
  wire  wb_req_arb_io_chosen;
  wire  replay_arb_clk;
  wire  replay_arb_reset;
  wire  replay_arb_io_in_0_ready;
  wire  replay_arb_io_in_0_valid;
  wire [39:0] replay_arb_io_in_0_bits_addr;
  wire [6:0] replay_arb_io_in_0_bits_tag;
  wire [4:0] replay_arb_io_in_0_bits_cmd;
  wire [2:0] replay_arb_io_in_0_bits_typ;
  wire  replay_arb_io_in_0_bits_phys;
  wire [4:0] replay_arb_io_in_0_bits_sdq_id;
  wire  replay_arb_io_in_1_ready;
  wire  replay_arb_io_in_1_valid;
  wire [39:0] replay_arb_io_in_1_bits_addr;
  wire [6:0] replay_arb_io_in_1_bits_tag;
  wire [4:0] replay_arb_io_in_1_bits_cmd;
  wire [2:0] replay_arb_io_in_1_bits_typ;
  wire  replay_arb_io_in_1_bits_phys;
  wire [4:0] replay_arb_io_in_1_bits_sdq_id;
  wire  replay_arb_io_out_ready;
  wire  replay_arb_io_out_valid;
  wire [39:0] replay_arb_io_out_bits_addr;
  wire [6:0] replay_arb_io_out_bits_tag;
  wire [4:0] replay_arb_io_out_bits_cmd;
  wire [2:0] replay_arb_io_out_bits_typ;
  wire  replay_arb_io_out_bits_phys;
  wire [4:0] replay_arb_io_out_bits_sdq_id;
  wire  replay_arb_io_chosen;
  wire  alloc_arb_clk;
  wire  alloc_arb_reset;
  wire  alloc_arb_io_in_0_ready;
  wire  alloc_arb_io_in_0_valid;
  wire  alloc_arb_io_in_0_bits;
  wire  alloc_arb_io_in_1_ready;
  wire  alloc_arb_io_in_1_valid;
  wire  alloc_arb_io_in_1_bits;
  wire  alloc_arb_io_out_ready;
  wire  alloc_arb_io_out_valid;
  wire  alloc_arb_io_out_bits;
  wire  alloc_arb_io_chosen;
  wire  MSHR_2_clk;
  wire  MSHR_2_reset;
  wire  MSHR_2_io_req_pri_val;
  wire  MSHR_2_io_req_pri_rdy;
  wire  MSHR_2_io_req_sec_val;
  wire  MSHR_2_io_req_sec_rdy;
  wire [39:0] MSHR_2_io_req_bits_addr;
  wire [6:0] MSHR_2_io_req_bits_tag;
  wire [4:0] MSHR_2_io_req_bits_cmd;
  wire [2:0] MSHR_2_io_req_bits_typ;
  wire  MSHR_2_io_req_bits_phys;
  wire [4:0] MSHR_2_io_req_bits_sdq_id;
  wire  MSHR_2_io_req_bits_tag_match;
  wire [19:0] MSHR_2_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_2_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_2_io_req_bits_way_en;
  wire  MSHR_2_io_idx_match;
  wire [19:0] MSHR_2_io_tag;
  wire  MSHR_2_io_mem_req_ready;
  wire  MSHR_2_io_mem_req_valid;
  wire [25:0] MSHR_2_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_2_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_2_io_mem_req_bits_addr_beat;
  wire  MSHR_2_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_2_io_mem_req_bits_a_type;
  wire [10:0] MSHR_2_io_mem_req_bits_union;
  wire [63:0] MSHR_2_io_mem_req_bits_data;
  wire [3:0] MSHR_2_io_refill_way_en;
  wire [11:0] MSHR_2_io_refill_addr;
  wire  MSHR_2_io_meta_read_ready;
  wire  MSHR_2_io_meta_read_valid;
  wire [5:0] MSHR_2_io_meta_read_bits_idx;
  wire [3:0] MSHR_2_io_meta_read_bits_way_en;
  wire [19:0] MSHR_2_io_meta_read_bits_tag;
  wire  MSHR_2_io_meta_write_ready;
  wire  MSHR_2_io_meta_write_valid;
  wire [5:0] MSHR_2_io_meta_write_bits_idx;
  wire [3:0] MSHR_2_io_meta_write_bits_way_en;
  wire [19:0] MSHR_2_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_2_io_meta_write_bits_data_coh_state;
  wire  MSHR_2_io_replay_ready;
  wire  MSHR_2_io_replay_valid;
  wire [39:0] MSHR_2_io_replay_bits_addr;
  wire [6:0] MSHR_2_io_replay_bits_tag;
  wire [4:0] MSHR_2_io_replay_bits_cmd;
  wire [2:0] MSHR_2_io_replay_bits_typ;
  wire  MSHR_2_io_replay_bits_phys;
  wire [4:0] MSHR_2_io_replay_bits_sdq_id;
  wire  MSHR_2_io_mem_grant_valid;
  wire [2:0] MSHR_2_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_2_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_2_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_2_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_2_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_2_io_mem_grant_bits_data;
  wire  MSHR_2_io_mem_grant_bits_manager_id;
  wire  MSHR_2_io_mem_finish_ready;
  wire  MSHR_2_io_mem_finish_valid;
  wire [2:0] MSHR_2_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_2_io_mem_finish_bits_manager_id;
  wire  MSHR_2_io_wb_req_ready;
  wire  MSHR_2_io_wb_req_valid;
  wire [2:0] MSHR_2_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_2_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_2_io_wb_req_bits_client_xact_id;
  wire  MSHR_2_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_2_io_wb_req_bits_r_type;
  wire [63:0] MSHR_2_io_wb_req_bits_data;
  wire [3:0] MSHR_2_io_wb_req_bits_way_en;
  wire  MSHR_2_io_probe_rdy;
  wire [19:0] T_3427;
  wire  T_3428;
  wire  T_3429;
  wire  T_3431;
  wire  T_3432;
  wire  T_3433;
  wire  T_3434;
  wire  T_3435;
  wire  T_3437;
  wire  GEN_7;
  wire  T_3440;
  wire  GEN_8;
  wire  MSHR_1_1_clk;
  wire  MSHR_1_1_reset;
  wire  MSHR_1_1_io_req_pri_val;
  wire  MSHR_1_1_io_req_pri_rdy;
  wire  MSHR_1_1_io_req_sec_val;
  wire  MSHR_1_1_io_req_sec_rdy;
  wire [39:0] MSHR_1_1_io_req_bits_addr;
  wire [6:0] MSHR_1_1_io_req_bits_tag;
  wire [4:0] MSHR_1_1_io_req_bits_cmd;
  wire [2:0] MSHR_1_1_io_req_bits_typ;
  wire  MSHR_1_1_io_req_bits_phys;
  wire [4:0] MSHR_1_1_io_req_bits_sdq_id;
  wire  MSHR_1_1_io_req_bits_tag_match;
  wire [19:0] MSHR_1_1_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_1_1_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_1_1_io_req_bits_way_en;
  wire  MSHR_1_1_io_idx_match;
  wire [19:0] MSHR_1_1_io_tag;
  wire  MSHR_1_1_io_mem_req_ready;
  wire  MSHR_1_1_io_mem_req_valid;
  wire [25:0] MSHR_1_1_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_1_1_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_1_1_io_mem_req_bits_addr_beat;
  wire  MSHR_1_1_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_1_1_io_mem_req_bits_a_type;
  wire [10:0] MSHR_1_1_io_mem_req_bits_union;
  wire [63:0] MSHR_1_1_io_mem_req_bits_data;
  wire [3:0] MSHR_1_1_io_refill_way_en;
  wire [11:0] MSHR_1_1_io_refill_addr;
  wire  MSHR_1_1_io_meta_read_ready;
  wire  MSHR_1_1_io_meta_read_valid;
  wire [5:0] MSHR_1_1_io_meta_read_bits_idx;
  wire [3:0] MSHR_1_1_io_meta_read_bits_way_en;
  wire [19:0] MSHR_1_1_io_meta_read_bits_tag;
  wire  MSHR_1_1_io_meta_write_ready;
  wire  MSHR_1_1_io_meta_write_valid;
  wire [5:0] MSHR_1_1_io_meta_write_bits_idx;
  wire [3:0] MSHR_1_1_io_meta_write_bits_way_en;
  wire [19:0] MSHR_1_1_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_1_1_io_meta_write_bits_data_coh_state;
  wire  MSHR_1_1_io_replay_ready;
  wire  MSHR_1_1_io_replay_valid;
  wire [39:0] MSHR_1_1_io_replay_bits_addr;
  wire [6:0] MSHR_1_1_io_replay_bits_tag;
  wire [4:0] MSHR_1_1_io_replay_bits_cmd;
  wire [2:0] MSHR_1_1_io_replay_bits_typ;
  wire  MSHR_1_1_io_replay_bits_phys;
  wire [4:0] MSHR_1_1_io_replay_bits_sdq_id;
  wire  MSHR_1_1_io_mem_grant_valid;
  wire [2:0] MSHR_1_1_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_1_1_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_1_1_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_1_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_1_1_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_1_1_io_mem_grant_bits_data;
  wire  MSHR_1_1_io_mem_grant_bits_manager_id;
  wire  MSHR_1_1_io_mem_finish_ready;
  wire  MSHR_1_1_io_mem_finish_valid;
  wire [2:0] MSHR_1_1_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_1_1_io_mem_finish_bits_manager_id;
  wire  MSHR_1_1_io_wb_req_ready;
  wire  MSHR_1_1_io_wb_req_valid;
  wire [2:0] MSHR_1_1_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_1_1_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_1_1_io_wb_req_bits_client_xact_id;
  wire  MSHR_1_1_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_1_1_io_wb_req_bits_r_type;
  wire [63:0] MSHR_1_1_io_wb_req_bits_data;
  wire [3:0] MSHR_1_1_io_wb_req_bits_way_en;
  wire  MSHR_1_1_io_probe_rdy;
  wire [19:0] T_3442;
  wire  T_3446;
  wire  T_3447;
  wire  pri_rdy;
  wire  sec_rdy;
  wire  idx_match;
  wire  T_3449;
  wire  GEN_9;
  wire  T_3452;
  wire  GEN_10;
  wire  T_3455;
  wire  T_3457;
  wire  T_3458;
  wire  mmio_alloc_arb_clk;
  wire  mmio_alloc_arb_reset;
  wire  mmio_alloc_arb_io_in_0_ready;
  wire  mmio_alloc_arb_io_in_0_valid;
  wire  mmio_alloc_arb_io_in_0_bits;
  wire  mmio_alloc_arb_io_out_ready;
  wire  mmio_alloc_arb_io_out_valid;
  wire  mmio_alloc_arb_io_out_bits;
  wire  mmio_alloc_arb_io_chosen;
  wire  resp_arb_clk;
  wire  resp_arb_reset;
  wire  resp_arb_io_in_0_ready;
  wire  resp_arb_io_in_0_valid;
  wire [39:0] resp_arb_io_in_0_bits_addr;
  wire [6:0] resp_arb_io_in_0_bits_tag;
  wire [4:0] resp_arb_io_in_0_bits_cmd;
  wire [2:0] resp_arb_io_in_0_bits_typ;
  wire [63:0] resp_arb_io_in_0_bits_data;
  wire  resp_arb_io_in_0_bits_replay;
  wire  resp_arb_io_in_0_bits_has_data;
  wire [63:0] resp_arb_io_in_0_bits_data_word_bypass;
  wire [63:0] resp_arb_io_in_0_bits_store_data;
  wire  resp_arb_io_out_ready;
  wire  resp_arb_io_out_valid;
  wire [39:0] resp_arb_io_out_bits_addr;
  wire [6:0] resp_arb_io_out_bits_tag;
  wire [4:0] resp_arb_io_out_bits_cmd;
  wire [2:0] resp_arb_io_out_bits_typ;
  wire [63:0] resp_arb_io_out_bits_data;
  wire  resp_arb_io_out_bits_replay;
  wire  resp_arb_io_out_bits_has_data;
  wire [63:0] resp_arb_io_out_bits_data_word_bypass;
  wire [63:0] resp_arb_io_out_bits_store_data;
  wire  resp_arb_io_chosen;
  wire  IOMSHR_1_clk;
  wire  IOMSHR_1_reset;
  wire  IOMSHR_1_io_req_ready;
  wire  IOMSHR_1_io_req_valid;
  wire [39:0] IOMSHR_1_io_req_bits_addr;
  wire [6:0] IOMSHR_1_io_req_bits_tag;
  wire [4:0] IOMSHR_1_io_req_bits_cmd;
  wire [2:0] IOMSHR_1_io_req_bits_typ;
  wire  IOMSHR_1_io_req_bits_phys;
  wire [63:0] IOMSHR_1_io_req_bits_data;
  wire  IOMSHR_1_io_acquire_ready;
  wire  IOMSHR_1_io_acquire_valid;
  wire [25:0] IOMSHR_1_io_acquire_bits_addr_block;
  wire [1:0] IOMSHR_1_io_acquire_bits_client_xact_id;
  wire [2:0] IOMSHR_1_io_acquire_bits_addr_beat;
  wire  IOMSHR_1_io_acquire_bits_is_builtin_type;
  wire [2:0] IOMSHR_1_io_acquire_bits_a_type;
  wire [10:0] IOMSHR_1_io_acquire_bits_union;
  wire [63:0] IOMSHR_1_io_acquire_bits_data;
  wire  IOMSHR_1_io_grant_valid;
  wire [2:0] IOMSHR_1_io_grant_bits_addr_beat;
  wire [1:0] IOMSHR_1_io_grant_bits_client_xact_id;
  wire [2:0] IOMSHR_1_io_grant_bits_manager_xact_id;
  wire  IOMSHR_1_io_grant_bits_is_builtin_type;
  wire [3:0] IOMSHR_1_io_grant_bits_g_type;
  wire [63:0] IOMSHR_1_io_grant_bits_data;
  wire  IOMSHR_1_io_grant_bits_manager_id;
  wire  IOMSHR_1_io_finish_ready;
  wire  IOMSHR_1_io_finish_valid;
  wire [2:0] IOMSHR_1_io_finish_bits_manager_xact_id;
  wire  IOMSHR_1_io_finish_bits_manager_id;
  wire  IOMSHR_1_io_resp_ready;
  wire  IOMSHR_1_io_resp_valid;
  wire [39:0] IOMSHR_1_io_resp_bits_addr;
  wire [6:0] IOMSHR_1_io_resp_bits_tag;
  wire [4:0] IOMSHR_1_io_resp_bits_cmd;
  wire [2:0] IOMSHR_1_io_resp_bits_typ;
  wire [63:0] IOMSHR_1_io_resp_bits_data;
  wire  IOMSHR_1_io_resp_bits_replay;
  wire  IOMSHR_1_io_resp_bits_has_data;
  wire [63:0] IOMSHR_1_io_resp_bits_data_word_bypass;
  wire [63:0] IOMSHR_1_io_resp_bits_store_data;
  wire  IOMSHR_1_io_replay_next;
  wire  mmio_rdy;
  wire  T_3533;
  wire  T_3534;
  wire  T_3536;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_3540;
  wire  T_3541;
  wire  T_3544;
  wire  T_3545;
  wire  T_3546;
  wire  T_3547;
  wire [3:0] GEN_0_way_en;
  wire [11:0] GEN_0_addr;
  wire [3:0] GEN_13;
  wire [11:0] GEN_14;
  wire [3:0] GEN_1_way_en;
  wire [11:0] GEN_1_addr;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire  T_3616;
  wire  T_3617;
  wire  free_sdq;
  reg [4:0] T_3618;
  reg [31:0] GEN_16;
  wire [4:0] GEN_17;
  wire  T_3620;
  wire [31:0] T_3622;
  wire [16:0] T_3626;
  wire [31:0] GEN_1;
  wire [31:0] T_3627;
  wire [31:0] T_3628;
  wire [31:0] GEN_19;
  wire [31:0] T_3629;
  wire [16:0] T_3668;
  wire [16:0] T_3669;
  wire [16:0] T_3670;
  wire [16:0] T_3671;
  wire [16:0] T_3672;
  wire [16:0] T_3673;
  wire [16:0] T_3674;
  wire [16:0] T_3675;
  wire [16:0] T_3676;
  wire [16:0] T_3677;
  wire [16:0] T_3678;
  wire [16:0] T_3679;
  wire [16:0] T_3680;
  wire [16:0] T_3681;
  wire [16:0] T_3682;
  wire [16:0] T_3683;
  wire [16:0] T_3684;
  wire [16:0] T_3688;
  wire [16:0] T_3689;
  wire [31:0] GEN_20;
  wire [31:0] T_3690;
  wire [31:0] GEN_18;
  wire  GEN_2;
  reg [31:0] GEN_21;
  wire  GEN_3;
  reg [31:0] GEN_22;
  wire  GEN_4;
  reg [31:0] GEN_23;
  Arbiter meta_read_arb (
    .clk(meta_read_arb_clk),
    .reset(meta_read_arb_reset),
    .io_in_0_ready(meta_read_arb_io_in_0_ready),
    .io_in_0_valid(meta_read_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_read_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_read_arb_io_in_0_bits_way_en),
    .io_in_0_bits_tag(meta_read_arb_io_in_0_bits_tag),
    .io_in_1_ready(meta_read_arb_io_in_1_ready),
    .io_in_1_valid(meta_read_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_read_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_read_arb_io_in_1_bits_way_en),
    .io_in_1_bits_tag(meta_read_arb_io_in_1_bits_tag),
    .io_out_ready(meta_read_arb_io_out_ready),
    .io_out_valid(meta_read_arb_io_out_valid),
    .io_out_bits_idx(meta_read_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_read_arb_io_out_bits_way_en),
    .io_out_bits_tag(meta_read_arb_io_out_bits_tag),
    .io_chosen(meta_read_arb_io_chosen)
  );
  Arbiter_1 meta_write_arb (
    .clk(meta_write_arb_clk),
    .reset(meta_write_arb_reset),
    .io_in_0_ready(meta_write_arb_io_in_0_ready),
    .io_in_0_valid(meta_write_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_write_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_write_arb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(meta_write_arb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(meta_write_arb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(meta_write_arb_io_in_1_ready),
    .io_in_1_valid(meta_write_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_write_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_write_arb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(meta_write_arb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(meta_write_arb_io_in_1_bits_data_coh_state),
    .io_out_ready(meta_write_arb_io_out_ready),
    .io_out_valid(meta_write_arb_io_out_valid),
    .io_out_bits_idx(meta_write_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_write_arb_io_out_bits_way_en),
    .io_out_bits_data_tag(meta_write_arb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(meta_write_arb_io_out_bits_data_coh_state),
    .io_chosen(meta_write_arb_io_chosen)
  );
  LockingArbiter mem_req_arb (
    .clk(mem_req_arb_clk),
    .reset(mem_req_arb_reset),
    .io_in_0_ready(mem_req_arb_io_in_0_ready),
    .io_in_0_valid(mem_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_block(mem_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(mem_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(mem_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(mem_req_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(mem_req_arb_io_in_0_bits_a_type),
    .io_in_0_bits_union(mem_req_arb_io_in_0_bits_union),
    .io_in_0_bits_data(mem_req_arb_io_in_0_bits_data),
    .io_in_1_ready(mem_req_arb_io_in_1_ready),
    .io_in_1_valid(mem_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_block(mem_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(mem_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(mem_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(mem_req_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(mem_req_arb_io_in_1_bits_a_type),
    .io_in_1_bits_union(mem_req_arb_io_in_1_bits_union),
    .io_in_1_bits_data(mem_req_arb_io_in_1_bits_data),
    .io_in_2_ready(mem_req_arb_io_in_2_ready),
    .io_in_2_valid(mem_req_arb_io_in_2_valid),
    .io_in_2_bits_addr_block(mem_req_arb_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(mem_req_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(mem_req_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(mem_req_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(mem_req_arb_io_in_2_bits_a_type),
    .io_in_2_bits_union(mem_req_arb_io_in_2_bits_union),
    .io_in_2_bits_data(mem_req_arb_io_in_2_bits_data),
    .io_out_ready(mem_req_arb_io_out_ready),
    .io_out_valid(mem_req_arb_io_out_valid),
    .io_out_bits_addr_block(mem_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(mem_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(mem_req_arb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(mem_req_arb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(mem_req_arb_io_out_bits_a_type),
    .io_out_bits_union(mem_req_arb_io_out_bits_union),
    .io_out_bits_data(mem_req_arb_io_out_bits_data),
    .io_chosen(mem_req_arb_io_chosen)
  );
  Arbiter_2 mem_finish_arb (
    .clk(mem_finish_arb_clk),
    .reset(mem_finish_arb_reset),
    .io_in_0_ready(mem_finish_arb_io_in_0_ready),
    .io_in_0_valid(mem_finish_arb_io_in_0_valid),
    .io_in_0_bits_manager_xact_id(mem_finish_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_manager_id(mem_finish_arb_io_in_0_bits_manager_id),
    .io_in_1_ready(mem_finish_arb_io_in_1_ready),
    .io_in_1_valid(mem_finish_arb_io_in_1_valid),
    .io_in_1_bits_manager_xact_id(mem_finish_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_manager_id(mem_finish_arb_io_in_1_bits_manager_id),
    .io_in_2_ready(mem_finish_arb_io_in_2_ready),
    .io_in_2_valid(mem_finish_arb_io_in_2_valid),
    .io_in_2_bits_manager_xact_id(mem_finish_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_manager_id(mem_finish_arb_io_in_2_bits_manager_id),
    .io_out_ready(mem_finish_arb_io_out_ready),
    .io_out_valid(mem_finish_arb_io_out_valid),
    .io_out_bits_manager_xact_id(mem_finish_arb_io_out_bits_manager_xact_id),
    .io_out_bits_manager_id(mem_finish_arb_io_out_bits_manager_id),
    .io_chosen(mem_finish_arb_io_chosen)
  );
  Arbiter_3 wb_req_arb (
    .clk(wb_req_arb_clk),
    .reset(wb_req_arb_reset),
    .io_in_0_ready(wb_req_arb_io_in_0_ready),
    .io_in_0_valid(wb_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wb_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wb_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wb_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wb_req_arb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wb_req_arb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wb_req_arb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wb_req_arb_io_in_0_bits_way_en),
    .io_in_1_ready(wb_req_arb_io_in_1_ready),
    .io_in_1_valid(wb_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wb_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wb_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wb_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wb_req_arb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wb_req_arb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wb_req_arb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wb_req_arb_io_in_1_bits_way_en),
    .io_out_ready(wb_req_arb_io_out_ready),
    .io_out_valid(wb_req_arb_io_out_valid),
    .io_out_bits_addr_beat(wb_req_arb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wb_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wb_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wb_req_arb_io_out_bits_voluntary),
    .io_out_bits_r_type(wb_req_arb_io_out_bits_r_type),
    .io_out_bits_data(wb_req_arb_io_out_bits_data),
    .io_out_bits_way_en(wb_req_arb_io_out_bits_way_en),
    .io_chosen(wb_req_arb_io_chosen)
  );
  Arbiter_4 replay_arb (
    .clk(replay_arb_clk),
    .reset(replay_arb_reset),
    .io_in_0_ready(replay_arb_io_in_0_ready),
    .io_in_0_valid(replay_arb_io_in_0_valid),
    .io_in_0_bits_addr(replay_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(replay_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(replay_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(replay_arb_io_in_0_bits_typ),
    .io_in_0_bits_phys(replay_arb_io_in_0_bits_phys),
    .io_in_0_bits_sdq_id(replay_arb_io_in_0_bits_sdq_id),
    .io_in_1_ready(replay_arb_io_in_1_ready),
    .io_in_1_valid(replay_arb_io_in_1_valid),
    .io_in_1_bits_addr(replay_arb_io_in_1_bits_addr),
    .io_in_1_bits_tag(replay_arb_io_in_1_bits_tag),
    .io_in_1_bits_cmd(replay_arb_io_in_1_bits_cmd),
    .io_in_1_bits_typ(replay_arb_io_in_1_bits_typ),
    .io_in_1_bits_phys(replay_arb_io_in_1_bits_phys),
    .io_in_1_bits_sdq_id(replay_arb_io_in_1_bits_sdq_id),
    .io_out_ready(replay_arb_io_out_ready),
    .io_out_valid(replay_arb_io_out_valid),
    .io_out_bits_addr(replay_arb_io_out_bits_addr),
    .io_out_bits_tag(replay_arb_io_out_bits_tag),
    .io_out_bits_cmd(replay_arb_io_out_bits_cmd),
    .io_out_bits_typ(replay_arb_io_out_bits_typ),
    .io_out_bits_phys(replay_arb_io_out_bits_phys),
    .io_out_bits_sdq_id(replay_arb_io_out_bits_sdq_id),
    .io_chosen(replay_arb_io_chosen)
  );
  Arbiter_5 alloc_arb (
    .clk(alloc_arb_clk),
    .reset(alloc_arb_reset),
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_0_bits(alloc_arb_io_in_0_bits),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_in_1_bits(alloc_arb_io_in_1_bits),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid),
    .io_out_bits(alloc_arb_io_out_bits),
    .io_chosen(alloc_arb_io_chosen)
  );
  MSHR MSHR_2 (
    .clk(MSHR_2_clk),
    .reset(MSHR_2_reset),
    .io_req_pri_val(MSHR_2_io_req_pri_val),
    .io_req_pri_rdy(MSHR_2_io_req_pri_rdy),
    .io_req_sec_val(MSHR_2_io_req_sec_val),
    .io_req_sec_rdy(MSHR_2_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_2_io_req_bits_addr),
    .io_req_bits_tag(MSHR_2_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_2_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_2_io_req_bits_typ),
    .io_req_bits_phys(MSHR_2_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_2_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_2_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_2_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_2_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_2_io_req_bits_way_en),
    .io_idx_match(MSHR_2_io_idx_match),
    .io_tag(MSHR_2_io_tag),
    .io_mem_req_ready(MSHR_2_io_mem_req_ready),
    .io_mem_req_valid(MSHR_2_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_2_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_2_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_2_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_2_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_2_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_2_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_2_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_2_io_refill_way_en),
    .io_refill_addr(MSHR_2_io_refill_addr),
    .io_meta_read_ready(MSHR_2_io_meta_read_ready),
    .io_meta_read_valid(MSHR_2_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_2_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_2_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_2_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_2_io_meta_write_ready),
    .io_meta_write_valid(MSHR_2_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_2_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_2_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_2_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_2_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_2_io_replay_ready),
    .io_replay_valid(MSHR_2_io_replay_valid),
    .io_replay_bits_addr(MSHR_2_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_2_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_2_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_2_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_2_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_2_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_2_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_2_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_2_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_2_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_2_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_2_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_2_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_2_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_2_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_2_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_2_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_2_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_2_io_wb_req_ready),
    .io_wb_req_valid(MSHR_2_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_2_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_2_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_2_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_2_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_2_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_2_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_2_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_2_io_probe_rdy)
  );
  MSHR_1 MSHR_1_1 (
    .clk(MSHR_1_1_clk),
    .reset(MSHR_1_1_reset),
    .io_req_pri_val(MSHR_1_1_io_req_pri_val),
    .io_req_pri_rdy(MSHR_1_1_io_req_pri_rdy),
    .io_req_sec_val(MSHR_1_1_io_req_sec_val),
    .io_req_sec_rdy(MSHR_1_1_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_1_1_io_req_bits_addr),
    .io_req_bits_tag(MSHR_1_1_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_1_1_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_1_1_io_req_bits_typ),
    .io_req_bits_phys(MSHR_1_1_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_1_1_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_1_1_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_1_1_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_1_1_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_1_1_io_req_bits_way_en),
    .io_idx_match(MSHR_1_1_io_idx_match),
    .io_tag(MSHR_1_1_io_tag),
    .io_mem_req_ready(MSHR_1_1_io_mem_req_ready),
    .io_mem_req_valid(MSHR_1_1_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_1_1_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_1_1_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_1_1_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_1_1_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_1_1_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_1_1_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_1_1_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_1_1_io_refill_way_en),
    .io_refill_addr(MSHR_1_1_io_refill_addr),
    .io_meta_read_ready(MSHR_1_1_io_meta_read_ready),
    .io_meta_read_valid(MSHR_1_1_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_1_1_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_1_1_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_1_1_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_1_1_io_meta_write_ready),
    .io_meta_write_valid(MSHR_1_1_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_1_1_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_1_1_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_1_1_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_1_1_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_1_1_io_replay_ready),
    .io_replay_valid(MSHR_1_1_io_replay_valid),
    .io_replay_bits_addr(MSHR_1_1_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_1_1_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_1_1_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_1_1_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_1_1_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_1_1_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_1_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_1_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_1_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_1_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_1_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_1_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_1_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_1_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_1_1_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_1_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_1_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_1_1_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_1_1_io_wb_req_ready),
    .io_wb_req_valid(MSHR_1_1_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_1_1_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_1_1_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_1_1_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_1_1_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_1_1_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_1_1_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_1_1_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_1_1_io_probe_rdy)
  );
  Arbiter_6 mmio_alloc_arb (
    .clk(mmio_alloc_arb_clk),
    .reset(mmio_alloc_arb_reset),
    .io_in_0_ready(mmio_alloc_arb_io_in_0_ready),
    .io_in_0_valid(mmio_alloc_arb_io_in_0_valid),
    .io_in_0_bits(mmio_alloc_arb_io_in_0_bits),
    .io_out_ready(mmio_alloc_arb_io_out_ready),
    .io_out_valid(mmio_alloc_arb_io_out_valid),
    .io_out_bits(mmio_alloc_arb_io_out_bits),
    .io_chosen(mmio_alloc_arb_io_chosen)
  );
  Arbiter_7 resp_arb (
    .clk(resp_arb_clk),
    .reset(resp_arb_reset),
    .io_in_0_ready(resp_arb_io_in_0_ready),
    .io_in_0_valid(resp_arb_io_in_0_valid),
    .io_in_0_bits_addr(resp_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(resp_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(resp_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(resp_arb_io_in_0_bits_typ),
    .io_in_0_bits_data(resp_arb_io_in_0_bits_data),
    .io_in_0_bits_replay(resp_arb_io_in_0_bits_replay),
    .io_in_0_bits_has_data(resp_arb_io_in_0_bits_has_data),
    .io_in_0_bits_data_word_bypass(resp_arb_io_in_0_bits_data_word_bypass),
    .io_in_0_bits_store_data(resp_arb_io_in_0_bits_store_data),
    .io_out_ready(resp_arb_io_out_ready),
    .io_out_valid(resp_arb_io_out_valid),
    .io_out_bits_addr(resp_arb_io_out_bits_addr),
    .io_out_bits_tag(resp_arb_io_out_bits_tag),
    .io_out_bits_cmd(resp_arb_io_out_bits_cmd),
    .io_out_bits_typ(resp_arb_io_out_bits_typ),
    .io_out_bits_data(resp_arb_io_out_bits_data),
    .io_out_bits_replay(resp_arb_io_out_bits_replay),
    .io_out_bits_has_data(resp_arb_io_out_bits_has_data),
    .io_out_bits_data_word_bypass(resp_arb_io_out_bits_data_word_bypass),
    .io_out_bits_store_data(resp_arb_io_out_bits_store_data),
    .io_chosen(resp_arb_io_chosen)
  );
  IOMSHR IOMSHR_1 (
    .clk(IOMSHR_1_clk),
    .reset(IOMSHR_1_reset),
    .io_req_ready(IOMSHR_1_io_req_ready),
    .io_req_valid(IOMSHR_1_io_req_valid),
    .io_req_bits_addr(IOMSHR_1_io_req_bits_addr),
    .io_req_bits_tag(IOMSHR_1_io_req_bits_tag),
    .io_req_bits_cmd(IOMSHR_1_io_req_bits_cmd),
    .io_req_bits_typ(IOMSHR_1_io_req_bits_typ),
    .io_req_bits_phys(IOMSHR_1_io_req_bits_phys),
    .io_req_bits_data(IOMSHR_1_io_req_bits_data),
    .io_acquire_ready(IOMSHR_1_io_acquire_ready),
    .io_acquire_valid(IOMSHR_1_io_acquire_valid),
    .io_acquire_bits_addr_block(IOMSHR_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(IOMSHR_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(IOMSHR_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(IOMSHR_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(IOMSHR_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(IOMSHR_1_io_acquire_bits_union),
    .io_acquire_bits_data(IOMSHR_1_io_acquire_bits_data),
    .io_grant_valid(IOMSHR_1_io_grant_valid),
    .io_grant_bits_addr_beat(IOMSHR_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(IOMSHR_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(IOMSHR_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(IOMSHR_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(IOMSHR_1_io_grant_bits_g_type),
    .io_grant_bits_data(IOMSHR_1_io_grant_bits_data),
    .io_grant_bits_manager_id(IOMSHR_1_io_grant_bits_manager_id),
    .io_finish_ready(IOMSHR_1_io_finish_ready),
    .io_finish_valid(IOMSHR_1_io_finish_valid),
    .io_finish_bits_manager_xact_id(IOMSHR_1_io_finish_bits_manager_xact_id),
    .io_finish_bits_manager_id(IOMSHR_1_io_finish_bits_manager_id),
    .io_resp_ready(IOMSHR_1_io_resp_ready),
    .io_resp_valid(IOMSHR_1_io_resp_valid),
    .io_resp_bits_addr(IOMSHR_1_io_resp_bits_addr),
    .io_resp_bits_tag(IOMSHR_1_io_resp_bits_tag),
    .io_resp_bits_cmd(IOMSHR_1_io_resp_bits_cmd),
    .io_resp_bits_typ(IOMSHR_1_io_resp_bits_typ),
    .io_resp_bits_data(IOMSHR_1_io_resp_bits_data),
    .io_resp_bits_replay(IOMSHR_1_io_resp_bits_replay),
    .io_resp_bits_has_data(IOMSHR_1_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(IOMSHR_1_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(IOMSHR_1_io_resp_bits_store_data),
    .io_replay_next(IOMSHR_1_io_replay_next)
  );
  assign io_req_ready = T_3547;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_secondary_miss = idx_match;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_refill_way_en = GEN_0_way_en;
  assign io_refill_addr = GEN_1_addr;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_bits_way_en = meta_read_arb_io_out_bits_way_en;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_data = sdq_T_3619_data;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_mem_finish_bits_manager_xact_id = mem_finish_arb_io_out_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mem_finish_arb_io_out_bits_manager_id;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_probe_rdy = GEN_10;
  assign io_fence_rdy = GEN_11;
  assign io_replay_next = GEN_12;
  assign T_2312 = 40'h80000000 <= io_req_bits_addr;
  assign T_2314 = io_req_bits_addr < 40'h90000000;
  assign T_2315 = T_2312 & T_2314;
  assign T_2319 = ~ sdq_val;
  assign T_2320 = T_2319[0];
  assign T_2321 = T_2319[1];
  assign T_2322 = T_2319[2];
  assign T_2323 = T_2319[3];
  assign T_2324 = T_2319[4];
  assign T_2325 = T_2319[5];
  assign T_2326 = T_2319[6];
  assign T_2327 = T_2319[7];
  assign T_2328 = T_2319[8];
  assign T_2329 = T_2319[9];
  assign T_2330 = T_2319[10];
  assign T_2331 = T_2319[11];
  assign T_2332 = T_2319[12];
  assign T_2333 = T_2319[13];
  assign T_2334 = T_2319[14];
  assign T_2335 = T_2319[15];
  assign T_2336 = T_2319[16];
  assign T_2354 = T_2335 ? 5'hf : 5'h10;
  assign T_2355 = T_2334 ? 5'he : T_2354;
  assign T_2356 = T_2333 ? 5'hd : T_2355;
  assign T_2357 = T_2332 ? 5'hc : T_2356;
  assign T_2358 = T_2331 ? 5'hb : T_2357;
  assign T_2359 = T_2330 ? 5'ha : T_2358;
  assign T_2360 = T_2329 ? 5'h9 : T_2359;
  assign T_2361 = T_2328 ? 5'h8 : T_2360;
  assign T_2362 = T_2327 ? 5'h7 : T_2361;
  assign T_2363 = T_2326 ? 5'h6 : T_2362;
  assign T_2364 = T_2325 ? 5'h5 : T_2363;
  assign T_2365 = T_2324 ? 5'h4 : T_2364;
  assign T_2366 = T_2323 ? 5'h3 : T_2365;
  assign T_2367 = T_2322 ? 5'h2 : T_2366;
  assign T_2368 = T_2321 ? 5'h1 : T_2367;
  assign sdq_alloc_id = T_2320 ? 5'h0 : T_2368;
  assign T_2371 = T_2319 == 17'h0;
  assign sdq_rdy = T_2371 == 1'h0;
  assign T_2373 = io_req_valid & io_req_ready;
  assign T_2374 = T_2373 & T_2315;
  assign T_2375 = io_req_bits_cmd == 5'h1;
  assign T_2376 = io_req_bits_cmd == 5'h7;
  assign T_2377 = T_2375 | T_2376;
  assign T_2378 = io_req_bits_cmd[3];
  assign T_2379 = io_req_bits_cmd == 5'h4;
  assign T_2380 = T_2378 | T_2379;
  assign T_2381 = T_2377 | T_2380;
  assign sdq_enq = T_2374 & T_2381;
  assign sdq_T_3619_addr = T_3618;
  assign sdq_T_3619_en = 1'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign sdq_T_3619_data = sdq[sdq_T_3619_addr];
  `else
  assign sdq_T_3619_data = sdq_T_3619_addr >= 5'h11 ? GEN_15[63:0] : sdq[sdq_T_3619_addr];
  `endif
  assign sdq_T_2383_data = io_req_bits_data;
  assign sdq_T_2383_addr = sdq_alloc_id;
  assign sdq_T_2383_mask = sdq_enq;
  assign sdq_T_2383_en = sdq_enq;
  assign idxMatch_0 = MSHR_2_io_idx_match;
  assign idxMatch_1 = MSHR_1_1_io_idx_match;
  assign tagList_0 = MSHR_2_io_tag;
  assign tagList_1 = MSHR_1_1_io_tag;
  assign T_2399 = idxMatch_0 ? tagList_0 : 20'h0;
  assign T_2401 = idxMatch_1 ? tagList_1 : 20'h0;
  assign T_2403 = T_2399 | T_2401;
  assign T_2404 = T_2403;
  assign T_2405 = io_req_bits_addr[39:12];
  assign GEN_0 = {{8'd0}, T_2404};
  assign tag_match = GEN_0 == T_2405;
  assign wbTagList_0 = T_3427;
  assign wbTagList_1 = T_3442;
  assign refillMux_0_way_en = MSHR_2_io_refill_way_en;
  assign refillMux_0_addr = MSHR_2_io_refill_addr;
  assign refillMux_1_way_en = MSHR_1_1_io_refill_way_en;
  assign refillMux_1_addr = MSHR_1_1_io_refill_addr;
  assign meta_read_arb_clk = clk;
  assign meta_read_arb_reset = reset;
  assign meta_read_arb_io_in_0_valid = MSHR_2_io_meta_read_valid;
  assign meta_read_arb_io_in_0_bits_idx = MSHR_2_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_0_bits_way_en = MSHR_2_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_0_bits_tag = MSHR_2_io_meta_read_bits_tag;
  assign meta_read_arb_io_in_1_valid = MSHR_1_1_io_meta_read_valid;
  assign meta_read_arb_io_in_1_bits_idx = MSHR_1_1_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_1_bits_way_en = MSHR_1_1_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_1_bits_tag = MSHR_1_1_io_meta_read_bits_tag;
  assign meta_read_arb_io_out_ready = io_meta_read_ready;
  assign meta_write_arb_clk = clk;
  assign meta_write_arb_reset = reset;
  assign meta_write_arb_io_in_0_valid = MSHR_2_io_meta_write_valid;
  assign meta_write_arb_io_in_0_bits_idx = MSHR_2_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_0_bits_way_en = MSHR_2_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_0_bits_data_tag = MSHR_2_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_0_bits_data_coh_state = MSHR_2_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_in_1_valid = MSHR_1_1_io_meta_write_valid;
  assign meta_write_arb_io_in_1_bits_idx = MSHR_1_1_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_1_bits_way_en = MSHR_1_1_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_1_bits_data_tag = MSHR_1_1_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_1_bits_data_coh_state = MSHR_1_1_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_out_ready = io_meta_write_ready;
  assign mem_req_arb_clk = clk;
  assign mem_req_arb_reset = reset;
  assign mem_req_arb_io_in_0_valid = MSHR_2_io_mem_req_valid;
  assign mem_req_arb_io_in_0_bits_addr_block = MSHR_2_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_0_bits_client_xact_id = MSHR_2_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_0_bits_addr_beat = MSHR_2_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_0_bits_is_builtin_type = MSHR_2_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_0_bits_a_type = MSHR_2_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_0_bits_union = MSHR_2_io_mem_req_bits_union;
  assign mem_req_arb_io_in_0_bits_data = MSHR_2_io_mem_req_bits_data;
  assign mem_req_arb_io_in_1_valid = MSHR_1_1_io_mem_req_valid;
  assign mem_req_arb_io_in_1_bits_addr_block = MSHR_1_1_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_1_bits_client_xact_id = MSHR_1_1_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_1_bits_addr_beat = MSHR_1_1_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_1_bits_is_builtin_type = MSHR_1_1_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_1_bits_a_type = MSHR_1_1_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_1_bits_union = MSHR_1_1_io_mem_req_bits_union;
  assign mem_req_arb_io_in_1_bits_data = MSHR_1_1_io_mem_req_bits_data;
  assign mem_req_arb_io_in_2_valid = IOMSHR_1_io_acquire_valid;
  assign mem_req_arb_io_in_2_bits_addr_block = IOMSHR_1_io_acquire_bits_addr_block;
  assign mem_req_arb_io_in_2_bits_client_xact_id = IOMSHR_1_io_acquire_bits_client_xact_id;
  assign mem_req_arb_io_in_2_bits_addr_beat = IOMSHR_1_io_acquire_bits_addr_beat;
  assign mem_req_arb_io_in_2_bits_is_builtin_type = IOMSHR_1_io_acquire_bits_is_builtin_type;
  assign mem_req_arb_io_in_2_bits_a_type = IOMSHR_1_io_acquire_bits_a_type;
  assign mem_req_arb_io_in_2_bits_union = IOMSHR_1_io_acquire_bits_union;
  assign mem_req_arb_io_in_2_bits_data = IOMSHR_1_io_acquire_bits_data;
  assign mem_req_arb_io_out_ready = io_mem_req_ready;
  assign mem_finish_arb_clk = clk;
  assign mem_finish_arb_reset = reset;
  assign mem_finish_arb_io_in_0_valid = MSHR_2_io_mem_finish_valid;
  assign mem_finish_arb_io_in_0_bits_manager_xact_id = MSHR_2_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_0_bits_manager_id = MSHR_2_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_1_valid = MSHR_1_1_io_mem_finish_valid;
  assign mem_finish_arb_io_in_1_bits_manager_xact_id = MSHR_1_1_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_1_bits_manager_id = MSHR_1_1_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_2_valid = IOMSHR_1_io_finish_valid;
  assign mem_finish_arb_io_in_2_bits_manager_xact_id = IOMSHR_1_io_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_2_bits_manager_id = IOMSHR_1_io_finish_bits_manager_id;
  assign mem_finish_arb_io_out_ready = io_mem_finish_ready;
  assign wb_req_arb_clk = clk;
  assign wb_req_arb_reset = reset;
  assign wb_req_arb_io_in_0_valid = MSHR_2_io_wb_req_valid;
  assign wb_req_arb_io_in_0_bits_addr_beat = MSHR_2_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_0_bits_addr_block = MSHR_2_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_0_bits_client_xact_id = MSHR_2_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_0_bits_voluntary = MSHR_2_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_0_bits_r_type = MSHR_2_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_0_bits_data = MSHR_2_io_wb_req_bits_data;
  assign wb_req_arb_io_in_0_bits_way_en = MSHR_2_io_wb_req_bits_way_en;
  assign wb_req_arb_io_in_1_valid = MSHR_1_1_io_wb_req_valid;
  assign wb_req_arb_io_in_1_bits_addr_beat = MSHR_1_1_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_1_bits_addr_block = MSHR_1_1_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_1_bits_client_xact_id = MSHR_1_1_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_1_bits_voluntary = MSHR_1_1_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_1_bits_r_type = MSHR_1_1_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_1_bits_data = MSHR_1_1_io_wb_req_bits_data;
  assign wb_req_arb_io_in_1_bits_way_en = MSHR_1_1_io_wb_req_bits_way_en;
  assign wb_req_arb_io_out_ready = io_wb_req_ready;
  assign replay_arb_clk = clk;
  assign replay_arb_reset = reset;
  assign replay_arb_io_in_0_valid = MSHR_2_io_replay_valid;
  assign replay_arb_io_in_0_bits_addr = MSHR_2_io_replay_bits_addr;
  assign replay_arb_io_in_0_bits_tag = MSHR_2_io_replay_bits_tag;
  assign replay_arb_io_in_0_bits_cmd = MSHR_2_io_replay_bits_cmd;
  assign replay_arb_io_in_0_bits_typ = MSHR_2_io_replay_bits_typ;
  assign replay_arb_io_in_0_bits_phys = MSHR_2_io_replay_bits_phys;
  assign replay_arb_io_in_0_bits_sdq_id = MSHR_2_io_replay_bits_sdq_id;
  assign replay_arb_io_in_1_valid = MSHR_1_1_io_replay_valid;
  assign replay_arb_io_in_1_bits_addr = MSHR_1_1_io_replay_bits_addr;
  assign replay_arb_io_in_1_bits_tag = MSHR_1_1_io_replay_bits_tag;
  assign replay_arb_io_in_1_bits_cmd = MSHR_1_1_io_replay_bits_cmd;
  assign replay_arb_io_in_1_bits_typ = MSHR_1_1_io_replay_bits_typ;
  assign replay_arb_io_in_1_bits_phys = MSHR_1_1_io_replay_bits_phys;
  assign replay_arb_io_in_1_bits_sdq_id = MSHR_1_1_io_replay_bits_sdq_id;
  assign replay_arb_io_out_ready = io_replay_ready;
  assign alloc_arb_clk = clk;
  assign alloc_arb_reset = reset;
  assign alloc_arb_io_in_0_valid = MSHR_2_io_req_pri_rdy;
  assign alloc_arb_io_in_0_bits = GEN_2;
  assign alloc_arb_io_in_1_valid = MSHR_1_1_io_req_pri_rdy;
  assign alloc_arb_io_in_1_bits = GEN_3;
  assign alloc_arb_io_out_ready = T_3458;
  assign MSHR_2_clk = clk;
  assign MSHR_2_reset = reset;
  assign MSHR_2_io_req_pri_val = alloc_arb_io_in_0_ready;
  assign MSHR_2_io_req_sec_val = T_3429;
  assign MSHR_2_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_2_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_2_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_2_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_2_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_2_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_2_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_2_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_2_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_2_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_2_io_mem_req_ready = mem_req_arb_io_in_0_ready;
  assign MSHR_2_io_meta_read_ready = meta_read_arb_io_in_0_ready;
  assign MSHR_2_io_meta_write_ready = meta_write_arb_io_in_0_ready;
  assign MSHR_2_io_replay_ready = replay_arb_io_in_0_ready;
  assign MSHR_2_io_mem_grant_valid = T_3432;
  assign MSHR_2_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_2_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_2_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_2_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_2_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_2_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_2_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_2_io_mem_finish_ready = mem_finish_arb_io_in_0_ready;
  assign MSHR_2_io_wb_req_ready = wb_req_arb_io_in_0_ready;
  assign T_3427 = MSHR_2_io_wb_req_bits_addr_block[25:6];
  assign T_3428 = io_req_valid & sdq_rdy;
  assign T_3429 = T_3428 & tag_match;
  assign T_3431 = io_mem_grant_bits_client_xact_id == 2'h0;
  assign T_3432 = io_mem_grant_valid & T_3431;
  assign T_3433 = MSHR_2_io_req_pri_rdy;
  assign T_3434 = MSHR_2_io_req_sec_rdy;
  assign T_3435 = MSHR_2_io_idx_match;
  assign T_3437 = MSHR_2_io_req_pri_rdy == 1'h0;
  assign GEN_7 = T_3437 ? 1'h0 : 1'h1;
  assign T_3440 = MSHR_2_io_probe_rdy == 1'h0;
  assign GEN_8 = T_3440 ? 1'h0 : 1'h1;
  assign MSHR_1_1_clk = clk;
  assign MSHR_1_1_reset = reset;
  assign MSHR_1_1_io_req_pri_val = alloc_arb_io_in_1_ready;
  assign MSHR_1_1_io_req_sec_val = T_3429;
  assign MSHR_1_1_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_1_1_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_1_1_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_1_1_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_1_1_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_1_1_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_1_1_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_1_1_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_1_1_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_1_1_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_1_1_io_mem_req_ready = mem_req_arb_io_in_1_ready;
  assign MSHR_1_1_io_meta_read_ready = meta_read_arb_io_in_1_ready;
  assign MSHR_1_1_io_meta_write_ready = meta_write_arb_io_in_1_ready;
  assign MSHR_1_1_io_replay_ready = replay_arb_io_in_1_ready;
  assign MSHR_1_1_io_mem_grant_valid = T_3447;
  assign MSHR_1_1_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_1_1_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_1_1_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_1_1_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_1_1_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_1_1_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_1_1_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_1_1_io_mem_finish_ready = mem_finish_arb_io_in_1_ready;
  assign MSHR_1_1_io_wb_req_ready = wb_req_arb_io_in_1_ready;
  assign T_3442 = MSHR_1_1_io_wb_req_bits_addr_block[25:6];
  assign T_3446 = io_mem_grant_bits_client_xact_id == 2'h1;
  assign T_3447 = io_mem_grant_valid & T_3446;
  assign pri_rdy = T_3433 | MSHR_1_1_io_req_pri_rdy;
  assign sec_rdy = T_3434 | MSHR_1_1_io_req_sec_rdy;
  assign idx_match = T_3435 | MSHR_1_1_io_idx_match;
  assign T_3449 = MSHR_1_1_io_req_pri_rdy == 1'h0;
  assign GEN_9 = T_3449 ? 1'h0 : GEN_7;
  assign T_3452 = MSHR_1_1_io_probe_rdy == 1'h0;
  assign GEN_10 = T_3452 ? 1'h0 : GEN_8;
  assign T_3455 = T_3428 & T_2315;
  assign T_3457 = idx_match == 1'h0;
  assign T_3458 = T_3455 & T_3457;
  assign mmio_alloc_arb_clk = clk;
  assign mmio_alloc_arb_reset = reset;
  assign mmio_alloc_arb_io_in_0_valid = IOMSHR_1_io_req_ready;
  assign mmio_alloc_arb_io_in_0_bits = GEN_4;
  assign mmio_alloc_arb_io_out_ready = T_3541;
  assign resp_arb_clk = clk;
  assign resp_arb_reset = reset;
  assign resp_arb_io_in_0_valid = IOMSHR_1_io_resp_valid;
  assign resp_arb_io_in_0_bits_addr = IOMSHR_1_io_resp_bits_addr;
  assign resp_arb_io_in_0_bits_tag = IOMSHR_1_io_resp_bits_tag;
  assign resp_arb_io_in_0_bits_cmd = IOMSHR_1_io_resp_bits_cmd;
  assign resp_arb_io_in_0_bits_typ = IOMSHR_1_io_resp_bits_typ;
  assign resp_arb_io_in_0_bits_data = IOMSHR_1_io_resp_bits_data;
  assign resp_arb_io_in_0_bits_replay = IOMSHR_1_io_resp_bits_replay;
  assign resp_arb_io_in_0_bits_has_data = IOMSHR_1_io_resp_bits_has_data;
  assign resp_arb_io_in_0_bits_data_word_bypass = IOMSHR_1_io_resp_bits_data_word_bypass;
  assign resp_arb_io_in_0_bits_store_data = IOMSHR_1_io_resp_bits_store_data;
  assign resp_arb_io_out_ready = io_resp_ready;
  assign IOMSHR_1_clk = clk;
  assign IOMSHR_1_reset = reset;
  assign IOMSHR_1_io_req_valid = mmio_alloc_arb_io_in_0_ready;
  assign IOMSHR_1_io_req_bits_addr = io_req_bits_addr;
  assign IOMSHR_1_io_req_bits_tag = io_req_bits_tag;
  assign IOMSHR_1_io_req_bits_cmd = io_req_bits_cmd;
  assign IOMSHR_1_io_req_bits_typ = io_req_bits_typ;
  assign IOMSHR_1_io_req_bits_phys = io_req_bits_phys;
  assign IOMSHR_1_io_req_bits_data = io_req_bits_data;
  assign IOMSHR_1_io_acquire_ready = mem_req_arb_io_in_2_ready;
  assign IOMSHR_1_io_grant_valid = T_3534;
  assign IOMSHR_1_io_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign IOMSHR_1_io_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign IOMSHR_1_io_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign IOMSHR_1_io_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign IOMSHR_1_io_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign IOMSHR_1_io_grant_bits_data = io_mem_grant_bits_data;
  assign IOMSHR_1_io_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign IOMSHR_1_io_finish_ready = mem_finish_arb_io_in_2_ready;
  assign IOMSHR_1_io_resp_ready = resp_arb_io_in_0_ready;
  assign mmio_rdy = IOMSHR_1_io_req_ready;
  assign T_3533 = io_mem_grant_bits_client_xact_id == 2'h2;
  assign T_3534 = io_mem_grant_valid & T_3533;
  assign T_3536 = IOMSHR_1_io_req_ready == 1'h0;
  assign GEN_11 = T_3536 ? 1'h0 : GEN_9;
  assign GEN_12 = IOMSHR_1_io_replay_next;
  assign T_3540 = T_2315 == 1'h0;
  assign T_3541 = io_req_valid & T_3540;
  assign T_3544 = tag_match & sec_rdy;
  assign T_3545 = idx_match ? T_3544 : pri_rdy;
  assign T_3546 = T_3545 & sdq_rdy;
  assign T_3547 = T_3540 ? mmio_rdy : T_3546;
  assign GEN_0_way_en = GEN_13;
  assign GEN_0_addr = GEN_14;
  assign GEN_13 = 2'h1 == io_mem_grant_bits_client_xact_id ? refillMux_1_way_en : refillMux_0_way_en;
  assign GEN_14 = 2'h1 == io_mem_grant_bits_client_xact_id ? refillMux_1_addr : refillMux_0_addr;
  assign GEN_1_way_en = GEN_13;
  assign GEN_1_addr = GEN_14;
  assign T_3610 = io_replay_ready & io_replay_valid;
  assign T_3611 = io_replay_bits_cmd == 5'h1;
  assign T_3612 = io_replay_bits_cmd == 5'h7;
  assign T_3613 = T_3611 | T_3612;
  assign T_3614 = io_replay_bits_cmd[3];
  assign T_3615 = io_replay_bits_cmd == 5'h4;
  assign T_3616 = T_3614 | T_3615;
  assign T_3617 = T_3613 | T_3616;
  assign free_sdq = T_3610 & T_3617;
  assign GEN_17 = free_sdq ? replay_arb_io_out_bits_sdq_id : T_3618;
  assign T_3620 = io_replay_valid | sdq_enq;
  assign T_3622 = 32'h1 << replay_arb_io_out_bits_sdq_id;
  assign T_3626 = free_sdq ? 17'h1ffff : 17'h0;
  assign GEN_1 = {{15'd0}, T_3626};
  assign T_3627 = T_3622 & GEN_1;
  assign T_3628 = ~ T_3627;
  assign GEN_19 = {{15'd0}, sdq_val};
  assign T_3629 = GEN_19 & T_3628;
  assign T_3668 = T_2336 ? 17'h10000 : 17'h0;
  assign T_3669 = T_2335 ? 17'h8000 : T_3668;
  assign T_3670 = T_2334 ? 17'h4000 : T_3669;
  assign T_3671 = T_2333 ? 17'h2000 : T_3670;
  assign T_3672 = T_2332 ? 17'h1000 : T_3671;
  assign T_3673 = T_2331 ? 17'h800 : T_3672;
  assign T_3674 = T_2330 ? 17'h400 : T_3673;
  assign T_3675 = T_2329 ? 17'h200 : T_3674;
  assign T_3676 = T_2328 ? 17'h100 : T_3675;
  assign T_3677 = T_2327 ? 17'h80 : T_3676;
  assign T_3678 = T_2326 ? 17'h40 : T_3677;
  assign T_3679 = T_2325 ? 17'h20 : T_3678;
  assign T_3680 = T_2324 ? 17'h10 : T_3679;
  assign T_3681 = T_2323 ? 17'h8 : T_3680;
  assign T_3682 = T_2322 ? 17'h4 : T_3681;
  assign T_3683 = T_2321 ? 17'h2 : T_3682;
  assign T_3684 = T_2320 ? 17'h1 : T_3683;
  assign T_3688 = sdq_enq ? 17'h1ffff : 17'h0;
  assign T_3689 = T_3684 & T_3688;
  assign GEN_20 = {{15'd0}, T_3689};
  assign T_3690 = T_3629 | GEN_20;
  assign GEN_18 = T_3620 ? T_3690 : {{15'd0}, sdq_val};
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_21[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_23[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  sdq_val = GEN_5[16:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    sdq[initvar] = GEN_6[63:0];
  `endif
  GEN_15 = {2{$random}};
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  T_3618 = GEN_16[4:0];
  `endif
  GEN_21 = {1{$random}};
  GEN_22 = {1{$random}};
  GEN_23 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      sdq_val <= 17'h0;
    end else begin
      sdq_val <= GEN_18[16:0];
    end
    if(sdq_T_2383_en & sdq_T_2383_mask) begin
      sdq[sdq_T_2383_addr] <= sdq_T_2383_data;
    end
    if(1'h0) begin
    end else begin
      if(free_sdq) begin
        T_3618 <= replay_arb_io_out_bits_sdq_id;
      end
    end
  end
endmodule
module MetadataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [5:0] io_read_bits_idx,
  input  [3:0] io_read_bits_way_en,
  output  io_write_ready,
  input   io_write_valid,
  input  [5:0] io_write_bits_idx,
  input  [3:0] io_write_bits_way_en,
  input  [19:0] io_write_bits_data_tag,
  input  [1:0] io_write_bits_data_coh_state,
  output [19:0] io_resp_0_tag,
  output [1:0] io_resp_0_coh_state,
  output [19:0] io_resp_1_tag,
  output [1:0] io_resp_1_coh_state,
  output [19:0] io_resp_2_tag,
  output [1:0] io_resp_2_coh_state,
  output [19:0] io_resp_3_tag,
  output [1:0] io_resp_3_coh_state
);
  wire [1:0] T_44_state;
  wire [19:0] rstVal_tag;
  wire [1:0] rstVal_coh_state;
  reg [6:0] rst_cnt;
  reg [31:0] GEN_1;
  wire  rst;
  wire [6:0] waddr;
  wire [19:0] T_2067_tag;
  wire [1:0] T_2067_coh_state;
  wire [21:0] wdata;
  wire [3:0] T_2154;
  wire [3:0] T_2155;
  wire  wmask_0;
  wire  wmask_1;
  wire  wmask_2;
  wire  wmask_3;
  wire [7:0] T_2162;
  wire [6:0] T_2163;
  wire [6:0] GEN_0;
  reg [21:0] T_2172_0 [0:63];
  reg [31:0] GEN_2;
  wire [21:0] T_2172_0_T_2189_data;
  wire [5:0] T_2172_0_T_2189_addr;
  wire  T_2172_0_T_2189_en;
  reg [5:0] GEN_3;
  reg [31:0] GEN_4;
  wire [21:0] T_2172_0_T_2183_data;
  wire [5:0] T_2172_0_T_2183_addr;
  wire  T_2172_0_T_2183_mask;
  wire  T_2172_0_T_2183_en;
  reg [21:0] T_2172_1 [0:63];
  reg [31:0] GEN_5;
  wire [21:0] T_2172_1_T_2189_data;
  wire [5:0] T_2172_1_T_2189_addr;
  wire  T_2172_1_T_2189_en;
  reg [5:0] GEN_6;
  reg [31:0] GEN_7;
  wire [21:0] T_2172_1_T_2183_data;
  wire [5:0] T_2172_1_T_2183_addr;
  wire  T_2172_1_T_2183_mask;
  wire  T_2172_1_T_2183_en;
  reg [21:0] T_2172_2 [0:63];
  reg [31:0] GEN_8;
  wire [21:0] T_2172_2_T_2189_data;
  wire [5:0] T_2172_2_T_2189_addr;
  wire  T_2172_2_T_2189_en;
  reg [5:0] GEN_9;
  reg [31:0] GEN_10;
  wire [21:0] T_2172_2_T_2183_data;
  wire [5:0] T_2172_2_T_2183_addr;
  wire  T_2172_2_T_2183_mask;
  wire  T_2172_2_T_2183_en;
  reg [21:0] T_2172_3 [0:63];
  reg [31:0] GEN_11;
  wire [21:0] T_2172_3_T_2189_data;
  wire [5:0] T_2172_3_T_2189_addr;
  wire  T_2172_3_T_2189_en;
  reg [5:0] GEN_12;
  reg [31:0] GEN_13;
  wire [21:0] T_2172_3_T_2183_data;
  wire [5:0] T_2172_3_T_2183_addr;
  wire  T_2172_3_T_2183_mask;
  wire  T_2172_3_T_2183_en;
  wire  T_2173;
  wire [21:0] T_2179_0;
  wire [21:0] T_2179_1;
  wire [21:0] T_2179_2;
  wire [21:0] T_2179_3;
  wire  GEN_17;
  wire  GEN_19;
  wire  GEN_21;
  wire  GEN_23;
  wire [5:0] T_2186;
  wire [19:0] T_2275_tag;
  wire [1:0] T_2275_coh_state;
  wire [1:0] T_2359;
  wire [19:0] T_2360;
  wire [19:0] T_2445_tag;
  wire [1:0] T_2445_coh_state;
  wire [1:0] T_2529;
  wire [19:0] T_2530;
  wire [19:0] T_2615_tag;
  wire [1:0] T_2615_coh_state;
  wire [1:0] T_2699;
  wire [19:0] T_2700;
  wire [19:0] T_2785_tag;
  wire [1:0] T_2785_coh_state;
  wire [1:0] T_2869;
  wire [19:0] T_2870;
  wire  T_2872;
  wire  T_2874;
  wire  T_2875;
  assign io_read_ready = T_2875;
  assign io_write_ready = T_2872;
  assign io_resp_0_tag = T_2275_tag;
  assign io_resp_0_coh_state = T_2275_coh_state;
  assign io_resp_1_tag = T_2445_tag;
  assign io_resp_1_coh_state = T_2445_coh_state;
  assign io_resp_2_tag = T_2615_tag;
  assign io_resp_2_coh_state = T_2615_coh_state;
  assign io_resp_3_tag = T_2785_tag;
  assign io_resp_3_coh_state = T_2785_coh_state;
  assign T_44_state = 2'h0;
  assign rstVal_tag = 20'h0;
  assign rstVal_coh_state = T_44_state;
  assign rst = rst_cnt < 7'h40;
  assign waddr = rst ? rst_cnt : {{1'd0}, io_write_bits_idx};
  assign T_2067_tag = rst ? rstVal_tag : io_write_bits_data_tag;
  assign T_2067_coh_state = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign wdata = {T_2067_tag,T_2067_coh_state};
  assign T_2154 = $signed(io_write_bits_way_en);
  assign T_2155 = rst ? $signed(4'shf) : $signed(T_2154);
  assign wmask_0 = T_2155[0];
  assign wmask_1 = T_2155[1];
  assign wmask_2 = T_2155[2];
  assign wmask_3 = T_2155[3];
  assign T_2162 = rst_cnt + 7'h1;
  assign T_2163 = T_2162[6:0];
  assign GEN_0 = rst ? T_2163 : rst_cnt;
  assign T_2172_0_T_2189_addr = T_2186;
  assign T_2172_0_T_2189_en = io_read_valid;
  assign T_2172_0_T_2189_data = T_2172_0[GEN_3];
  assign T_2172_0_T_2183_data = T_2179_0;
  assign T_2172_0_T_2183_addr = waddr[5:0];
  assign T_2172_0_T_2183_mask = GEN_17;
  assign T_2172_0_T_2183_en = T_2173;
  assign T_2172_1_T_2189_addr = T_2186;
  assign T_2172_1_T_2189_en = io_read_valid;
  assign T_2172_1_T_2189_data = T_2172_1[GEN_6];
  assign T_2172_1_T_2183_data = T_2179_1;
  assign T_2172_1_T_2183_addr = waddr[5:0];
  assign T_2172_1_T_2183_mask = GEN_19;
  assign T_2172_1_T_2183_en = T_2173;
  assign T_2172_2_T_2189_addr = T_2186;
  assign T_2172_2_T_2189_en = io_read_valid;
  assign T_2172_2_T_2189_data = T_2172_2[GEN_9];
  assign T_2172_2_T_2183_data = T_2179_2;
  assign T_2172_2_T_2183_addr = waddr[5:0];
  assign T_2172_2_T_2183_mask = GEN_21;
  assign T_2172_2_T_2183_en = T_2173;
  assign T_2172_3_T_2189_addr = T_2186;
  assign T_2172_3_T_2189_en = io_read_valid;
  assign T_2172_3_T_2189_data = T_2172_3[GEN_12];
  assign T_2172_3_T_2183_data = T_2179_3;
  assign T_2172_3_T_2183_addr = waddr[5:0];
  assign T_2172_3_T_2183_mask = GEN_23;
  assign T_2172_3_T_2183_en = T_2173;
  assign T_2173 = rst | io_write_valid;
  assign T_2179_0 = wdata;
  assign T_2179_1 = wdata;
  assign T_2179_2 = wdata;
  assign T_2179_3 = wdata;
  assign GEN_17 = T_2173 ? wmask_0 : 1'h0;
  assign GEN_19 = T_2173 ? wmask_1 : 1'h0;
  assign GEN_21 = T_2173 ? wmask_2 : 1'h0;
  assign GEN_23 = T_2173 ? wmask_3 : 1'h0;
  assign T_2186 = io_read_bits_idx;
  assign T_2275_tag = T_2360;
  assign T_2275_coh_state = T_2359;
  assign T_2359 = T_2172_0_T_2189_data[1:0];
  assign T_2360 = T_2172_0_T_2189_data[21:2];
  assign T_2445_tag = T_2530;
  assign T_2445_coh_state = T_2529;
  assign T_2529 = T_2172_1_T_2189_data[1:0];
  assign T_2530 = T_2172_1_T_2189_data[21:2];
  assign T_2615_tag = T_2700;
  assign T_2615_coh_state = T_2699;
  assign T_2699 = T_2172_2_T_2189_data[1:0];
  assign T_2700 = T_2172_2_T_2189_data[21:2];
  assign T_2785_tag = T_2870;
  assign T_2785_coh_state = T_2869;
  assign T_2869 = T_2172_3_T_2189_data[1:0];
  assign T_2870 = T_2172_3_T_2189_data[21:2];
  assign T_2872 = rst == 1'h0;
  assign T_2874 = io_write_valid == 1'h0;
  assign T_2875 = T_2872 & T_2874;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  rst_cnt = GEN_1[6:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2172_0[initvar] = GEN_2[21:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[5:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2172_1[initvar] = GEN_5[21:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  GEN_6 = GEN_7[5:0];
  `endif
  GEN_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2172_2[initvar] = GEN_8[21:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  GEN_9 = GEN_10[5:0];
  `endif
  GEN_11 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2172_3[initvar] = GEN_11[21:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_13 = {1{$random}};
  GEN_12 = GEN_13[5:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else begin
      if(rst) begin
        rst_cnt <= T_2163;
      end
    end
    if(T_2172_0_T_2189_en) begin
      GEN_3 <= T_2172_0_T_2189_addr;
    end
    if(T_2172_0_T_2183_en & T_2172_0_T_2183_mask) begin
      T_2172_0[T_2172_0_T_2183_addr] <= T_2172_0_T_2183_data;
    end
    if(T_2172_1_T_2189_en) begin
      GEN_6 <= T_2172_1_T_2189_addr;
    end
    if(T_2172_1_T_2183_en & T_2172_1_T_2183_mask) begin
      T_2172_1[T_2172_1_T_2183_addr] <= T_2172_1_T_2183_data;
    end
    if(T_2172_2_T_2189_en) begin
      GEN_9 <= T_2172_2_T_2189_addr;
    end
    if(T_2172_2_T_2183_en & T_2172_2_T_2183_mask) begin
      T_2172_2[T_2172_2_T_2183_addr] <= T_2172_2_T_2183_data;
    end
    if(T_2172_3_T_2189_en) begin
      GEN_12 <= T_2172_3_T_2189_addr;
    end
    if(T_2172_3_T_2183_en & T_2172_3_T_2183_mask) begin
      T_2172_3[T_2172_3_T_2183_addr] <= T_2172_3_T_2183_data;
    end
  end
endmodule
module Arbiter_8(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [5:0] io_in_2_bits_idx,
  input  [3:0] io_in_2_bits_way_en,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [5:0] io_in_3_bits_idx,
  input  [3:0] io_in_3_bits_way_en,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [5:0] io_in_4_bits_idx,
  input  [3:0] io_in_4_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [2:0] io_chosen
);
  wire [2:0] GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [2:0] GEN_3;
  wire [5:0] GEN_4;
  wire [3:0] GEN_5;
  wire [2:0] GEN_6;
  wire [5:0] GEN_7;
  wire [3:0] GEN_8;
  wire [2:0] GEN_9;
  wire [5:0] GEN_10;
  wire [3:0] GEN_11;
  wire  T_831;
  wire  T_832;
  wire  T_833;
  wire  grant_1;
  wire  grant_2;
  wire  grant_3;
  wire  grant_4;
  wire  T_839;
  wire  T_840;
  wire  T_841;
  wire  T_842;
  wire  T_844;
  wire  T_845;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_839;
  assign io_in_2_ready = T_840;
  assign io_in_3_ready = T_841;
  assign io_in_4_ready = T_842;
  assign io_out_valid = T_845;
  assign io_out_bits_idx = GEN_10;
  assign io_out_bits_way_en = GEN_11;
  assign io_chosen = GEN_9;
  assign GEN_0 = io_in_3_valid ? 3'h3 : 3'h4;
  assign GEN_1 = io_in_3_valid ? io_in_3_bits_idx : io_in_4_bits_idx;
  assign GEN_2 = io_in_3_valid ? io_in_3_bits_way_en : io_in_4_bits_way_en;
  assign GEN_3 = io_in_2_valid ? 3'h2 : GEN_0;
  assign GEN_4 = io_in_2_valid ? io_in_2_bits_idx : GEN_1;
  assign GEN_5 = io_in_2_valid ? io_in_2_bits_way_en : GEN_2;
  assign GEN_6 = io_in_1_valid ? 3'h1 : GEN_3;
  assign GEN_7 = io_in_1_valid ? io_in_1_bits_idx : GEN_4;
  assign GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : GEN_5;
  assign GEN_9 = io_in_0_valid ? 3'h0 : GEN_6;
  assign GEN_10 = io_in_0_valid ? io_in_0_bits_idx : GEN_7;
  assign GEN_11 = io_in_0_valid ? io_in_0_bits_way_en : GEN_8;
  assign T_831 = io_in_0_valid | io_in_1_valid;
  assign T_832 = T_831 | io_in_2_valid;
  assign T_833 = T_832 | io_in_3_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_831 == 1'h0;
  assign grant_3 = T_832 == 1'h0;
  assign grant_4 = T_833 == 1'h0;
  assign T_839 = grant_1 & io_out_ready;
  assign T_840 = grant_2 & io_out_ready;
  assign T_841 = grant_3 & io_out_ready;
  assign T_842 = grant_4 & io_out_ready;
  assign T_844 = grant_4 == 1'h0;
  assign T_845 = T_844 | io_in_4_valid;
endmodule
module DataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [3:0] io_read_bits_way_en,
  input  [11:0] io_read_bits_addr,
  output  io_write_ready,
  input   io_write_valid,
  input  [3:0] io_write_bits_way_en,
  input  [11:0] io_write_bits_addr,
  input   io_write_bits_wmask,
  input  [63:0] io_write_bits_data,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3
);
  wire [8:0] waddr;
  wire [8:0] raddr;
  wire  T_716;
  wire  T_717;
  wire [63:0] T_724_0;
  reg [11:0] T_726;
  reg [31:0] GEN_1;
  wire [11:0] GEN_0;
  reg [63:0] T_735_0 [0:511];
  reg [63:0] GEN_2;
  wire [63:0] T_735_0_T_761_data;
  wire [8:0] T_735_0_T_761_addr;
  wire  T_735_0_T_761_en;
  reg [8:0] GEN_3;
  reg [31:0] GEN_4;
  wire [63:0] T_735_0_T_752_data;
  wire [8:0] T_735_0_T_752_addr;
  wire  T_735_0_T_752_mask;
  wire  T_735_0_T_752_en;
  wire  T_738;
  wire  T_740;
  wire [63:0] T_747_0;
  wire  GEN_8;
  wire  T_756;
  wire [8:0] T_758;
  wire [63:0] T_769_0;
  wire  T_771;
  wire  T_772;
  wire [63:0] T_779_0;
  reg [11:0] T_781;
  reg [31:0] GEN_5;
  wire [11:0] GEN_11;
  reg [63:0] T_790_0 [0:511];
  reg [63:0] GEN_6;
  wire [63:0] T_790_0_T_816_data;
  wire [8:0] T_790_0_T_816_addr;
  wire  T_790_0_T_816_en;
  reg [8:0] GEN_7;
  reg [31:0] GEN_9;
  wire [63:0] T_790_0_T_807_data;
  wire [8:0] T_790_0_T_807_addr;
  wire  T_790_0_T_807_mask;
  wire  T_790_0_T_807_en;
  wire  T_793;
  wire  T_795;
  wire [63:0] T_802_0;
  wire  GEN_19;
  wire  T_811;
  wire [8:0] T_813;
  wire [63:0] T_824_0;
  wire  T_826;
  wire  T_827;
  wire [63:0] T_834_0;
  reg [11:0] T_836;
  reg [31:0] GEN_10;
  wire [11:0] GEN_22;
  reg [63:0] T_845_0 [0:511];
  reg [63:0] GEN_12;
  wire [63:0] T_845_0_T_871_data;
  wire [8:0] T_845_0_T_871_addr;
  wire  T_845_0_T_871_en;
  reg [8:0] GEN_13;
  reg [31:0] GEN_14;
  wire [63:0] T_845_0_T_862_data;
  wire [8:0] T_845_0_T_862_addr;
  wire  T_845_0_T_862_mask;
  wire  T_845_0_T_862_en;
  wire  T_848;
  wire  T_850;
  wire [63:0] T_857_0;
  wire  GEN_30;
  wire  T_866;
  wire [8:0] T_868;
  wire [63:0] T_879_0;
  wire  T_881;
  wire  T_882;
  wire [63:0] T_889_0;
  reg [11:0] T_891;
  reg [31:0] GEN_15;
  wire [11:0] GEN_33;
  reg [63:0] T_900_0 [0:511];
  reg [63:0] GEN_16;
  wire [63:0] T_900_0_T_926_data;
  wire [8:0] T_900_0_T_926_addr;
  wire  T_900_0_T_926_en;
  reg [8:0] GEN_17;
  reg [31:0] GEN_18;
  wire [63:0] T_900_0_T_917_data;
  wire [8:0] T_900_0_T_917_addr;
  wire  T_900_0_T_917_mask;
  wire  T_900_0_T_917_en;
  wire  T_903;
  wire  T_905;
  wire [63:0] T_912_0;
  wire  GEN_41;
  wire  T_921;
  wire [8:0] T_923;
  wire [63:0] T_934_0;
  assign io_read_ready = 1'h1;
  assign io_write_ready = 1'h1;
  assign io_resp_0 = T_769_0;
  assign io_resp_1 = T_824_0;
  assign io_resp_2 = T_879_0;
  assign io_resp_3 = T_934_0;
  assign waddr = io_write_bits_addr[11:3];
  assign raddr = io_read_bits_addr[11:3];
  assign T_716 = io_write_bits_way_en[0];
  assign T_717 = io_read_bits_way_en[0];
  assign T_724_0 = T_735_0_T_761_data;
  assign GEN_0 = io_read_valid ? io_read_bits_addr : T_726;
  assign T_735_0_T_761_addr = T_758;
  assign T_735_0_T_761_en = T_756;
  assign T_735_0_T_761_data = T_735_0[GEN_3];
  assign T_735_0_T_752_data = T_747_0;
  assign T_735_0_T_752_addr = waddr;
  assign T_735_0_T_752_mask = GEN_8;
  assign T_735_0_T_752_en = T_740;
  assign T_738 = T_716 & io_write_valid;
  assign T_740 = T_738 & io_write_bits_wmask;
  assign T_747_0 = io_write_bits_data;
  assign GEN_8 = T_740 ? T_716 : 1'h0;
  assign T_756 = T_717 & io_read_valid;
  assign T_758 = raddr;
  assign T_769_0 = T_724_0;
  assign T_771 = io_write_bits_way_en[1];
  assign T_772 = io_read_bits_way_en[1];
  assign T_779_0 = T_790_0_T_816_data;
  assign GEN_11 = io_read_valid ? io_read_bits_addr : T_781;
  assign T_790_0_T_816_addr = T_813;
  assign T_790_0_T_816_en = T_811;
  assign T_790_0_T_816_data = T_790_0[GEN_7];
  assign T_790_0_T_807_data = T_802_0;
  assign T_790_0_T_807_addr = waddr;
  assign T_790_0_T_807_mask = GEN_19;
  assign T_790_0_T_807_en = T_795;
  assign T_793 = T_771 & io_write_valid;
  assign T_795 = T_793 & io_write_bits_wmask;
  assign T_802_0 = io_write_bits_data;
  assign GEN_19 = T_795 ? T_771 : 1'h0;
  assign T_811 = T_772 & io_read_valid;
  assign T_813 = raddr;
  assign T_824_0 = T_779_0;
  assign T_826 = io_write_bits_way_en[2];
  assign T_827 = io_read_bits_way_en[2];
  assign T_834_0 = T_845_0_T_871_data;
  assign GEN_22 = io_read_valid ? io_read_bits_addr : T_836;
  assign T_845_0_T_871_addr = T_868;
  assign T_845_0_T_871_en = T_866;
  assign T_845_0_T_871_data = T_845_0[GEN_13];
  assign T_845_0_T_862_data = T_857_0;
  assign T_845_0_T_862_addr = waddr;
  assign T_845_0_T_862_mask = GEN_30;
  assign T_845_0_T_862_en = T_850;
  assign T_848 = T_826 & io_write_valid;
  assign T_850 = T_848 & io_write_bits_wmask;
  assign T_857_0 = io_write_bits_data;
  assign GEN_30 = T_850 ? T_826 : 1'h0;
  assign T_866 = T_827 & io_read_valid;
  assign T_868 = raddr;
  assign T_879_0 = T_834_0;
  assign T_881 = io_write_bits_way_en[3];
  assign T_882 = io_read_bits_way_en[3];
  assign T_889_0 = T_900_0_T_926_data;
  assign GEN_33 = io_read_valid ? io_read_bits_addr : T_891;
  assign T_900_0_T_926_addr = T_923;
  assign T_900_0_T_926_en = T_921;
  assign T_900_0_T_926_data = T_900_0[GEN_17];
  assign T_900_0_T_917_data = T_912_0;
  assign T_900_0_T_917_addr = waddr;
  assign T_900_0_T_917_mask = GEN_41;
  assign T_900_0_T_917_en = T_905;
  assign T_903 = T_881 & io_write_valid;
  assign T_905 = T_903 & io_write_bits_wmask;
  assign T_912_0 = io_write_bits_data;
  assign GEN_41 = T_905 ? T_881 : 1'h0;
  assign T_921 = T_882 & io_read_valid;
  assign T_923 = raddr;
  assign T_934_0 = T_889_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_726 = GEN_1[11:0];
  `endif
  GEN_2 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_735_0[initvar] = GEN_2[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_781 = GEN_5[11:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_790_0[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  GEN_7 = GEN_9[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  T_836 = GEN_10[11:0];
  `endif
  GEN_12 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_845_0[initvar] = GEN_12[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  T_891 = GEN_15[11:0];
  `endif
  GEN_16 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_900_0[initvar] = GEN_16[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_18 = {1{$random}};
  GEN_17 = GEN_18[8:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_726 <= io_read_bits_addr;
      end
    end
    if(T_735_0_T_761_en) begin
      GEN_3 <= T_735_0_T_761_addr;
    end
    if(T_735_0_T_752_en & T_735_0_T_752_mask) begin
      T_735_0[T_735_0_T_752_addr] <= T_735_0_T_752_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_781 <= io_read_bits_addr;
      end
    end
    if(T_790_0_T_816_en) begin
      GEN_7 <= T_790_0_T_816_addr;
    end
    if(T_790_0_T_807_en & T_790_0_T_807_mask) begin
      T_790_0[T_790_0_T_807_addr] <= T_790_0_T_807_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_836 <= io_read_bits_addr;
      end
    end
    if(T_845_0_T_871_en) begin
      GEN_13 <= T_845_0_T_871_addr;
    end
    if(T_845_0_T_862_en & T_845_0_T_862_mask) begin
      T_845_0[T_845_0_T_862_addr] <= T_845_0_T_862_data;
    end
    if(1'h0) begin
    end else begin
      if(io_read_valid) begin
        T_891 <= io_read_bits_addr;
      end
    end
    if(T_900_0_T_926_en) begin
      GEN_17 <= T_900_0_T_926_addr;
    end
    if(T_900_0_T_917_en & T_900_0_T_917_mask) begin
      T_900_0[T_900_0_T_917_addr] <= T_900_0_T_917_data;
    end
  end
endmodule
module Arbiter_10(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [3:0] io_in_2_bits_way_en,
  input  [11:0] io_in_2_bits_addr,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [3:0] io_in_3_bits_way_en,
  input  [11:0] io_in_3_bits_addr,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire [1:0] GEN_3;
  wire [3:0] GEN_4;
  wire [11:0] GEN_5;
  wire [1:0] GEN_6;
  wire [3:0] GEN_7;
  wire [11:0] GEN_8;
  wire  T_1934;
  wire  T_1935;
  wire  grant_1;
  wire  grant_2;
  wire  grant_3;
  wire  T_1940;
  wire  T_1941;
  wire  T_1942;
  wire  T_1944;
  wire  T_1945;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1940;
  assign io_in_2_ready = T_1941;
  assign io_in_3_ready = T_1942;
  assign io_out_valid = T_1945;
  assign io_out_bits_way_en = GEN_7;
  assign io_out_bits_addr = GEN_8;
  assign io_chosen = GEN_6;
  assign GEN_0 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_1 = io_in_2_valid ? io_in_2_bits_way_en : io_in_3_bits_way_en;
  assign GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign GEN_3 = io_in_1_valid ? 2'h1 : GEN_0;
  assign GEN_4 = io_in_1_valid ? io_in_1_bits_way_en : GEN_1;
  assign GEN_5 = io_in_1_valid ? io_in_1_bits_addr : GEN_2;
  assign GEN_6 = io_in_0_valid ? 2'h0 : GEN_3;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : GEN_4;
  assign GEN_8 = io_in_0_valid ? io_in_0_bits_addr : GEN_5;
  assign T_1934 = io_in_0_valid | io_in_1_valid;
  assign T_1935 = T_1934 | io_in_2_valid;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign grant_2 = T_1934 == 1'h0;
  assign grant_3 = T_1935 == 1'h0;
  assign T_1940 = grant_1 & io_out_ready;
  assign T_1941 = grant_2 & io_out_ready;
  assign T_1942 = grant_3 & io_out_ready;
  assign T_1944 = grant_3 == 1'h0;
  assign T_1945 = T_1944 | io_in_3_valid;
endmodule
module Arbiter_11(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  input   io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  input   io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output  io_out_bits_wmask,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire  GEN_3;
  wire [63:0] GEN_4;
  wire  grant_1;
  wire  T_1466;
  wire  T_1468;
  wire  T_1469;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1466;
  assign io_out_valid = T_1469;
  assign io_out_bits_way_en = GEN_1;
  assign io_out_bits_addr = GEN_2;
  assign io_out_bits_wmask = GEN_3;
  assign io_out_bits_data = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign grant_1 = io_in_0_valid == 1'h0;
  assign T_1466 = grant_1 & io_out_ready;
  assign T_1468 = grant_1 == 1'h0;
  assign T_1469 = T_1468 | io_in_1_valid;
endmodule
module AMOALU(
  input   clk,
  input   reset,
  input  [2:0] io_addr,
  input  [4:0] io_cmd,
  input  [1:0] io_typ,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out
);
  wire  T_8;
  wire [31:0] T_9;
  wire [63:0] T_10;
  wire [63:0] rhs;
  wire  T_11;
  wire  T_12;
  wire  sgned;
  wire  T_14;
  wire  max;
  wire  T_16;
  wire  min;
  wire  T_19;
  wire [31:0] GEN_0;
  wire [31:0] T_20;
  wire [63:0] GEN_1;
  wire [63:0] T_21;
  wire [63:0] T_22;
  wire [63:0] T_23;
  wire [64:0] T_24;
  wire [63:0] adder_out;
  wire  T_25;
  wire  T_27;
  wire  T_30;
  wire  T_31;
  wire  T_32;
  wire  T_33;
  wire  T_34;
  wire  T_39;
  wire  T_40;
  wire  T_41;
  wire [31:0] T_42;
  wire [31:0] T_43;
  wire  T_44;
  wire [31:0] T_45;
  wire [31:0] T_46;
  wire  T_47;
  wire  T_50;
  wire  T_52;
  wire  T_53;
  wire  T_54;
  wire  T_55;
  wire  T_56;
  wire  T_57;
  wire  less;
  wire  T_58;
  wire  T_59;
  wire [63:0] T_60;
  wire  T_61;
  wire [63:0] T_62;
  wire  T_63;
  wire [63:0] T_64;
  wire  T_65;
  wire  T_67;
  wire [7:0] T_68;
  wire [15:0] T_69;
  wire [31:0] T_70;
  wire [63:0] T_71;
  wire  T_73;
  wire [15:0] T_74;
  wire [31:0] T_75;
  wire [63:0] T_76;
  wire [63:0] T_82;
  wire [63:0] T_83;
  wire [63:0] T_84;
  wire [63:0] T_85;
  wire [63:0] T_86;
  wire [63:0] T_87;
  wire [63:0] out;
  wire  T_89;
  wire  T_93;
  wire  T_97;
  wire  T_100;
  wire [1:0] T_101;
  wire  T_102;
  wire [1:0] T_104;
  wire  T_106;
  wire [1:0] T_109;
  wire [1:0] T_110;
  wire [1:0] T_113;
  wire [3:0] T_114;
  wire [3:0] T_117;
  wire  T_119;
  wire [3:0] T_122;
  wire [3:0] T_123;
  wire [3:0] T_126;
  wire [7:0] T_127;
  wire  T_128;
  wire  T_129;
  wire  T_130;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire  T_134;
  wire  T_135;
  wire [7:0] T_139;
  wire [7:0] T_143;
  wire [7:0] T_147;
  wire [7:0] T_151;
  wire [7:0] T_155;
  wire [7:0] T_159;
  wire [7:0] T_163;
  wire [7:0] T_167;
  wire [15:0] T_168;
  wire [15:0] T_169;
  wire [31:0] T_170;
  wire [15:0] T_171;
  wire [15:0] T_172;
  wire [31:0] T_173;
  wire [63:0] wmask;
  wire [63:0] T_174;
  wire [63:0] T_175;
  wire [63:0] T_176;
  wire [63:0] T_177;
  assign io_out = T_177;
  assign T_8 = io_typ == 2'h2;
  assign T_9 = io_rhs[31:0];
  assign T_10 = {T_9,T_9};
  assign rhs = T_8 ? T_10 : io_rhs;
  assign T_11 = io_cmd == 5'hc;
  assign T_12 = io_cmd == 5'hd;
  assign sgned = T_11 | T_12;
  assign T_14 = io_cmd == 5'hf;
  assign max = T_12 | T_14;
  assign T_16 = io_cmd == 5'he;
  assign min = T_11 | T_16;
  assign T_19 = io_addr[2];
  assign GEN_0 = {{31'd0}, T_19};
  assign T_20 = GEN_0 << 31;
  assign GEN_1 = {{32'd0}, T_20};
  assign T_21 = 64'hffffffffffffffff ^ GEN_1;
  assign T_22 = io_lhs & T_21;
  assign T_23 = rhs & T_21;
  assign T_24 = T_22 + T_23;
  assign adder_out = T_24[63:0];
  assign T_25 = io_typ[0];
  assign T_27 = T_25 == 1'h0;
  assign T_30 = T_19 == 1'h0;
  assign T_31 = T_27 & T_30;
  assign T_32 = io_lhs[31];
  assign T_33 = io_lhs[63];
  assign T_34 = T_31 ? T_32 : T_33;
  assign T_39 = rhs[31];
  assign T_40 = rhs[63];
  assign T_41 = T_31 ? T_39 : T_40;
  assign T_42 = io_lhs[31:0];
  assign T_43 = rhs[31:0];
  assign T_44 = T_42 < T_43;
  assign T_45 = io_lhs[63:32];
  assign T_46 = rhs[63:32];
  assign T_47 = T_45 < T_46;
  assign T_50 = T_45 == T_46;
  assign T_52 = T_19 ? T_47 : T_44;
  assign T_53 = T_50 & T_44;
  assign T_54 = T_47 | T_53;
  assign T_55 = T_27 ? T_52 : T_54;
  assign T_56 = T_34 == T_41;
  assign T_57 = sgned ? T_34 : T_41;
  assign less = T_56 ? T_55 : T_57;
  assign T_58 = io_cmd == 5'h8;
  assign T_59 = io_cmd == 5'hb;
  assign T_60 = io_lhs & rhs;
  assign T_61 = io_cmd == 5'ha;
  assign T_62 = io_lhs | rhs;
  assign T_63 = io_cmd == 5'h9;
  assign T_64 = io_lhs ^ rhs;
  assign T_65 = less ? min : max;
  assign T_67 = io_typ == 2'h0;
  assign T_68 = io_rhs[7:0];
  assign T_69 = {T_68,T_68};
  assign T_70 = {T_69,T_69};
  assign T_71 = {T_70,T_70};
  assign T_73 = io_typ == 2'h1;
  assign T_74 = io_rhs[15:0];
  assign T_75 = {T_74,T_74};
  assign T_76 = {T_75,T_75};
  assign T_82 = T_73 ? T_76 : rhs;
  assign T_83 = T_67 ? T_71 : T_82;
  assign T_84 = T_65 ? io_lhs : T_83;
  assign T_85 = T_63 ? T_64 : T_84;
  assign T_86 = T_61 ? T_62 : T_85;
  assign T_87 = T_59 ? T_60 : T_86;
  assign out = T_58 ? adder_out : T_87;
  assign T_89 = io_addr[0];
  assign T_93 = io_typ >= 2'h1;
  assign T_97 = T_89 | T_93;
  assign T_100 = T_89 ? 1'h0 : 1'h1;
  assign T_101 = {T_97,T_100};
  assign T_102 = io_addr[1];
  assign T_104 = T_102 ? T_101 : 2'h0;
  assign T_106 = io_typ >= 2'h2;
  assign T_109 = T_106 ? 2'h3 : 2'h0;
  assign T_110 = T_104 | T_109;
  assign T_113 = T_102 ? 2'h0 : T_101;
  assign T_114 = {T_110,T_113};
  assign T_117 = T_19 ? T_114 : 4'h0;
  assign T_119 = io_typ >= 2'h3;
  assign T_122 = T_119 ? 4'hf : 4'h0;
  assign T_123 = T_117 | T_122;
  assign T_126 = T_19 ? 4'h0 : T_114;
  assign T_127 = {T_123,T_126};
  assign T_128 = T_127[0];
  assign T_129 = T_127[1];
  assign T_130 = T_127[2];
  assign T_131 = T_127[3];
  assign T_132 = T_127[4];
  assign T_133 = T_127[5];
  assign T_134 = T_127[6];
  assign T_135 = T_127[7];
  assign T_139 = T_128 ? 8'hff : 8'h0;
  assign T_143 = T_129 ? 8'hff : 8'h0;
  assign T_147 = T_130 ? 8'hff : 8'h0;
  assign T_151 = T_131 ? 8'hff : 8'h0;
  assign T_155 = T_132 ? 8'hff : 8'h0;
  assign T_159 = T_133 ? 8'hff : 8'h0;
  assign T_163 = T_134 ? 8'hff : 8'h0;
  assign T_167 = T_135 ? 8'hff : 8'h0;
  assign T_168 = {T_143,T_139};
  assign T_169 = {T_151,T_147};
  assign T_170 = {T_169,T_168};
  assign T_171 = {T_159,T_155};
  assign T_172 = {T_167,T_163};
  assign T_173 = {T_172,T_171};
  assign wmask = {T_173,T_170};
  assign T_174 = wmask & out;
  assign T_175 = ~ wmask;
  assign T_176 = T_175 & io_lhs;
  assign T_177 = T_174 | T_176;
endmodule
module LockingArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_voluntary;
  wire [2:0] GEN_0_bits_r_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [25:0] GEN_10;
  wire [1:0] GEN_11;
  wire  GEN_12;
  wire [2:0] GEN_13;
  wire [63:0] GEN_14;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_voluntary;
  wire [2:0] GEN_1_bits_r_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_voluntary;
  wire [2:0] GEN_2_bits_r_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_voluntary;
  wire [2:0] GEN_3_bits_r_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [25:0] GEN_4_bits_addr_block;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_voluntary;
  wire [2:0] GEN_4_bits_r_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [25:0] GEN_5_bits_addr_block;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_voluntary;
  wire [2:0] GEN_5_bits_r_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [25:0] GEN_6_bits_addr_block;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_voluntary;
  wire [2:0] GEN_6_bits_r_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_740;
  reg [31:0] GEN_0;
  reg  T_742;
  reg [31:0] GEN_1;
  wire  T_744;
  wire  T_746;
  wire  T_747;
  wire  T_748;
  wire  T_749;
  wire  T_750;
  wire  T_752;
  wire  T_753;
  wire [3:0] T_757;
  wire [2:0] T_758;
  wire  GEN_63;
  wire [2:0] GEN_64;
  wire  GEN_65;
  wire  T_761;
  wire  T_763;
  wire  T_764;
  wire  T_765;
  wire  T_768;
  wire  T_769;
  wire  GEN_66;
  assign io_in_0_ready = T_765;
  assign io_in_1_ready = T_769;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_addr_block = GEN_2_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_3_bits_client_xact_id;
  assign io_out_bits_voluntary = GEN_4_bits_voluntary;
  assign io_out_bits_r_type = GEN_5_bits_r_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_65;
  assign choice = GEN_66;
  assign GEN_0_ready = GEN_7;
  assign GEN_0_valid = GEN_8;
  assign GEN_0_bits_addr_beat = GEN_9;
  assign GEN_0_bits_addr_block = GEN_10;
  assign GEN_0_bits_client_xact_id = GEN_11;
  assign GEN_0_bits_voluntary = GEN_12;
  assign GEN_0_bits_r_type = GEN_13;
  assign GEN_0_bits_data = GEN_14;
  assign GEN_7 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_10 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_13 = io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_14 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_1_ready = GEN_7;
  assign GEN_1_valid = GEN_8;
  assign GEN_1_bits_addr_beat = GEN_9;
  assign GEN_1_bits_addr_block = GEN_10;
  assign GEN_1_bits_client_xact_id = GEN_11;
  assign GEN_1_bits_voluntary = GEN_12;
  assign GEN_1_bits_r_type = GEN_13;
  assign GEN_1_bits_data = GEN_14;
  assign GEN_2_ready = GEN_7;
  assign GEN_2_valid = GEN_8;
  assign GEN_2_bits_addr_beat = GEN_9;
  assign GEN_2_bits_addr_block = GEN_10;
  assign GEN_2_bits_client_xact_id = GEN_11;
  assign GEN_2_bits_voluntary = GEN_12;
  assign GEN_2_bits_r_type = GEN_13;
  assign GEN_2_bits_data = GEN_14;
  assign GEN_3_ready = GEN_7;
  assign GEN_3_valid = GEN_8;
  assign GEN_3_bits_addr_beat = GEN_9;
  assign GEN_3_bits_addr_block = GEN_10;
  assign GEN_3_bits_client_xact_id = GEN_11;
  assign GEN_3_bits_voluntary = GEN_12;
  assign GEN_3_bits_r_type = GEN_13;
  assign GEN_3_bits_data = GEN_14;
  assign GEN_4_ready = GEN_7;
  assign GEN_4_valid = GEN_8;
  assign GEN_4_bits_addr_beat = GEN_9;
  assign GEN_4_bits_addr_block = GEN_10;
  assign GEN_4_bits_client_xact_id = GEN_11;
  assign GEN_4_bits_voluntary = GEN_12;
  assign GEN_4_bits_r_type = GEN_13;
  assign GEN_4_bits_data = GEN_14;
  assign GEN_5_ready = GEN_7;
  assign GEN_5_valid = GEN_8;
  assign GEN_5_bits_addr_beat = GEN_9;
  assign GEN_5_bits_addr_block = GEN_10;
  assign GEN_5_bits_client_xact_id = GEN_11;
  assign GEN_5_bits_voluntary = GEN_12;
  assign GEN_5_bits_r_type = GEN_13;
  assign GEN_5_bits_data = GEN_14;
  assign GEN_6_ready = GEN_7;
  assign GEN_6_valid = GEN_8;
  assign GEN_6_bits_addr_beat = GEN_9;
  assign GEN_6_bits_addr_block = GEN_10;
  assign GEN_6_bits_client_xact_id = GEN_11;
  assign GEN_6_bits_voluntary = GEN_12;
  assign GEN_6_bits_r_type = GEN_13;
  assign GEN_6_bits_data = GEN_14;
  assign T_744 = T_740 != 3'h0;
  assign T_746 = io_out_bits_r_type == 3'h0;
  assign T_747 = io_out_bits_r_type == 3'h1;
  assign T_748 = io_out_bits_r_type == 3'h2;
  assign T_749 = T_746 | T_747;
  assign T_750 = T_749 | T_748;
  assign T_752 = io_out_ready & io_out_valid;
  assign T_753 = T_752 & T_750;
  assign T_757 = T_740 + 3'h1;
  assign T_758 = T_757[2:0];
  assign GEN_63 = T_753 ? io_chosen : T_742;
  assign GEN_64 = T_753 ? T_758 : T_740;
  assign GEN_65 = T_744 ? T_742 : choice;
  assign T_761 = io_in_0_valid == 1'h0;
  assign T_763 = T_742 == 1'h0;
  assign T_764 = T_744 ? T_763 : 1'h1;
  assign T_765 = T_764 & io_out_ready;
  assign T_768 = T_744 ? T_742 : T_761;
  assign T_769 = T_768 & io_out_ready;
  assign GEN_66 = io_in_0_valid ? 1'h0 : 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_740 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_742 = GEN_1[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_740 <= 3'h0;
    end else begin
      if(T_753) begin
        T_740 <= T_758;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_753) begin
        T_742 <= io_chosen;
      end
    end
  end
endmodule
module FlowThroughSerializer_1(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_in_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_manager_id,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_manager_id = io_in_bits_manager_id;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module HellaCache(
  input   clk,
  input   reset,
  output  io_cpu_req_ready,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [6:0] io_cpu_req_bits_tag,
  input  [4:0] io_cpu_req_bits_cmd,
  input  [2:0] io_cpu_req_bits_typ,
  input   io_cpu_req_bits_phys,
  input  [63:0] io_cpu_req_bits_data,
  input   io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data,
  output  io_cpu_s2_nack,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_addr,
  output [6:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [2:0] io_cpu_resp_bits_typ,
  output [63:0] io_cpu_resp_bits_data,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_store_data,
  output  io_cpu_replay_next,
  output  io_cpu_xcpt_ma_ld,
  output  io_cpu_xcpt_ma_st,
  output  io_cpu_xcpt_pf_ld,
  output  io_cpu_xcpt_pf_st,
  input   io_cpu_invalidate_lr,
  output  io_cpu_ordered,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [26:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [37:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [10:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_probe_ready,
  input   io_mem_probe_valid,
  input  [25:0] io_mem_probe_bits_addr_block,
  input  [1:0] io_mem_probe_bits_p_type,
  input   io_mem_release_ready,
  output  io_mem_release_valid,
  output [2:0] io_mem_release_bits_addr_beat,
  output [25:0] io_mem_release_bits_addr_block,
  output [1:0] io_mem_release_bits_client_xact_id,
  output  io_mem_release_bits_voluntary,
  output [2:0] io_mem_release_bits_r_type,
  output [63:0] io_mem_release_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id
);
  wire  wb_clk;
  wire  wb_reset;
  wire  wb_io_req_ready;
  wire  wb_io_req_valid;
  wire [2:0] wb_io_req_bits_addr_beat;
  wire [25:0] wb_io_req_bits_addr_block;
  wire [1:0] wb_io_req_bits_client_xact_id;
  wire  wb_io_req_bits_voluntary;
  wire [2:0] wb_io_req_bits_r_type;
  wire [63:0] wb_io_req_bits_data;
  wire [3:0] wb_io_req_bits_way_en;
  wire  wb_io_meta_read_ready;
  wire  wb_io_meta_read_valid;
  wire [5:0] wb_io_meta_read_bits_idx;
  wire [3:0] wb_io_meta_read_bits_way_en;
  wire [19:0] wb_io_meta_read_bits_tag;
  wire  wb_io_data_req_ready;
  wire  wb_io_data_req_valid;
  wire [3:0] wb_io_data_req_bits_way_en;
  wire [11:0] wb_io_data_req_bits_addr;
  wire [63:0] wb_io_data_resp;
  wire  wb_io_release_ready;
  wire  wb_io_release_valid;
  wire [2:0] wb_io_release_bits_addr_beat;
  wire [25:0] wb_io_release_bits_addr_block;
  wire [1:0] wb_io_release_bits_client_xact_id;
  wire  wb_io_release_bits_voluntary;
  wire [2:0] wb_io_release_bits_r_type;
  wire [63:0] wb_io_release_bits_data;
  wire  prober_clk;
  wire  prober_reset;
  wire  prober_io_req_ready;
  wire  prober_io_req_valid;
  wire [25:0] prober_io_req_bits_addr_block;
  wire [1:0] prober_io_req_bits_p_type;
  wire [1:0] prober_io_req_bits_client_xact_id;
  wire  prober_io_rep_ready;
  wire  prober_io_rep_valid;
  wire [2:0] prober_io_rep_bits_addr_beat;
  wire [25:0] prober_io_rep_bits_addr_block;
  wire [1:0] prober_io_rep_bits_client_xact_id;
  wire  prober_io_rep_bits_voluntary;
  wire [2:0] prober_io_rep_bits_r_type;
  wire [63:0] prober_io_rep_bits_data;
  wire  prober_io_meta_read_ready;
  wire  prober_io_meta_read_valid;
  wire [5:0] prober_io_meta_read_bits_idx;
  wire [3:0] prober_io_meta_read_bits_way_en;
  wire [19:0] prober_io_meta_read_bits_tag;
  wire  prober_io_meta_write_ready;
  wire  prober_io_meta_write_valid;
  wire [5:0] prober_io_meta_write_bits_idx;
  wire [3:0] prober_io_meta_write_bits_way_en;
  wire [19:0] prober_io_meta_write_bits_data_tag;
  wire [1:0] prober_io_meta_write_bits_data_coh_state;
  wire  prober_io_wb_req_ready;
  wire  prober_io_wb_req_valid;
  wire [2:0] prober_io_wb_req_bits_addr_beat;
  wire [25:0] prober_io_wb_req_bits_addr_block;
  wire [1:0] prober_io_wb_req_bits_client_xact_id;
  wire  prober_io_wb_req_bits_voluntary;
  wire [2:0] prober_io_wb_req_bits_r_type;
  wire [63:0] prober_io_wb_req_bits_data;
  wire [3:0] prober_io_wb_req_bits_way_en;
  wire [3:0] prober_io_way_en;
  wire  prober_io_mshr_rdy;
  wire [1:0] prober_io_block_state_state;
  wire  mshrs_clk;
  wire  mshrs_reset;
  wire  mshrs_io_req_ready;
  wire  mshrs_io_req_valid;
  wire [39:0] mshrs_io_req_bits_addr;
  wire [6:0] mshrs_io_req_bits_tag;
  wire [4:0] mshrs_io_req_bits_cmd;
  wire [2:0] mshrs_io_req_bits_typ;
  wire  mshrs_io_req_bits_phys;
  wire [63:0] mshrs_io_req_bits_data;
  wire  mshrs_io_req_bits_tag_match;
  wire [19:0] mshrs_io_req_bits_old_meta_tag;
  wire [1:0] mshrs_io_req_bits_old_meta_coh_state;
  wire [3:0] mshrs_io_req_bits_way_en;
  wire  mshrs_io_resp_ready;
  wire  mshrs_io_resp_valid;
  wire [39:0] mshrs_io_resp_bits_addr;
  wire [6:0] mshrs_io_resp_bits_tag;
  wire [4:0] mshrs_io_resp_bits_cmd;
  wire [2:0] mshrs_io_resp_bits_typ;
  wire [63:0] mshrs_io_resp_bits_data;
  wire  mshrs_io_resp_bits_replay;
  wire  mshrs_io_resp_bits_has_data;
  wire [63:0] mshrs_io_resp_bits_data_word_bypass;
  wire [63:0] mshrs_io_resp_bits_store_data;
  wire  mshrs_io_secondary_miss;
  wire  mshrs_io_mem_req_ready;
  wire  mshrs_io_mem_req_valid;
  wire [25:0] mshrs_io_mem_req_bits_addr_block;
  wire [1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_req_bits_addr_beat;
  wire  mshrs_io_mem_req_bits_is_builtin_type;
  wire [2:0] mshrs_io_mem_req_bits_a_type;
  wire [10:0] mshrs_io_mem_req_bits_union;
  wire [63:0] mshrs_io_mem_req_bits_data;
  wire [3:0] mshrs_io_refill_way_en;
  wire [11:0] mshrs_io_refill_addr;
  wire  mshrs_io_meta_read_ready;
  wire  mshrs_io_meta_read_valid;
  wire [5:0] mshrs_io_meta_read_bits_idx;
  wire [3:0] mshrs_io_meta_read_bits_way_en;
  wire [19:0] mshrs_io_meta_read_bits_tag;
  wire  mshrs_io_meta_write_ready;
  wire  mshrs_io_meta_write_valid;
  wire [5:0] mshrs_io_meta_write_bits_idx;
  wire [3:0] mshrs_io_meta_write_bits_way_en;
  wire [19:0] mshrs_io_meta_write_bits_data_tag;
  wire [1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire  mshrs_io_replay_ready;
  wire  mshrs_io_replay_valid;
  wire [39:0] mshrs_io_replay_bits_addr;
  wire [6:0] mshrs_io_replay_bits_tag;
  wire [4:0] mshrs_io_replay_bits_cmd;
  wire [2:0] mshrs_io_replay_bits_typ;
  wire  mshrs_io_replay_bits_phys;
  wire [63:0] mshrs_io_replay_bits_data;
  wire  mshrs_io_mem_grant_valid;
  wire [2:0] mshrs_io_mem_grant_bits_addr_beat;
  wire [1:0] mshrs_io_mem_grant_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_grant_bits_manager_xact_id;
  wire  mshrs_io_mem_grant_bits_is_builtin_type;
  wire [3:0] mshrs_io_mem_grant_bits_g_type;
  wire [63:0] mshrs_io_mem_grant_bits_data;
  wire  mshrs_io_mem_grant_bits_manager_id;
  wire  mshrs_io_mem_finish_ready;
  wire  mshrs_io_mem_finish_valid;
  wire [2:0] mshrs_io_mem_finish_bits_manager_xact_id;
  wire  mshrs_io_mem_finish_bits_manager_id;
  wire  mshrs_io_wb_req_ready;
  wire  mshrs_io_wb_req_valid;
  wire [2:0] mshrs_io_wb_req_bits_addr_beat;
  wire [25:0] mshrs_io_wb_req_bits_addr_block;
  wire [1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire  mshrs_io_wb_req_bits_voluntary;
  wire [2:0] mshrs_io_wb_req_bits_r_type;
  wire [63:0] mshrs_io_wb_req_bits_data;
  wire [3:0] mshrs_io_wb_req_bits_way_en;
  wire  mshrs_io_probe_rdy;
  wire  mshrs_io_fence_rdy;
  wire  mshrs_io_replay_next;
  wire  T_1901;
  reg  s1_valid;
  reg [31:0] GEN_94;
  reg [39:0] s1_req_addr;
  reg [63:0] GEN_95;
  reg [6:0] s1_req_tag;
  reg [31:0] GEN_96;
  reg [4:0] s1_req_cmd;
  reg [31:0] GEN_97;
  reg [2:0] s1_req_typ;
  reg [31:0] GEN_98;
  reg  s1_req_phys;
  reg [31:0] GEN_99;
  reg [63:0] s1_req_data;
  reg [63:0] GEN_100;
  wire  T_1970;
  wire  T_1971;
  wire [1:0] T_1972;
  wire [1:0] T_1973;
  wire [3:0] T_1974;
  wire  T_1976;
  wire  T_1978;
  wire  s1_valid_masked;
  reg  s1_replay;
  reg [31:0] GEN_101;
  reg  s1_clk_en;
  reg [31:0] GEN_102;
  reg  s2_valid;
  reg [31:0] GEN_103;
  reg [39:0] s2_req_addr;
  reg [63:0] GEN_104;
  reg [6:0] s2_req_tag;
  reg [31:0] GEN_105;
  reg [4:0] s2_req_cmd;
  reg [31:0] GEN_106;
  reg [2:0] s2_req_typ;
  reg [31:0] GEN_107;
  reg  s2_req_phys;
  reg [31:0] GEN_108;
  reg [63:0] s2_req_data;
  reg [63:0] GEN_109;
  reg  T_2049;
  reg [31:0] GEN_110;
  wire  T_2050;
  wire  s2_replay;
  wire  s2_recycle;
  wire  s2_valid_masked;
  reg  s3_valid;
  reg [31:0] GEN_111;
  reg [39:0] s3_req_addr;
  reg [63:0] GEN_112;
  reg [6:0] s3_req_tag;
  reg [31:0] GEN_113;
  reg [4:0] s3_req_cmd;
  reg [31:0] GEN_114;
  reg [2:0] s3_req_typ;
  reg [31:0] GEN_115;
  reg  s3_req_phys;
  reg [31:0] GEN_116;
  reg [63:0] s3_req_data;
  reg [63:0] GEN_117;
  reg [3:0] s3_way;
  reg [31:0] GEN_118;
  reg  s1_recycled;
  reg [31:0] GEN_119;
  wire  GEN_0;
  wire  T_2122;
  wire  T_2123;
  wire  T_2124;
  wire  T_2125;
  wire  T_2126;
  wire  T_2127;
  wire  T_2128;
  wire  T_2129;
  wire  s1_read;
  wire  T_2130;
  wire  T_2132;
  wire  s1_write;
  wire  T_2136;
  wire  T_2137;
  wire  T_2138;
  wire  T_2139;
  wire  s1_readwrite;
  wire  dtlb_clk;
  wire  dtlb_reset;
  wire  dtlb_io_req_ready;
  wire  dtlb_io_req_valid;
  wire [27:0] dtlb_io_req_bits_vpn;
  wire  dtlb_io_req_bits_passthrough;
  wire  dtlb_io_req_bits_instruction;
  wire  dtlb_io_req_bits_store;
  wire  dtlb_io_resp_miss;
  wire [19:0] dtlb_io_resp_ppn;
  wire  dtlb_io_resp_xcpt_ld;
  wire  dtlb_io_resp_xcpt_st;
  wire  dtlb_io_resp_xcpt_if;
  wire  dtlb_io_resp_cacheable;
  wire  dtlb_io_ptw_req_ready;
  wire  dtlb_io_ptw_req_valid;
  wire [1:0] dtlb_io_ptw_req_bits_prv;
  wire  dtlb_io_ptw_req_bits_pum;
  wire  dtlb_io_ptw_req_bits_mxr;
  wire [26:0] dtlb_io_ptw_req_bits_addr;
  wire  dtlb_io_ptw_req_bits_store;
  wire  dtlb_io_ptw_req_bits_fetch;
  wire  dtlb_io_ptw_resp_valid;
  wire [15:0] dtlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] dtlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] dtlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  dtlb_io_ptw_resp_bits_pte_d;
  wire  dtlb_io_ptw_resp_bits_pte_a;
  wire  dtlb_io_ptw_resp_bits_pte_g;
  wire  dtlb_io_ptw_resp_bits_pte_u;
  wire  dtlb_io_ptw_resp_bits_pte_x;
  wire  dtlb_io_ptw_resp_bits_pte_w;
  wire  dtlb_io_ptw_resp_bits_pte_r;
  wire  dtlb_io_ptw_resp_bits_pte_v;
  wire [6:0] dtlb_io_ptw_ptbr_asid;
  wire [37:0] dtlb_io_ptw_ptbr_ppn;
  wire  dtlb_io_ptw_invalidate;
  wire  dtlb_io_ptw_status_debug;
  wire [1:0] dtlb_io_ptw_status_prv;
  wire  dtlb_io_ptw_status_sd;
  wire [30:0] dtlb_io_ptw_status_zero3;
  wire  dtlb_io_ptw_status_sd_rv32;
  wire [1:0] dtlb_io_ptw_status_zero2;
  wire [4:0] dtlb_io_ptw_status_vm;
  wire [3:0] dtlb_io_ptw_status_zero1;
  wire  dtlb_io_ptw_status_mxr;
  wire  dtlb_io_ptw_status_pum;
  wire  dtlb_io_ptw_status_mprv;
  wire [1:0] dtlb_io_ptw_status_xs;
  wire [1:0] dtlb_io_ptw_status_fs;
  wire [1:0] dtlb_io_ptw_status_mpp;
  wire [1:0] dtlb_io_ptw_status_hpp;
  wire  dtlb_io_ptw_status_spp;
  wire  dtlb_io_ptw_status_mpie;
  wire  dtlb_io_ptw_status_hpie;
  wire  dtlb_io_ptw_status_spie;
  wire  dtlb_io_ptw_status_upie;
  wire  dtlb_io_ptw_status_mie;
  wire  dtlb_io_ptw_status_hie;
  wire  dtlb_io_ptw_status_sie;
  wire  dtlb_io_ptw_status_uie;
  wire  T_2140;
  wire [27:0] T_2141;
  wire  T_2144;
  wire  T_2146;
  wire  T_2147;
  wire  GEN_1;
  wire [39:0] GEN_2;
  wire [6:0] GEN_3;
  wire [4:0] GEN_4;
  wire [2:0] GEN_5;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire [25:0] T_2149;
  wire [31:0] GEN_83;
  wire [31:0] T_2150;
  wire [39:0] GEN_8;
  wire  GEN_9;
  wire [25:0] T_2152;
  wire [31:0] GEN_84;
  wire [31:0] T_2153;
  wire [39:0] GEN_10;
  wire  GEN_11;
  wire [39:0] GEN_12;
  wire [6:0] GEN_13;
  wire [4:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire [63:0] GEN_17;
  wire [39:0] GEN_18;
  wire [6:0] GEN_19;
  wire [4:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [63:0] GEN_23;
  wire [11:0] T_2155;
  wire [31:0] s1_addr;
  wire [63:0] T_2156;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_27;
  wire [39:0] GEN_28;
  wire [63:0] GEN_29;
  wire [6:0] GEN_30;
  wire [4:0] GEN_31;
  wire [1:0] T_2158;
  wire [3:0] T_2160;
  wire [4:0] T_2162;
  wire [3:0] T_2163;
  wire [2:0] T_2164;
  wire [39:0] GEN_85;
  wire [39:0] T_2165;
  wire  misaligned;
  wire  T_2167;
  wire  T_2168;
  wire  T_2169;
  wire  T_2170;
  wire  meta_clk;
  wire  meta_reset;
  wire  meta_io_read_ready;
  wire  meta_io_read_valid;
  wire [5:0] meta_io_read_bits_idx;
  wire [3:0] meta_io_read_bits_way_en;
  wire  meta_io_write_ready;
  wire  meta_io_write_valid;
  wire [5:0] meta_io_write_bits_idx;
  wire [3:0] meta_io_write_bits_way_en;
  wire [19:0] meta_io_write_bits_data_tag;
  wire [1:0] meta_io_write_bits_data_coh_state;
  wire [19:0] meta_io_resp_0_tag;
  wire [1:0] meta_io_resp_0_coh_state;
  wire [19:0] meta_io_resp_1_tag;
  wire [1:0] meta_io_resp_1_coh_state;
  wire [19:0] meta_io_resp_2_tag;
  wire [1:0] meta_io_resp_2_coh_state;
  wire [19:0] meta_io_resp_3_tag;
  wire [1:0] meta_io_resp_3_coh_state;
  wire  metaReadArb_clk;
  wire  metaReadArb_reset;
  wire  metaReadArb_io_in_0_ready;
  wire  metaReadArb_io_in_0_valid;
  wire [5:0] metaReadArb_io_in_0_bits_idx;
  wire [3:0] metaReadArb_io_in_0_bits_way_en;
  wire  metaReadArb_io_in_1_ready;
  wire  metaReadArb_io_in_1_valid;
  wire [5:0] metaReadArb_io_in_1_bits_idx;
  wire [3:0] metaReadArb_io_in_1_bits_way_en;
  wire  metaReadArb_io_in_2_ready;
  wire  metaReadArb_io_in_2_valid;
  wire [5:0] metaReadArb_io_in_2_bits_idx;
  wire [3:0] metaReadArb_io_in_2_bits_way_en;
  wire  metaReadArb_io_in_3_ready;
  wire  metaReadArb_io_in_3_valid;
  wire [5:0] metaReadArb_io_in_3_bits_idx;
  wire [3:0] metaReadArb_io_in_3_bits_way_en;
  wire  metaReadArb_io_in_4_ready;
  wire  metaReadArb_io_in_4_valid;
  wire [5:0] metaReadArb_io_in_4_bits_idx;
  wire [3:0] metaReadArb_io_in_4_bits_way_en;
  wire  metaReadArb_io_out_ready;
  wire  metaReadArb_io_out_valid;
  wire [5:0] metaReadArb_io_out_bits_idx;
  wire [3:0] metaReadArb_io_out_bits_way_en;
  wire [2:0] metaReadArb_io_chosen;
  wire  metaWriteArb_clk;
  wire  metaWriteArb_reset;
  wire  metaWriteArb_io_in_0_ready;
  wire  metaWriteArb_io_in_0_valid;
  wire [5:0] metaWriteArb_io_in_0_bits_idx;
  wire [3:0] metaWriteArb_io_in_0_bits_way_en;
  wire [19:0] metaWriteArb_io_in_0_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_0_bits_data_coh_state;
  wire  metaWriteArb_io_in_1_ready;
  wire  metaWriteArb_io_in_1_valid;
  wire [5:0] metaWriteArb_io_in_1_bits_idx;
  wire [3:0] metaWriteArb_io_in_1_bits_way_en;
  wire [19:0] metaWriteArb_io_in_1_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_1_bits_data_coh_state;
  wire  metaWriteArb_io_out_ready;
  wire  metaWriteArb_io_out_valid;
  wire [5:0] metaWriteArb_io_out_bits_idx;
  wire [3:0] metaWriteArb_io_out_bits_way_en;
  wire [19:0] metaWriteArb_io_out_bits_data_tag;
  wire [1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire  metaWriteArb_io_chosen;
  wire  data_clk;
  wire  data_reset;
  wire  data_io_read_ready;
  wire  data_io_read_valid;
  wire [3:0] data_io_read_bits_way_en;
  wire [11:0] data_io_read_bits_addr;
  wire  data_io_write_ready;
  wire  data_io_write_valid;
  wire [3:0] data_io_write_bits_way_en;
  wire [11:0] data_io_write_bits_addr;
  wire  data_io_write_bits_wmask;
  wire [63:0] data_io_write_bits_data;
  wire [63:0] data_io_resp_0;
  wire [63:0] data_io_resp_1;
  wire [63:0] data_io_resp_2;
  wire [63:0] data_io_resp_3;
  wire  readArb_clk;
  wire  readArb_reset;
  wire  readArb_io_in_0_ready;
  wire  readArb_io_in_0_valid;
  wire [3:0] readArb_io_in_0_bits_way_en;
  wire [11:0] readArb_io_in_0_bits_addr;
  wire  readArb_io_in_1_ready;
  wire  readArb_io_in_1_valid;
  wire [3:0] readArb_io_in_1_bits_way_en;
  wire [11:0] readArb_io_in_1_bits_addr;
  wire  readArb_io_in_2_ready;
  wire  readArb_io_in_2_valid;
  wire [3:0] readArb_io_in_2_bits_way_en;
  wire [11:0] readArb_io_in_2_bits_addr;
  wire  readArb_io_in_3_ready;
  wire  readArb_io_in_3_valid;
  wire [3:0] readArb_io_in_3_bits_way_en;
  wire [11:0] readArb_io_in_3_bits_addr;
  wire  readArb_io_out_ready;
  wire  readArb_io_out_valid;
  wire [3:0] readArb_io_out_bits_way_en;
  wire [11:0] readArb_io_out_bits_addr;
  wire [1:0] readArb_io_chosen;
  wire  writeArb_clk;
  wire  writeArb_reset;
  wire  writeArb_io_in_0_ready;
  wire  writeArb_io_in_0_valid;
  wire [3:0] writeArb_io_in_0_bits_way_en;
  wire [11:0] writeArb_io_in_0_bits_addr;
  wire  writeArb_io_in_0_bits_wmask;
  wire [63:0] writeArb_io_in_0_bits_data;
  wire  writeArb_io_in_1_ready;
  wire  writeArb_io_in_1_valid;
  wire [3:0] writeArb_io_in_1_bits_way_en;
  wire [11:0] writeArb_io_in_1_bits_addr;
  wire  writeArb_io_in_1_bits_wmask;
  wire [63:0] writeArb_io_in_1_bits_data;
  wire  writeArb_io_out_ready;
  wire  writeArb_io_out_valid;
  wire [3:0] writeArb_io_out_bits_way_en;
  wire [11:0] writeArb_io_out_bits_addr;
  wire  writeArb_io_out_bits_wmask;
  wire [63:0] writeArb_io_out_bits_data;
  wire  writeArb_io_chosen;
  wire [63:0] wdata_encoded_0;
  wire [33:0] T_2513;
  wire  T_2515;
  wire  GEN_32;
  wire  T_2520;
  wire  GEN_33;
  wire [33:0] T_2522;
  wire [19:0] T_2525;
  wire  T_2526;
  wire  T_2528;
  wire  T_2530;
  wire  T_2532;
  wire  T_2538_0;
  wire  T_2538_1;
  wire  T_2538_2;
  wire  T_2538_3;
  wire [1:0] T_2540;
  wire [1:0] T_2541;
  wire [3:0] s1_tag_eq_way;
  wire  T_2542;
  wire  T_2543;
  wire  T_2544;
  wire  T_2545;
  wire  T_2546;
  wire  T_2547;
  wire  T_2548;
  wire  T_2549;
  wire  T_2550;
  wire  T_2551;
  wire  T_2552;
  wire  T_2553;
  wire  T_2559_0;
  wire  T_2559_1;
  wire  T_2559_2;
  wire  T_2559_3;
  wire [1:0] T_2561;
  wire [1:0] T_2562;
  wire [3:0] s1_tag_match_way;
  wire  T_2564;
  reg [3:0] s2_tag_match_way;
  reg [31:0] GEN_120;
  wire [3:0] GEN_34;
  wire  s2_tag_match;
  reg [1:0] T_2569_state;
  reg [31:0] GEN_121;
  wire [1:0] GEN_35;
  reg [1:0] T_2591_state;
  reg [31:0] GEN_122;
  wire [1:0] GEN_36;
  reg [1:0] T_2613_state;
  reg [31:0] GEN_123;
  wire [1:0] GEN_37;
  reg [1:0] T_2635_state;
  reg [31:0] GEN_124;
  wire [1:0] GEN_38;
  wire [1:0] T_2830_0_state;
  wire [1:0] T_2830_1_state;
  wire [1:0] T_2830_2_state;
  wire [1:0] T_2830_3_state;
  wire  T_2937;
  wire  T_2938;
  wire  T_2939;
  wire  T_2940;
  wire [1:0] T_2942;
  wire [1:0] T_2944;
  wire [1:0] T_2946;
  wire [1:0] T_2948;
  wire [1:0] T_2971;
  wire [1:0] T_2972;
  wire [1:0] T_2973;
  wire [1:0] s2_hit_state_state;
  wire  T_3018;
  wire  T_3019;
  wire  T_3020;
  wire  T_3021;
  wire  T_3022;
  wire  T_3023;
  wire  T_3024;
  wire  T_3025;
  wire  T_3026;
  wire  T_3027;
  wire  T_3028;
  wire  T_3029;
  wire  T_3030;
  wire  T_3031;
  wire  T_3035;
  wire  T_3036;
  wire [1:0] T_3044;
  wire [1:0] T_3067_state;
  wire  T_3089;
  wire  s2_hit;
  reg [4:0] lrsc_count;
  reg [31:0] GEN_125;
  wire  lrsc_valid;
  reg [33:0] lrsc_addr;
  reg [63:0] GEN_126;
  wire  T_3094;
  wire  s2_lrsc_addr_match;
  wire  T_3096;
  wire  s2_sc_fail;
  wire [5:0] T_3098;
  wire [4:0] T_3099;
  wire [4:0] GEN_39;
  wire  T_3100;
  wire  T_3101;
  wire  T_3103;
  wire [4:0] GEN_40;
  wire [4:0] GEN_41;
  wire [33:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [33:0] GEN_45;
  wire [4:0] GEN_46;
  wire [63:0] s2_data_0;
  wire [63:0] s2_data_1;
  wire [63:0] s2_data_2;
  wire [63:0] s2_data_3;
  reg [63:0] T_3121_0;
  reg [63:0] GEN_127;
  wire  T_3124;
  wire [63:0] T_3132;
  wire [63:0] GEN_47;
  reg [63:0] T_3139_0;
  reg [63:0] GEN_128;
  wire  T_3142;
  wire [63:0] T_3150;
  wire [63:0] GEN_48;
  reg [63:0] T_3157_0;
  reg [63:0] GEN_129;
  wire  T_3160;
  wire [63:0] T_3168;
  wire [63:0] GEN_49;
  reg [63:0] T_3175_0;
  reg [63:0] GEN_130;
  wire  T_3178;
  wire [63:0] T_3186;
  wire [63:0] GEN_50;
  wire [63:0] T_3192;
  wire [63:0] T_3194;
  wire [63:0] T_3196;
  wire [63:0] T_3198;
  wire [63:0] T_3200;
  wire [63:0] T_3201;
  wire [63:0] T_3202;
  wire [63:0] s2_data_muxed;
  wire  T_3204;
  wire  T_3208;
  wire  T_3209;
  wire  T_3217;
  wire  amoalu_clk;
  wire  amoalu_reset;
  wire [2:0] amoalu_io_addr;
  wire [4:0] amoalu_io_cmd;
  wire [1:0] amoalu_io_typ;
  wire [63:0] amoalu_io_lhs;
  wire [63:0] amoalu_io_rhs;
  wire [63:0] amoalu_io_out;
  wire  T_3218;
  wire  T_3226;
  wire  T_3227;
  wire [63:0] T_3228;
  wire [39:0] GEN_51;
  wire [6:0] GEN_52;
  wire [4:0] GEN_53;
  wire [2:0] GEN_54;
  wire  GEN_55;
  wire [63:0] GEN_56;
  wire [3:0] GEN_57;
  wire [1:0] T_3231;
  wire  T_3233;
  reg [15:0] T_3236;
  reg [31:0] GEN_131;
  wire  T_3237;
  wire  T_3238;
  wire  T_3239;
  wire  T_3240;
  wire  T_3241;
  wire  T_3242;
  wire  T_3243;
  wire [14:0] T_3244;
  wire [15:0] T_3245;
  wire [15:0] GEN_58;
  wire [1:0] T_3246;
  wire [3:0] s1_replaced_way_en;
  reg [1:0] T_3249;
  reg [31:0] GEN_132;
  wire [1:0] GEN_59;
  wire [3:0] s2_replaced_way_en;
  wire  T_3251;
  wire  T_3252;
  reg [19:0] T_3253_tag;
  reg [31:0] GEN_133;
  reg [1:0] T_3253_coh_state;
  reg [31:0] GEN_134;
  wire [19:0] GEN_60;
  wire [1:0] GEN_61;
  wire  T_3337;
  wire  T_3338;
  reg [19:0] T_3339_tag;
  reg [31:0] GEN_135;
  reg [1:0] T_3339_coh_state;
  reg [31:0] GEN_136;
  wire [19:0] GEN_62;
  wire [1:0] GEN_63;
  wire  T_3423;
  wire  T_3424;
  reg [19:0] T_3425_tag;
  reg [31:0] GEN_137;
  reg [1:0] T_3425_coh_state;
  reg [31:0] GEN_138;
  wire [19:0] GEN_64;
  wire [1:0] GEN_65;
  wire  T_3509;
  wire  T_3510;
  reg [19:0] T_3511_tag;
  reg [31:0] GEN_139;
  reg [1:0] T_3511_coh_state;
  reg [31:0] GEN_140;
  wire [19:0] GEN_66;
  wire [1:0] GEN_67;
  wire [19:0] T_4264_0_tag;
  wire [1:0] T_4264_0_coh_state;
  wire [19:0] T_4264_1_tag;
  wire [1:0] T_4264_1_coh_state;
  wire [19:0] T_4264_2_tag;
  wire [1:0] T_4264_2_coh_state;
  wire [19:0] T_4264_3_tag;
  wire [1:0] T_4264_3_coh_state;
  wire  T_4681;
  wire  T_4682;
  wire  T_4683;
  wire  T_4684;
  wire [21:0] T_4685;
  wire [21:0] T_4687;
  wire [21:0] T_4688;
  wire [21:0] T_4690;
  wire [21:0] T_4691;
  wire [21:0] T_4693;
  wire [21:0] T_4694;
  wire [21:0] T_4696;
  wire [21:0] T_4781;
  wire [21:0] T_4782;
  wire [21:0] T_4783;
  wire [19:0] s2_repl_meta_tag;
  wire [1:0] s2_repl_meta_coh_state;
  wire [1:0] T_4951;
  wire [19:0] T_4952;
  wire  T_4954;
  wire  T_4955;
  wire  T_4956;
  wire  T_4958;
  wire  T_4959;
  wire  T_4961;
  wire  T_4963;
  wire  T_4967;
  wire  T_4968;
  wire  T_4976;
  wire  T_4977;
  wire [19:0] T_5062_tag;
  wire [1:0] T_5062_coh_state;
  wire [19:0] T_5146_tag;
  wire [1:0] T_5146_coh_state;
  wire [3:0] T_5230;
  wire  T_5231;
  wire  T_5235;
  wire  releaseArb_clk;
  wire  releaseArb_reset;
  wire  releaseArb_io_in_0_ready;
  wire  releaseArb_io_in_0_valid;
  wire [2:0] releaseArb_io_in_0_bits_addr_beat;
  wire [25:0] releaseArb_io_in_0_bits_addr_block;
  wire [1:0] releaseArb_io_in_0_bits_client_xact_id;
  wire  releaseArb_io_in_0_bits_voluntary;
  wire [2:0] releaseArb_io_in_0_bits_r_type;
  wire [63:0] releaseArb_io_in_0_bits_data;
  wire  releaseArb_io_in_1_ready;
  wire  releaseArb_io_in_1_valid;
  wire [2:0] releaseArb_io_in_1_bits_addr_beat;
  wire [25:0] releaseArb_io_in_1_bits_addr_block;
  wire [1:0] releaseArb_io_in_1_bits_client_xact_id;
  wire  releaseArb_io_in_1_bits_voluntary;
  wire [2:0] releaseArb_io_in_1_bits_r_type;
  wire [63:0] releaseArb_io_in_1_bits_data;
  wire  releaseArb_io_out_ready;
  wire  releaseArb_io_out_valid;
  wire [2:0] releaseArb_io_out_bits_addr_beat;
  wire [25:0] releaseArb_io_out_bits_addr_block;
  wire [1:0] releaseArb_io_out_bits_client_xact_id;
  wire  releaseArb_io_out_bits_voluntary;
  wire [2:0] releaseArb_io_out_bits_r_type;
  wire [63:0] releaseArb_io_out_bits_data;
  wire  releaseArb_io_chosen;
  wire  T_5265;
  wire  T_5268;
  wire  FlowThroughSerializer_1_1_clk;
  wire  FlowThroughSerializer_1_1_reset;
  wire  FlowThroughSerializer_1_1_io_in_ready;
  wire  FlowThroughSerializer_1_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_1_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_1_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_1_io_in_bits_manager_id;
  wire  FlowThroughSerializer_1_1_io_out_ready;
  wire  FlowThroughSerializer_1_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_1_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_1_1_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_1_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_1_io_out_bits_manager_id;
  wire  FlowThroughSerializer_1_1_io_cnt;
  wire  FlowThroughSerializer_1_1_io_done;
  wire  T_5269;
  wire [2:0] T_5277_0;
  wire [2:0] T_5277_1;
  wire [3:0] GEN_86;
  wire  T_5279;
  wire [3:0] GEN_87;
  wire  T_5280;
  wire  T_5281;
  wire  T_5282;
  wire  T_5283;
  wire  T_5285;
  wire  T_5286;
  wire [2:0] T_5294_0;
  wire [2:0] T_5294_1;
  wire [3:0] GEN_88;
  wire  T_5296;
  wire [3:0] GEN_89;
  wire  T_5297;
  wire  T_5298;
  wire  T_5300;
  wire  T_5301;
  wire  T_5303;
  wire  T_5304;
  wire [63:0] T_5307;
  wire  T_5309;
  wire  T_5310;
  wire  wbArb_clk;
  wire  wbArb_reset;
  wire  wbArb_io_in_0_ready;
  wire  wbArb_io_in_0_valid;
  wire [2:0] wbArb_io_in_0_bits_addr_beat;
  wire [25:0] wbArb_io_in_0_bits_addr_block;
  wire [1:0] wbArb_io_in_0_bits_client_xact_id;
  wire  wbArb_io_in_0_bits_voluntary;
  wire [2:0] wbArb_io_in_0_bits_r_type;
  wire [63:0] wbArb_io_in_0_bits_data;
  wire [3:0] wbArb_io_in_0_bits_way_en;
  wire  wbArb_io_in_1_ready;
  wire  wbArb_io_in_1_valid;
  wire [2:0] wbArb_io_in_1_bits_addr_beat;
  wire [25:0] wbArb_io_in_1_bits_addr_block;
  wire [1:0] wbArb_io_in_1_bits_client_xact_id;
  wire  wbArb_io_in_1_bits_voluntary;
  wire [2:0] wbArb_io_in_1_bits_r_type;
  wire [63:0] wbArb_io_in_1_bits_data;
  wire [3:0] wbArb_io_in_1_bits_way_en;
  wire  wbArb_io_out_ready;
  wire  wbArb_io_out_valid;
  wire [2:0] wbArb_io_out_bits_addr_beat;
  wire [25:0] wbArb_io_out_bits_addr_block;
  wire [1:0] wbArb_io_out_bits_client_xact_id;
  wire  wbArb_io_out_bits_voluntary;
  wire [2:0] wbArb_io_out_bits_r_type;
  wire [63:0] wbArb_io_out_bits_data;
  wire [3:0] wbArb_io_out_bits_way_en;
  wire  wbArb_io_chosen;
  reg  s4_valid;
  reg [31:0] GEN_141;
  wire  T_5360;
  reg [39:0] s4_req_addr;
  reg [63:0] GEN_142;
  reg [6:0] s4_req_tag;
  reg [31:0] GEN_143;
  reg [4:0] s4_req_cmd;
  reg [31:0] GEN_144;
  reg [2:0] s4_req_typ;
  reg [31:0] GEN_145;
  reg  s4_req_phys;
  reg [31:0] GEN_146;
  reg [63:0] s4_req_data;
  reg [63:0] GEN_147;
  wire [39:0] GEN_69;
  wire [6:0] GEN_70;
  wire [4:0] GEN_71;
  wire [2:0] GEN_72;
  wire  GEN_73;
  wire [63:0] GEN_74;
  wire  T_5427;
  wire  T_5430;
  wire [28:0] T_5431;
  wire [36:0] T_5432;
  wire [36:0] GEN_90;
  wire  T_5433;
  wire  T_5434;
  wire  T_5442;
  wire [36:0] T_5444;
  wire  T_5445;
  wire  T_5446;
  wire  T_5447;
  wire  T_5448;
  wire  T_5449;
  wire  T_5450;
  wire  T_5451;
  wire  T_5452;
  wire  T_5453;
  wire  T_5454;
  wire [36:0] T_5456;
  wire  T_5457;
  wire  T_5458;
  wire  T_5459;
  wire  T_5460;
  wire  T_5461;
  wire  T_5462;
  wire  T_5463;
  wire  T_5464;
  wire  T_5465;
  wire  T_5466;
  reg [63:0] s2_store_bypass_data;
  reg [63:0] GEN_148;
  reg  s2_store_bypass;
  reg [31:0] GEN_149;
  wire  T_5470;
  wire  T_5471;
  wire [63:0] T_5472;
  wire [63:0] T_5473;
  wire [63:0] GEN_75;
  wire  GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] s2_data_word_prebypass;
  wire [63:0] s2_data_word;
  wire  T_5477;
  wire  T_5479;
  wire [1:0] T_5480;
  wire  T_5481;
  wire [5:0] T_5482;
  wire  T_5483;
  wire  T_5485;
  wire  T_5486;
  wire  s1_nack;
  wire  T_5487;
  reg  s2_nack_hit;
  reg [31:0] GEN_150;
  wire  GEN_79;
  wire  GEN_80;
  wire  s2_nack_victim;
  wire  T_5492;
  wire  s2_nack_miss;
  wire  T_5493;
  wire  s2_nack;
  wire  T_5495;
  wire  T_5496;
  wire  T_5498;
  wire  s2_recycle_ecc;
  reg  s2_recycle_next;
  reg [31:0] GEN_151;
  wire  GEN_81;
  wire  T_5501;
  reg  block_miss;
  reg [31:0] GEN_152;
  wire  T_5503;
  wire  T_5504;
  wire  GEN_82;
  wire  cache_resp_valid;
  wire [39:0] cache_resp_bits_addr;
  wire [6:0] cache_resp_bits_tag;
  wire [4:0] cache_resp_bits_cmd;
  wire [2:0] cache_resp_bits_typ;
  wire [63:0] cache_resp_bits_data;
  wire  cache_resp_bits_replay;
  wire  cache_resp_bits_has_data;
  wire [63:0] cache_resp_bits_data_word_bypass;
  wire [63:0] cache_resp_bits_store_data;
  wire  T_5860;
  wire  T_5862;
  wire  T_5863;
  wire  T_5873;
  wire [31:0] T_5874;
  wire [31:0] T_5875;
  wire [31:0] T_5876;
  wire  T_5882;
  wire  T_5884;
  wire  T_5885;
  wire [31:0] T_5889;
  wire [31:0] T_5891;
  wire [63:0] T_5892;
  wire  T_5893;
  wire [15:0] T_5894;
  wire [15:0] T_5895;
  wire [15:0] T_5896;
  wire  T_5902;
  wire  T_5904;
  wire  T_5905;
  wire [47:0] T_5909;
  wire [47:0] T_5910;
  wire [47:0] T_5911;
  wire [63:0] T_5912;
  wire  T_5913;
  wire [7:0] T_5914;
  wire [7:0] T_5915;
  wire [7:0] T_5916;
  wire [7:0] T_5920;
  wire  T_5922;
  wire  T_5923;
  wire  T_5924;
  wire  T_5925;
  wire [55:0] T_5929;
  wire [55:0] T_5930;
  wire [55:0] T_5931;
  wire [63:0] T_5932;
  wire [63:0] GEN_93;
  wire [63:0] T_5933;
  wire  uncache_resp_valid;
  wire [39:0] uncache_resp_bits_addr;
  wire [6:0] uncache_resp_bits_tag;
  wire [4:0] uncache_resp_bits_cmd;
  wire [2:0] uncache_resp_bits_typ;
  wire [63:0] uncache_resp_bits_data;
  wire  uncache_resp_bits_replay;
  wire  uncache_resp_bits_has_data;
  wire [63:0] uncache_resp_bits_data_word_bypass;
  wire [63:0] uncache_resp_bits_store_data;
  wire  T_6289;
  reg  T_6290;
  reg [31:0] GEN_153;
  wire  T_6291;
  wire  T_6292_valid;
  wire [39:0] T_6292_bits_addr;
  wire [6:0] T_6292_bits_tag;
  wire [4:0] T_6292_bits_cmd;
  wire [2:0] T_6292_bits_typ;
  wire [63:0] T_6292_bits_data;
  wire  T_6292_bits_replay;
  wire  T_6292_bits_has_data;
  wire [63:0] T_6292_bits_store_data;
  wire  T_6456;
  wire  T_6458;
  wire  T_6459;
  wire  T_6460;
  wire  T_6461;
  wire [1:0] GEN_68;
  reg [31:0] GEN_154;
  wire [3:0] GEN_76;
  reg [31:0] GEN_155;
  wire [3:0] GEN_91;
  reg [31:0] GEN_156;
  wire [63:0] GEN_92;
  reg [63:0] GEN_157;
  WritebackUnit wb (
    .clk(wb_clk),
    .reset(wb_reset),
    .io_req_ready(wb_io_req_ready),
    .io_req_valid(wb_io_req_valid),
    .io_req_bits_addr_beat(wb_io_req_bits_addr_beat),
    .io_req_bits_addr_block(wb_io_req_bits_addr_block),
    .io_req_bits_client_xact_id(wb_io_req_bits_client_xact_id),
    .io_req_bits_voluntary(wb_io_req_bits_voluntary),
    .io_req_bits_r_type(wb_io_req_bits_r_type),
    .io_req_bits_data(wb_io_req_bits_data),
    .io_req_bits_way_en(wb_io_req_bits_way_en),
    .io_meta_read_ready(wb_io_meta_read_ready),
    .io_meta_read_valid(wb_io_meta_read_valid),
    .io_meta_read_bits_idx(wb_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(wb_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(wb_io_meta_read_bits_tag),
    .io_data_req_ready(wb_io_data_req_ready),
    .io_data_req_valid(wb_io_data_req_valid),
    .io_data_req_bits_way_en(wb_io_data_req_bits_way_en),
    .io_data_req_bits_addr(wb_io_data_req_bits_addr),
    .io_data_resp(wb_io_data_resp),
    .io_release_ready(wb_io_release_ready),
    .io_release_valid(wb_io_release_valid),
    .io_release_bits_addr_beat(wb_io_release_bits_addr_beat),
    .io_release_bits_addr_block(wb_io_release_bits_addr_block),
    .io_release_bits_client_xact_id(wb_io_release_bits_client_xact_id),
    .io_release_bits_voluntary(wb_io_release_bits_voluntary),
    .io_release_bits_r_type(wb_io_release_bits_r_type),
    .io_release_bits_data(wb_io_release_bits_data)
  );
  ProbeUnit prober (
    .clk(prober_clk),
    .reset(prober_reset),
    .io_req_ready(prober_io_req_ready),
    .io_req_valid(prober_io_req_valid),
    .io_req_bits_addr_block(prober_io_req_bits_addr_block),
    .io_req_bits_p_type(prober_io_req_bits_p_type),
    .io_req_bits_client_xact_id(prober_io_req_bits_client_xact_id),
    .io_rep_ready(prober_io_rep_ready),
    .io_rep_valid(prober_io_rep_valid),
    .io_rep_bits_addr_beat(prober_io_rep_bits_addr_beat),
    .io_rep_bits_addr_block(prober_io_rep_bits_addr_block),
    .io_rep_bits_client_xact_id(prober_io_rep_bits_client_xact_id),
    .io_rep_bits_voluntary(prober_io_rep_bits_voluntary),
    .io_rep_bits_r_type(prober_io_rep_bits_r_type),
    .io_rep_bits_data(prober_io_rep_bits_data),
    .io_meta_read_ready(prober_io_meta_read_ready),
    .io_meta_read_valid(prober_io_meta_read_valid),
    .io_meta_read_bits_idx(prober_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(prober_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(prober_io_meta_read_bits_tag),
    .io_meta_write_ready(prober_io_meta_write_ready),
    .io_meta_write_valid(prober_io_meta_write_valid),
    .io_meta_write_bits_idx(prober_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(prober_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(prober_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(prober_io_meta_write_bits_data_coh_state),
    .io_wb_req_ready(prober_io_wb_req_ready),
    .io_wb_req_valid(prober_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(prober_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(prober_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(prober_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(prober_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(prober_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(prober_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(prober_io_wb_req_bits_way_en),
    .io_way_en(prober_io_way_en),
    .io_mshr_rdy(prober_io_mshr_rdy),
    .io_block_state_state(prober_io_block_state_state)
  );
  MSHRFile mshrs (
    .clk(mshrs_clk),
    .reset(mshrs_reset),
    .io_req_ready(mshrs_io_req_ready),
    .io_req_valid(mshrs_io_req_valid),
    .io_req_bits_addr(mshrs_io_req_bits_addr),
    .io_req_bits_tag(mshrs_io_req_bits_tag),
    .io_req_bits_cmd(mshrs_io_req_bits_cmd),
    .io_req_bits_typ(mshrs_io_req_bits_typ),
    .io_req_bits_phys(mshrs_io_req_bits_phys),
    .io_req_bits_data(mshrs_io_req_bits_data),
    .io_req_bits_tag_match(mshrs_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(mshrs_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(mshrs_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(mshrs_io_req_bits_way_en),
    .io_resp_ready(mshrs_io_resp_ready),
    .io_resp_valid(mshrs_io_resp_valid),
    .io_resp_bits_addr(mshrs_io_resp_bits_addr),
    .io_resp_bits_tag(mshrs_io_resp_bits_tag),
    .io_resp_bits_cmd(mshrs_io_resp_bits_cmd),
    .io_resp_bits_typ(mshrs_io_resp_bits_typ),
    .io_resp_bits_data(mshrs_io_resp_bits_data),
    .io_resp_bits_replay(mshrs_io_resp_bits_replay),
    .io_resp_bits_has_data(mshrs_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(mshrs_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(mshrs_io_resp_bits_store_data),
    .io_secondary_miss(mshrs_io_secondary_miss),
    .io_mem_req_ready(mshrs_io_mem_req_ready),
    .io_mem_req_valid(mshrs_io_mem_req_valid),
    .io_mem_req_bits_addr_block(mshrs_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(mshrs_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(mshrs_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(mshrs_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(mshrs_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(mshrs_io_mem_req_bits_union),
    .io_mem_req_bits_data(mshrs_io_mem_req_bits_data),
    .io_refill_way_en(mshrs_io_refill_way_en),
    .io_refill_addr(mshrs_io_refill_addr),
    .io_meta_read_ready(mshrs_io_meta_read_ready),
    .io_meta_read_valid(mshrs_io_meta_read_valid),
    .io_meta_read_bits_idx(mshrs_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(mshrs_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(mshrs_io_meta_read_bits_tag),
    .io_meta_write_ready(mshrs_io_meta_write_ready),
    .io_meta_write_valid(mshrs_io_meta_write_valid),
    .io_meta_write_bits_idx(mshrs_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(mshrs_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(mshrs_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(mshrs_io_meta_write_bits_data_coh_state),
    .io_replay_ready(mshrs_io_replay_ready),
    .io_replay_valid(mshrs_io_replay_valid),
    .io_replay_bits_addr(mshrs_io_replay_bits_addr),
    .io_replay_bits_tag(mshrs_io_replay_bits_tag),
    .io_replay_bits_cmd(mshrs_io_replay_bits_cmd),
    .io_replay_bits_typ(mshrs_io_replay_bits_typ),
    .io_replay_bits_phys(mshrs_io_replay_bits_phys),
    .io_replay_bits_data(mshrs_io_replay_bits_data),
    .io_mem_grant_valid(mshrs_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(mshrs_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(mshrs_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(mshrs_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(mshrs_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(mshrs_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(mshrs_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(mshrs_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(mshrs_io_mem_finish_ready),
    .io_mem_finish_valid(mshrs_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(mshrs_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(mshrs_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(mshrs_io_wb_req_ready),
    .io_wb_req_valid(mshrs_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(mshrs_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(mshrs_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(mshrs_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(mshrs_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(mshrs_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(mshrs_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(mshrs_io_wb_req_bits_way_en),
    .io_probe_rdy(mshrs_io_probe_rdy),
    .io_fence_rdy(mshrs_io_fence_rdy),
    .io_replay_next(mshrs_io_replay_next)
  );
  TLB dtlb (
    .clk(dtlb_clk),
    .reset(dtlb_reset),
    .io_req_ready(dtlb_io_req_ready),
    .io_req_valid(dtlb_io_req_valid),
    .io_req_bits_vpn(dtlb_io_req_bits_vpn),
    .io_req_bits_passthrough(dtlb_io_req_bits_passthrough),
    .io_req_bits_instruction(dtlb_io_req_bits_instruction),
    .io_req_bits_store(dtlb_io_req_bits_store),
    .io_resp_miss(dtlb_io_resp_miss),
    .io_resp_ppn(dtlb_io_resp_ppn),
    .io_resp_xcpt_ld(dtlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(dtlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(dtlb_io_resp_xcpt_if),
    .io_resp_cacheable(dtlb_io_resp_cacheable),
    .io_ptw_req_ready(dtlb_io_ptw_req_ready),
    .io_ptw_req_valid(dtlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(dtlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(dtlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(dtlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(dtlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(dtlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(dtlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(dtlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(dtlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(dtlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(dtlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(dtlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(dtlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(dtlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(dtlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(dtlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(dtlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(dtlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(dtlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(dtlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(dtlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(dtlb_io_ptw_invalidate),
    .io_ptw_status_debug(dtlb_io_ptw_status_debug),
    .io_ptw_status_prv(dtlb_io_ptw_status_prv),
    .io_ptw_status_sd(dtlb_io_ptw_status_sd),
    .io_ptw_status_zero3(dtlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(dtlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(dtlb_io_ptw_status_zero2),
    .io_ptw_status_vm(dtlb_io_ptw_status_vm),
    .io_ptw_status_zero1(dtlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(dtlb_io_ptw_status_mxr),
    .io_ptw_status_pum(dtlb_io_ptw_status_pum),
    .io_ptw_status_mprv(dtlb_io_ptw_status_mprv),
    .io_ptw_status_xs(dtlb_io_ptw_status_xs),
    .io_ptw_status_fs(dtlb_io_ptw_status_fs),
    .io_ptw_status_mpp(dtlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(dtlb_io_ptw_status_hpp),
    .io_ptw_status_spp(dtlb_io_ptw_status_spp),
    .io_ptw_status_mpie(dtlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(dtlb_io_ptw_status_hpie),
    .io_ptw_status_spie(dtlb_io_ptw_status_spie),
    .io_ptw_status_upie(dtlb_io_ptw_status_upie),
    .io_ptw_status_mie(dtlb_io_ptw_status_mie),
    .io_ptw_status_hie(dtlb_io_ptw_status_hie),
    .io_ptw_status_sie(dtlb_io_ptw_status_sie),
    .io_ptw_status_uie(dtlb_io_ptw_status_uie)
  );
  MetadataArray meta (
    .clk(meta_clk),
    .reset(meta_reset),
    .io_read_ready(meta_io_read_ready),
    .io_read_valid(meta_io_read_valid),
    .io_read_bits_idx(meta_io_read_bits_idx),
    .io_read_bits_way_en(meta_io_read_bits_way_en),
    .io_write_ready(meta_io_write_ready),
    .io_write_valid(meta_io_write_valid),
    .io_write_bits_idx(meta_io_write_bits_idx),
    .io_write_bits_way_en(meta_io_write_bits_way_en),
    .io_write_bits_data_tag(meta_io_write_bits_data_tag),
    .io_write_bits_data_coh_state(meta_io_write_bits_data_coh_state),
    .io_resp_0_tag(meta_io_resp_0_tag),
    .io_resp_0_coh_state(meta_io_resp_0_coh_state),
    .io_resp_1_tag(meta_io_resp_1_tag),
    .io_resp_1_coh_state(meta_io_resp_1_coh_state),
    .io_resp_2_tag(meta_io_resp_2_tag),
    .io_resp_2_coh_state(meta_io_resp_2_coh_state),
    .io_resp_3_tag(meta_io_resp_3_tag),
    .io_resp_3_coh_state(meta_io_resp_3_coh_state)
  );
  Arbiter_8 metaReadArb (
    .clk(metaReadArb_clk),
    .reset(metaReadArb_reset),
    .io_in_0_ready(metaReadArb_io_in_0_ready),
    .io_in_0_valid(metaReadArb_io_in_0_valid),
    .io_in_0_bits_idx(metaReadArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaReadArb_io_in_0_bits_way_en),
    .io_in_1_ready(metaReadArb_io_in_1_ready),
    .io_in_1_valid(metaReadArb_io_in_1_valid),
    .io_in_1_bits_idx(metaReadArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaReadArb_io_in_1_bits_way_en),
    .io_in_2_ready(metaReadArb_io_in_2_ready),
    .io_in_2_valid(metaReadArb_io_in_2_valid),
    .io_in_2_bits_idx(metaReadArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaReadArb_io_in_2_bits_way_en),
    .io_in_3_ready(metaReadArb_io_in_3_ready),
    .io_in_3_valid(metaReadArb_io_in_3_valid),
    .io_in_3_bits_idx(metaReadArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaReadArb_io_in_3_bits_way_en),
    .io_in_4_ready(metaReadArb_io_in_4_ready),
    .io_in_4_valid(metaReadArb_io_in_4_valid),
    .io_in_4_bits_idx(metaReadArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaReadArb_io_in_4_bits_way_en),
    .io_out_ready(metaReadArb_io_out_ready),
    .io_out_valid(metaReadArb_io_out_valid),
    .io_out_bits_idx(metaReadArb_io_out_bits_idx),
    .io_out_bits_way_en(metaReadArb_io_out_bits_way_en),
    .io_chosen(metaReadArb_io_chosen)
  );
  Arbiter_1 metaWriteArb (
    .clk(metaWriteArb_clk),
    .reset(metaWriteArb_reset),
    .io_in_0_ready(metaWriteArb_io_in_0_ready),
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_idx(metaWriteArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaWriteArb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(metaWriteArb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(metaWriteArb_io_in_1_ready),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_idx(metaWriteArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaWriteArb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(metaWriteArb_io_in_1_bits_data_coh_state),
    .io_out_ready(metaWriteArb_io_out_ready),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_idx(metaWriteArb_io_out_bits_idx),
    .io_out_bits_way_en(metaWriteArb_io_out_bits_way_en),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(metaWriteArb_io_out_bits_data_coh_state),
    .io_chosen(metaWriteArb_io_chosen)
  );
  DataArray data (
    .clk(data_clk),
    .reset(data_reset),
    .io_read_ready(data_io_read_ready),
    .io_read_valid(data_io_read_valid),
    .io_read_bits_way_en(data_io_read_bits_way_en),
    .io_read_bits_addr(data_io_read_bits_addr),
    .io_write_ready(data_io_write_ready),
    .io_write_valid(data_io_write_valid),
    .io_write_bits_way_en(data_io_write_bits_way_en),
    .io_write_bits_addr(data_io_write_bits_addr),
    .io_write_bits_wmask(data_io_write_bits_wmask),
    .io_write_bits_data(data_io_write_bits_data),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  Arbiter_10 readArb (
    .clk(readArb_clk),
    .reset(readArb_reset),
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_way_en(readArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(readArb_io_in_0_bits_addr),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_way_en(readArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(readArb_io_in_1_bits_addr),
    .io_in_2_ready(readArb_io_in_2_ready),
    .io_in_2_valid(readArb_io_in_2_valid),
    .io_in_2_bits_way_en(readArb_io_in_2_bits_way_en),
    .io_in_2_bits_addr(readArb_io_in_2_bits_addr),
    .io_in_3_ready(readArb_io_in_3_ready),
    .io_in_3_valid(readArb_io_in_3_valid),
    .io_in_3_bits_way_en(readArb_io_in_3_bits_way_en),
    .io_in_3_bits_addr(readArb_io_in_3_bits_addr),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_way_en(readArb_io_out_bits_way_en),
    .io_out_bits_addr(readArb_io_out_bits_addr),
    .io_chosen(readArb_io_chosen)
  );
  Arbiter_11 writeArb (
    .clk(writeArb_clk),
    .reset(writeArb_reset),
    .io_in_0_ready(writeArb_io_in_0_ready),
    .io_in_0_valid(writeArb_io_in_0_valid),
    .io_in_0_bits_way_en(writeArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(writeArb_io_in_0_bits_addr),
    .io_in_0_bits_wmask(writeArb_io_in_0_bits_wmask),
    .io_in_0_bits_data(writeArb_io_in_0_bits_data),
    .io_in_1_ready(writeArb_io_in_1_ready),
    .io_in_1_valid(writeArb_io_in_1_valid),
    .io_in_1_bits_way_en(writeArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(writeArb_io_in_1_bits_addr),
    .io_in_1_bits_wmask(writeArb_io_in_1_bits_wmask),
    .io_in_1_bits_data(writeArb_io_in_1_bits_data),
    .io_out_ready(writeArb_io_out_ready),
    .io_out_valid(writeArb_io_out_valid),
    .io_out_bits_way_en(writeArb_io_out_bits_way_en),
    .io_out_bits_addr(writeArb_io_out_bits_addr),
    .io_out_bits_wmask(writeArb_io_out_bits_wmask),
    .io_out_bits_data(writeArb_io_out_bits_data),
    .io_chosen(writeArb_io_chosen)
  );
  AMOALU amoalu (
    .clk(amoalu_clk),
    .reset(amoalu_reset),
    .io_addr(amoalu_io_addr),
    .io_cmd(amoalu_io_cmd),
    .io_typ(amoalu_io_typ),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  LockingArbiter_1 releaseArb (
    .clk(releaseArb_clk),
    .reset(releaseArb_reset),
    .io_in_0_ready(releaseArb_io_in_0_ready),
    .io_in_0_valid(releaseArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(releaseArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(releaseArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(releaseArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(releaseArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(releaseArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(releaseArb_io_in_0_bits_data),
    .io_in_1_ready(releaseArb_io_in_1_ready),
    .io_in_1_valid(releaseArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(releaseArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(releaseArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(releaseArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(releaseArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(releaseArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(releaseArb_io_in_1_bits_data),
    .io_out_ready(releaseArb_io_out_ready),
    .io_out_valid(releaseArb_io_out_valid),
    .io_out_bits_addr_beat(releaseArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(releaseArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(releaseArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(releaseArb_io_out_bits_voluntary),
    .io_out_bits_r_type(releaseArb_io_out_bits_r_type),
    .io_out_bits_data(releaseArb_io_out_bits_data),
    .io_chosen(releaseArb_io_chosen)
  );
  FlowThroughSerializer_1 FlowThroughSerializer_1_1 (
    .clk(FlowThroughSerializer_1_1_clk),
    .reset(FlowThroughSerializer_1_1_reset),
    .io_in_ready(FlowThroughSerializer_1_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_1_io_in_bits_data),
    .io_in_bits_manager_id(FlowThroughSerializer_1_1_io_in_bits_manager_id),
    .io_out_ready(FlowThroughSerializer_1_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_1_io_out_bits_data),
    .io_out_bits_manager_id(FlowThroughSerializer_1_1_io_out_bits_manager_id),
    .io_cnt(FlowThroughSerializer_1_1_io_cnt),
    .io_done(FlowThroughSerializer_1_1_io_done)
  );
  Arbiter_3 wbArb (
    .clk(wbArb_clk),
    .reset(wbArb_reset),
    .io_in_0_ready(wbArb_io_in_0_ready),
    .io_in_0_valid(wbArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wbArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wbArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wbArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wbArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wbArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wbArb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wbArb_io_in_0_bits_way_en),
    .io_in_1_ready(wbArb_io_in_1_ready),
    .io_in_1_valid(wbArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wbArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wbArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wbArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wbArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wbArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wbArb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wbArb_io_in_1_bits_way_en),
    .io_out_ready(wbArb_io_out_ready),
    .io_out_valid(wbArb_io_out_valid),
    .io_out_bits_addr_beat(wbArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wbArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wbArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wbArb_io_out_bits_voluntary),
    .io_out_bits_r_type(wbArb_io_out_bits_r_type),
    .io_out_bits_data(wbArb_io_out_bits_data),
    .io_out_bits_way_en(wbArb_io_out_bits_way_en),
    .io_chosen(wbArb_io_chosen)
  );
  assign io_cpu_req_ready = GEN_82;
  assign io_cpu_s2_nack = T_6291;
  assign io_cpu_resp_valid = T_6292_valid;
  assign io_cpu_resp_bits_addr = T_6292_bits_addr;
  assign io_cpu_resp_bits_tag = T_6292_bits_tag;
  assign io_cpu_resp_bits_cmd = T_6292_bits_cmd;
  assign io_cpu_resp_bits_typ = T_6292_bits_typ;
  assign io_cpu_resp_bits_data = T_6292_bits_data;
  assign io_cpu_resp_bits_replay = T_6292_bits_replay;
  assign io_cpu_resp_bits_has_data = T_6292_bits_has_data;
  assign io_cpu_resp_bits_data_word_bypass = T_5892;
  assign io_cpu_resp_bits_store_data = T_6292_bits_store_data;
  assign io_cpu_replay_next = T_6461;
  assign io_cpu_xcpt_ma_ld = T_2167;
  assign io_cpu_xcpt_ma_st = T_2168;
  assign io_cpu_xcpt_pf_ld = T_2169;
  assign io_cpu_xcpt_pf_st = T_2170;
  assign io_cpu_ordered = T_6459;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = dtlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = dtlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_probe_ready = T_5268;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_1_io_in_ready;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_finish_bits_manager_xact_id = mshrs_io_mem_finish_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mshrs_io_mem_finish_bits_manager_id;
  assign wb_clk = clk;
  assign wb_reset = reset;
  assign wb_io_req_valid = wbArb_io_out_valid;
  assign wb_io_req_bits_addr_beat = wbArb_io_out_bits_addr_beat;
  assign wb_io_req_bits_addr_block = wbArb_io_out_bits_addr_block;
  assign wb_io_req_bits_client_xact_id = wbArb_io_out_bits_client_xact_id;
  assign wb_io_req_bits_voluntary = wbArb_io_out_bits_voluntary;
  assign wb_io_req_bits_r_type = wbArb_io_out_bits_r_type;
  assign wb_io_req_bits_data = wbArb_io_out_bits_data;
  assign wb_io_req_bits_way_en = wbArb_io_out_bits_way_en;
  assign wb_io_meta_read_ready = metaReadArb_io_in_3_ready;
  assign wb_io_data_req_ready = readArb_io_in_2_ready;
  assign wb_io_data_resp = s2_data_muxed;
  assign wb_io_release_ready = releaseArb_io_in_0_ready;
  assign prober_clk = clk;
  assign prober_reset = reset;
  assign prober_io_req_valid = T_5265;
  assign prober_io_req_bits_addr_block = io_mem_probe_bits_addr_block;
  assign prober_io_req_bits_p_type = io_mem_probe_bits_p_type;
  assign prober_io_req_bits_client_xact_id = GEN_68;
  assign prober_io_rep_ready = releaseArb_io_in_1_ready;
  assign prober_io_meta_read_ready = metaReadArb_io_in_2_ready;
  assign prober_io_meta_write_ready = metaWriteArb_io_in_1_ready;
  assign prober_io_wb_req_ready = wbArb_io_in_0_ready;
  assign prober_io_way_en = s2_tag_match_way;
  assign prober_io_mshr_rdy = mshrs_io_probe_rdy;
  assign prober_io_block_state_state = s2_hit_state_state;
  assign mshrs_clk = clk;
  assign mshrs_reset = reset;
  assign mshrs_io_req_valid = GEN_80;
  assign mshrs_io_req_bits_addr = s2_req_addr;
  assign mshrs_io_req_bits_tag = s2_req_tag;
  assign mshrs_io_req_bits_cmd = s2_req_cmd;
  assign mshrs_io_req_bits_typ = s2_req_typ;
  assign mshrs_io_req_bits_phys = s2_req_phys;
  assign mshrs_io_req_bits_data = s2_req_data;
  assign mshrs_io_req_bits_tag_match = s2_tag_match;
  assign mshrs_io_req_bits_old_meta_tag = T_5146_tag;
  assign mshrs_io_req_bits_old_meta_coh_state = T_5146_coh_state;
  assign mshrs_io_req_bits_way_en = T_5230;
  assign mshrs_io_resp_ready = T_6290;
  assign mshrs_io_mem_req_ready = io_mem_acquire_ready;
  assign mshrs_io_meta_read_ready = metaReadArb_io_in_1_ready;
  assign mshrs_io_meta_write_ready = metaWriteArb_io_in_0_ready;
  assign mshrs_io_replay_ready = readArb_io_in_1_ready;
  assign mshrs_io_mem_grant_valid = T_5269;
  assign mshrs_io_mem_grant_bits_addr_beat = FlowThroughSerializer_1_1_io_out_bits_addr_beat;
  assign mshrs_io_mem_grant_bits_client_xact_id = FlowThroughSerializer_1_1_io_out_bits_client_xact_id;
  assign mshrs_io_mem_grant_bits_manager_xact_id = FlowThroughSerializer_1_1_io_out_bits_manager_xact_id;
  assign mshrs_io_mem_grant_bits_is_builtin_type = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type;
  assign mshrs_io_mem_grant_bits_g_type = FlowThroughSerializer_1_1_io_out_bits_g_type;
  assign mshrs_io_mem_grant_bits_data = FlowThroughSerializer_1_1_io_out_bits_data;
  assign mshrs_io_mem_grant_bits_manager_id = FlowThroughSerializer_1_1_io_out_bits_manager_id;
  assign mshrs_io_mem_finish_ready = io_mem_finish_ready;
  assign mshrs_io_wb_req_ready = wbArb_io_in_1_ready;
  assign T_1901 = io_cpu_req_ready & io_cpu_req_valid;
  assign T_1970 = io_cpu_s1_kill == 1'h0;
  assign T_1971 = s1_valid & T_1970;
  assign T_1972 = {io_cpu_xcpt_pf_ld,io_cpu_xcpt_pf_st};
  assign T_1973 = {io_cpu_xcpt_ma_ld,io_cpu_xcpt_ma_st};
  assign T_1974 = {T_1973,T_1972};
  assign T_1976 = T_1974 != 4'h0;
  assign T_1978 = T_1976 == 1'h0;
  assign s1_valid_masked = T_1971 & T_1978;
  assign T_2050 = s2_req_cmd != 5'h5;
  assign s2_replay = T_2049 & T_2050;
  assign s2_recycle = T_5501;
  assign s2_valid_masked = T_5496;
  assign GEN_0 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T_2122 = s1_req_cmd == 5'h0;
  assign T_2123 = s1_req_cmd == 5'h6;
  assign T_2124 = T_2122 | T_2123;
  assign T_2125 = s1_req_cmd == 5'h7;
  assign T_2126 = T_2124 | T_2125;
  assign T_2127 = s1_req_cmd[3];
  assign T_2128 = s1_req_cmd == 5'h4;
  assign T_2129 = T_2127 | T_2128;
  assign s1_read = T_2126 | T_2129;
  assign T_2130 = s1_req_cmd == 5'h1;
  assign T_2132 = T_2130 | T_2125;
  assign s1_write = T_2132 | T_2129;
  assign T_2136 = s1_read | s1_write;
  assign T_2137 = s1_req_cmd == 5'h2;
  assign T_2138 = s1_req_cmd == 5'h3;
  assign T_2139 = T_2137 | T_2138;
  assign s1_readwrite = T_2136 | T_2139;
  assign dtlb_clk = clk;
  assign dtlb_reset = reset;
  assign dtlb_io_req_valid = T_2140;
  assign dtlb_io_req_bits_vpn = T_2141;
  assign dtlb_io_req_bits_passthrough = s1_req_phys;
  assign dtlb_io_req_bits_instruction = 1'h0;
  assign dtlb_io_req_bits_store = s1_write;
  assign dtlb_io_ptw_req_ready = io_ptw_req_ready;
  assign dtlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign dtlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign dtlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign dtlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign dtlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign dtlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign dtlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign dtlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign dtlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign dtlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign dtlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign dtlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign dtlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign dtlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign dtlb_io_ptw_invalidate = io_ptw_invalidate;
  assign dtlb_io_ptw_status_debug = io_ptw_status_debug;
  assign dtlb_io_ptw_status_prv = io_ptw_status_prv;
  assign dtlb_io_ptw_status_sd = io_ptw_status_sd;
  assign dtlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign dtlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign dtlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign dtlb_io_ptw_status_vm = io_ptw_status_vm;
  assign dtlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign dtlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign dtlb_io_ptw_status_pum = io_ptw_status_pum;
  assign dtlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign dtlb_io_ptw_status_xs = io_ptw_status_xs;
  assign dtlb_io_ptw_status_fs = io_ptw_status_fs;
  assign dtlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign dtlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign dtlb_io_ptw_status_spp = io_ptw_status_spp;
  assign dtlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign dtlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign dtlb_io_ptw_status_spie = io_ptw_status_spie;
  assign dtlb_io_ptw_status_upie = io_ptw_status_upie;
  assign dtlb_io_ptw_status_mie = io_ptw_status_mie;
  assign dtlb_io_ptw_status_hie = io_ptw_status_hie;
  assign dtlb_io_ptw_status_sie = io_ptw_status_sie;
  assign dtlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_2140 = s1_valid_masked & s1_readwrite;
  assign T_2141 = s1_req_addr[39:12];
  assign T_2144 = dtlb_io_req_ready == 1'h0;
  assign T_2146 = io_cpu_req_bits_phys == 1'h0;
  assign T_2147 = T_2144 & T_2146;
  assign GEN_1 = T_2147 ? 1'h0 : 1'h1;
  assign GEN_2 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign GEN_3 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign GEN_4 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign GEN_5 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign GEN_6 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign GEN_7 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T_2149 = {wb_io_meta_read_bits_tag,wb_io_meta_read_bits_idx};
  assign GEN_83 = {{6'd0}, T_2149};
  assign T_2150 = GEN_83 << 6;
  assign GEN_8 = wb_io_meta_read_valid ? {{8'd0}, T_2150} : GEN_2;
  assign GEN_9 = wb_io_meta_read_valid ? 1'h1 : GEN_6;
  assign T_2152 = {prober_io_meta_read_bits_tag,prober_io_meta_read_bits_idx};
  assign GEN_84 = {{6'd0}, T_2152};
  assign T_2153 = GEN_84 << 6;
  assign GEN_10 = prober_io_meta_read_valid ? {{8'd0}, T_2153} : GEN_8;
  assign GEN_11 = prober_io_meta_read_valid ? 1'h1 : GEN_9;
  assign GEN_12 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : GEN_10;
  assign GEN_13 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : GEN_3;
  assign GEN_14 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : GEN_4;
  assign GEN_15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : GEN_5;
  assign GEN_16 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : GEN_11;
  assign GEN_17 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : GEN_7;
  assign GEN_18 = s2_recycle ? s2_req_addr : GEN_12;
  assign GEN_19 = s2_recycle ? s2_req_tag : GEN_13;
  assign GEN_20 = s2_recycle ? s2_req_cmd : GEN_14;
  assign GEN_21 = s2_recycle ? s2_req_typ : GEN_15;
  assign GEN_22 = s2_recycle ? s2_req_phys : GEN_16;
  assign GEN_23 = s2_recycle ? s2_req_data : GEN_17;
  assign T_2155 = s1_req_addr[11:0];
  assign s1_addr = {dtlb_io_resp_ppn,T_2155};
  assign T_2156 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_s1_data;
  assign GEN_24 = s1_write ? T_2156 : s2_req_data;
  assign GEN_25 = s1_recycled ? s1_req_data : GEN_24;
  assign GEN_26 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign GEN_27 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign GEN_28 = s1_clk_en ? {{8'd0}, s1_addr} : s2_req_addr;
  assign GEN_29 = s1_clk_en ? GEN_25 : s2_req_data;
  assign GEN_30 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign GEN_31 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign T_2158 = s1_req_typ[1:0];
  assign T_2160 = 4'h1 << T_2158;
  assign T_2162 = T_2160 - 4'h1;
  assign T_2163 = T_2162[3:0];
  assign T_2164 = T_2163[2:0];
  assign GEN_85 = {{37'd0}, T_2164};
  assign T_2165 = s1_req_addr & GEN_85;
  assign misaligned = T_2165 != 40'h0;
  assign T_2167 = s1_read & misaligned;
  assign T_2168 = s1_write & misaligned;
  assign T_2169 = s1_read & dtlb_io_resp_xcpt_ld;
  assign T_2170 = s1_write & dtlb_io_resp_xcpt_st;
  assign meta_clk = clk;
  assign meta_reset = reset;
  assign meta_io_read_valid = metaReadArb_io_out_valid;
  assign meta_io_read_bits_idx = metaReadArb_io_out_bits_idx;
  assign meta_io_read_bits_way_en = metaReadArb_io_out_bits_way_en;
  assign meta_io_write_valid = metaWriteArb_io_out_valid;
  assign meta_io_write_bits_idx = metaWriteArb_io_out_bits_idx;
  assign meta_io_write_bits_way_en = metaWriteArb_io_out_bits_way_en;
  assign meta_io_write_bits_data_tag = metaWriteArb_io_out_bits_data_tag;
  assign meta_io_write_bits_data_coh_state = metaWriteArb_io_out_bits_data_coh_state;
  assign metaReadArb_clk = clk;
  assign metaReadArb_reset = reset;
  assign metaReadArb_io_in_0_valid = s2_recycle;
  assign metaReadArb_io_in_0_bits_idx = T_2522[5:0];
  assign metaReadArb_io_in_0_bits_way_en = GEN_76;
  assign metaReadArb_io_in_1_valid = mshrs_io_meta_read_valid;
  assign metaReadArb_io_in_1_bits_idx = mshrs_io_meta_read_bits_idx;
  assign metaReadArb_io_in_1_bits_way_en = mshrs_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_2_valid = prober_io_meta_read_valid;
  assign metaReadArb_io_in_2_bits_idx = prober_io_meta_read_bits_idx;
  assign metaReadArb_io_in_2_bits_way_en = prober_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_3_valid = wb_io_meta_read_valid;
  assign metaReadArb_io_in_3_bits_idx = wb_io_meta_read_bits_idx;
  assign metaReadArb_io_in_3_bits_way_en = wb_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_4_valid = io_cpu_req_valid;
  assign metaReadArb_io_in_4_bits_idx = T_2513[5:0];
  assign metaReadArb_io_in_4_bits_way_en = GEN_91;
  assign metaReadArb_io_out_ready = meta_io_read_ready;
  assign metaWriteArb_clk = clk;
  assign metaWriteArb_reset = reset;
  assign metaWriteArb_io_in_0_valid = mshrs_io_meta_write_valid;
  assign metaWriteArb_io_in_0_bits_idx = mshrs_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_0_bits_way_en = mshrs_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_0_bits_data_tag = mshrs_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_0_bits_data_coh_state = mshrs_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_in_1_valid = prober_io_meta_write_valid;
  assign metaWriteArb_io_in_1_bits_idx = prober_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_1_bits_way_en = prober_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_1_bits_data_tag = prober_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_1_bits_data_coh_state = prober_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_out_ready = meta_io_write_ready;
  assign data_clk = clk;
  assign data_reset = reset;
  assign data_io_read_valid = readArb_io_out_valid;
  assign data_io_read_bits_way_en = readArb_io_out_bits_way_en;
  assign data_io_read_bits_addr = readArb_io_out_bits_addr;
  assign data_io_write_valid = writeArb_io_out_valid;
  assign data_io_write_bits_way_en = writeArb_io_out_bits_way_en;
  assign data_io_write_bits_addr = writeArb_io_out_bits_addr;
  assign data_io_write_bits_wmask = writeArb_io_out_bits_wmask;
  assign data_io_write_bits_data = wdata_encoded_0;
  assign readArb_clk = clk;
  assign readArb_reset = reset;
  assign readArb_io_in_0_valid = s2_recycle;
  assign readArb_io_in_0_bits_way_en = 4'hf;
  assign readArb_io_in_0_bits_addr = s2_req_addr[11:0];
  assign readArb_io_in_1_valid = mshrs_io_replay_valid;
  assign readArb_io_in_1_bits_way_en = 4'hf;
  assign readArb_io_in_1_bits_addr = mshrs_io_replay_bits_addr[11:0];
  assign readArb_io_in_2_valid = wb_io_data_req_valid;
  assign readArb_io_in_2_bits_way_en = wb_io_data_req_bits_way_en;
  assign readArb_io_in_2_bits_addr = wb_io_data_req_bits_addr;
  assign readArb_io_in_3_valid = io_cpu_req_valid;
  assign readArb_io_in_3_bits_way_en = 4'hf;
  assign readArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0];
  assign readArb_io_out_ready = T_5310;
  assign writeArb_clk = clk;
  assign writeArb_reset = reset;
  assign writeArb_io_in_0_valid = s3_valid;
  assign writeArb_io_in_0_bits_way_en = s3_way;
  assign writeArb_io_in_0_bits_addr = s3_req_addr[11:0];
  assign writeArb_io_in_0_bits_wmask = T_3231[0];
  assign writeArb_io_in_0_bits_data = s3_req_data;
  assign writeArb_io_in_1_valid = T_5304;
  assign writeArb_io_in_1_bits_way_en = mshrs_io_refill_way_en;
  assign writeArb_io_in_1_bits_addr = mshrs_io_refill_addr;
  assign writeArb_io_in_1_bits_wmask = 1'h1;
  assign writeArb_io_in_1_bits_data = T_5307;
  assign writeArb_io_out_ready = data_io_write_ready;
  assign wdata_encoded_0 = writeArb_io_out_bits_data;
  assign T_2513 = io_cpu_req_bits_addr[39:6];
  assign T_2515 = metaReadArb_io_in_4_ready == 1'h0;
  assign GEN_32 = T_2515 ? 1'h0 : GEN_1;
  assign T_2520 = readArb_io_in_3_ready == 1'h0;
  assign GEN_33 = T_2520 ? 1'h0 : GEN_32;
  assign T_2522 = s2_req_addr[39:6];
  assign T_2525 = s1_addr[31:12];
  assign T_2526 = meta_io_resp_0_tag == T_2525;
  assign T_2528 = meta_io_resp_1_tag == T_2525;
  assign T_2530 = meta_io_resp_2_tag == T_2525;
  assign T_2532 = meta_io_resp_3_tag == T_2525;
  assign T_2538_0 = T_2526;
  assign T_2538_1 = T_2528;
  assign T_2538_2 = T_2530;
  assign T_2538_3 = T_2532;
  assign T_2540 = {T_2538_1,T_2538_0};
  assign T_2541 = {T_2538_3,T_2538_2};
  assign s1_tag_eq_way = {T_2541,T_2540};
  assign T_2542 = s1_tag_eq_way[0];
  assign T_2543 = meta_io_resp_0_coh_state != 2'h0;
  assign T_2544 = T_2542 & T_2543;
  assign T_2545 = s1_tag_eq_way[1];
  assign T_2546 = meta_io_resp_1_coh_state != 2'h0;
  assign T_2547 = T_2545 & T_2546;
  assign T_2548 = s1_tag_eq_way[2];
  assign T_2549 = meta_io_resp_2_coh_state != 2'h0;
  assign T_2550 = T_2548 & T_2549;
  assign T_2551 = s1_tag_eq_way[3];
  assign T_2552 = meta_io_resp_3_coh_state != 2'h0;
  assign T_2553 = T_2551 & T_2552;
  assign T_2559_0 = T_2544;
  assign T_2559_1 = T_2547;
  assign T_2559_2 = T_2550;
  assign T_2559_3 = T_2553;
  assign T_2561 = {T_2559_1,T_2559_0};
  assign T_2562 = {T_2559_3,T_2559_2};
  assign s1_tag_match_way = {T_2562,T_2561};
  assign T_2564 = s1_valid == 1'h0;
  assign GEN_34 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s2_tag_match = s2_tag_match_way != 4'h0;
  assign GEN_35 = s1_clk_en ? meta_io_resp_0_coh_state : T_2569_state;
  assign GEN_36 = s1_clk_en ? meta_io_resp_1_coh_state : T_2591_state;
  assign GEN_37 = s1_clk_en ? meta_io_resp_2_coh_state : T_2613_state;
  assign GEN_38 = s1_clk_en ? meta_io_resp_3_coh_state : T_2635_state;
  assign T_2830_0_state = T_2569_state;
  assign T_2830_1_state = T_2591_state;
  assign T_2830_2_state = T_2613_state;
  assign T_2830_3_state = T_2635_state;
  assign T_2937 = s2_tag_match_way[0];
  assign T_2938 = s2_tag_match_way[1];
  assign T_2939 = s2_tag_match_way[2];
  assign T_2940 = s2_tag_match_way[3];
  assign T_2942 = T_2937 ? T_2830_0_state : 2'h0;
  assign T_2944 = T_2938 ? T_2830_1_state : 2'h0;
  assign T_2946 = T_2939 ? T_2830_2_state : 2'h0;
  assign T_2948 = T_2940 ? T_2830_3_state : 2'h0;
  assign T_2971 = T_2942 | T_2944;
  assign T_2972 = T_2971 | T_2946;
  assign T_2973 = T_2972 | T_2948;
  assign s2_hit_state_state = T_2973;
  assign T_3018 = s2_req_cmd == 5'h1;
  assign T_3019 = s2_req_cmd == 5'h7;
  assign T_3020 = T_3018 | T_3019;
  assign T_3021 = s2_req_cmd[3];
  assign T_3022 = s2_req_cmd == 5'h4;
  assign T_3023 = T_3021 | T_3022;
  assign T_3024 = T_3020 | T_3023;
  assign T_3025 = s2_req_cmd == 5'h3;
  assign T_3026 = T_3024 | T_3025;
  assign T_3027 = s2_req_cmd == 5'h6;
  assign T_3028 = T_3026 | T_3027;
  assign T_3029 = s2_hit_state_state == 2'h1;
  assign T_3030 = s2_hit_state_state == 2'h2;
  assign T_3031 = T_3029 | T_3030;
  assign T_3035 = T_3028 ? T_3031 : T_3031;
  assign T_3036 = s2_tag_match & T_3035;
  assign T_3044 = T_3024 ? 2'h2 : s2_hit_state_state;
  assign T_3067_state = T_3044;
  assign T_3089 = s2_hit_state_state == T_3067_state;
  assign s2_hit = T_3036 & T_3089;
  assign lrsc_valid = lrsc_count != 5'h0;
  assign T_3094 = lrsc_addr == T_2522;
  assign s2_lrsc_addr_match = lrsc_valid & T_3094;
  assign T_3096 = s2_lrsc_addr_match == 1'h0;
  assign s2_sc_fail = T_3019 & T_3096;
  assign T_3098 = lrsc_count - 5'h1;
  assign T_3099 = T_3098[4:0];
  assign GEN_39 = lrsc_valid ? T_3099 : lrsc_count;
  assign T_3100 = s2_valid_masked & s2_hit;
  assign T_3101 = T_3100 | s2_replay;
  assign T_3103 = lrsc_valid == 1'h0;
  assign GEN_40 = T_3103 ? 5'h1f : GEN_39;
  assign GEN_41 = T_3027 ? GEN_40 : GEN_39;
  assign GEN_42 = T_3027 ? T_2522 : lrsc_addr;
  assign GEN_43 = T_3019 ? 5'h0 : GEN_41;
  assign GEN_44 = T_3101 ? GEN_43 : GEN_39;
  assign GEN_45 = T_3101 ? GEN_42 : lrsc_addr;
  assign GEN_46 = io_cpu_invalidate_lr ? 5'h0 : GEN_44;
  assign s2_data_0 = T_3121_0;
  assign s2_data_1 = T_3139_0;
  assign s2_data_2 = T_3157_0;
  assign s2_data_3 = T_3175_0;
  assign T_3124 = s1_clk_en & T_2542;
  assign T_3132 = data_io_resp_0;
  assign GEN_47 = T_3124 ? T_3132 : T_3121_0;
  assign T_3142 = s1_clk_en & T_2545;
  assign T_3150 = data_io_resp_1;
  assign GEN_48 = T_3142 ? T_3150 : T_3139_0;
  assign T_3160 = s1_clk_en & T_2548;
  assign T_3168 = data_io_resp_2;
  assign GEN_49 = T_3160 ? T_3168 : T_3157_0;
  assign T_3178 = s1_clk_en & T_2551;
  assign T_3186 = data_io_resp_3;
  assign GEN_50 = T_3178 ? T_3186 : T_3175_0;
  assign T_3192 = T_2937 ? s2_data_0 : 64'h0;
  assign T_3194 = T_2938 ? s2_data_1 : 64'h0;
  assign T_3196 = T_2939 ? s2_data_2 : 64'h0;
  assign T_3198 = T_2940 ? s2_data_3 : 64'h0;
  assign T_3200 = T_3192 | T_3194;
  assign T_3201 = T_3200 | T_3196;
  assign T_3202 = T_3201 | T_3198;
  assign s2_data_muxed = T_3202;
  assign T_3204 = 1'h0 >> 1'h0;
  assign T_3208 = s2_sc_fail == 1'h0;
  assign T_3209 = T_3101 & T_3208;
  assign T_3217 = T_3209 & T_3024;
  assign amoalu_clk = clk;
  assign amoalu_reset = reset;
  assign amoalu_io_addr = s2_req_addr[2:0];
  assign amoalu_io_cmd = s2_req_cmd;
  assign amoalu_io_typ = s2_req_typ[1:0];
  assign amoalu_io_lhs = s2_data_word;
  assign amoalu_io_rhs = s2_req_data;
  assign T_3218 = s2_valid | s2_replay;
  assign T_3226 = T_3024 | T_3204;
  assign T_3227 = T_3218 & T_3226;
  assign T_3228 = T_3204 ? s2_data_muxed : amoalu_io_out;
  assign GEN_51 = T_3227 ? s2_req_addr : s3_req_addr;
  assign GEN_52 = T_3227 ? s2_req_tag : s3_req_tag;
  assign GEN_53 = T_3227 ? s2_req_cmd : s3_req_cmd;
  assign GEN_54 = T_3227 ? s2_req_typ : s3_req_typ;
  assign GEN_55 = T_3227 ? s2_req_phys : s3_req_phys;
  assign GEN_56 = T_3227 ? T_3228 : s3_req_data;
  assign GEN_57 = T_3227 ? s2_tag_match_way : s3_way;
  assign T_3231 = 2'h1 << 1'h0;
  assign T_3233 = T_5231;
  assign T_3237 = T_3236[0];
  assign T_3238 = T_3236[2];
  assign T_3239 = T_3237 ^ T_3238;
  assign T_3240 = T_3236[3];
  assign T_3241 = T_3239 ^ T_3240;
  assign T_3242 = T_3236[5];
  assign T_3243 = T_3241 ^ T_3242;
  assign T_3244 = T_3236[15:1];
  assign T_3245 = {T_3243,T_3244};
  assign GEN_58 = T_3233 ? T_3245 : T_3236;
  assign T_3246 = T_3236[1:0];
  assign s1_replaced_way_en = 4'h1 << T_3246;
  assign GEN_59 = s1_clk_en ? T_3246 : T_3249;
  assign s2_replaced_way_en = 4'h1 << T_3249;
  assign T_3251 = s1_replaced_way_en[0];
  assign T_3252 = s1_clk_en & T_3251;
  assign GEN_60 = T_3252 ? meta_io_resp_0_tag : T_3253_tag;
  assign GEN_61 = T_3252 ? meta_io_resp_0_coh_state : T_3253_coh_state;
  assign T_3337 = s1_replaced_way_en[1];
  assign T_3338 = s1_clk_en & T_3337;
  assign GEN_62 = T_3338 ? meta_io_resp_1_tag : T_3339_tag;
  assign GEN_63 = T_3338 ? meta_io_resp_1_coh_state : T_3339_coh_state;
  assign T_3423 = s1_replaced_way_en[2];
  assign T_3424 = s1_clk_en & T_3423;
  assign GEN_64 = T_3424 ? meta_io_resp_2_tag : T_3425_tag;
  assign GEN_65 = T_3424 ? meta_io_resp_2_coh_state : T_3425_coh_state;
  assign T_3509 = s1_replaced_way_en[3];
  assign T_3510 = s1_clk_en & T_3509;
  assign GEN_66 = T_3510 ? meta_io_resp_3_tag : T_3511_tag;
  assign GEN_67 = T_3510 ? meta_io_resp_3_coh_state : T_3511_coh_state;
  assign T_4264_0_tag = T_3253_tag;
  assign T_4264_0_coh_state = T_3253_coh_state;
  assign T_4264_1_tag = T_3339_tag;
  assign T_4264_1_coh_state = T_3339_coh_state;
  assign T_4264_2_tag = T_3425_tag;
  assign T_4264_2_coh_state = T_3425_coh_state;
  assign T_4264_3_tag = T_3511_tag;
  assign T_4264_3_coh_state = T_3511_coh_state;
  assign T_4681 = s2_replaced_way_en[0];
  assign T_4682 = s2_replaced_way_en[1];
  assign T_4683 = s2_replaced_way_en[2];
  assign T_4684 = s2_replaced_way_en[3];
  assign T_4685 = {T_4264_0_tag,T_4264_0_coh_state};
  assign T_4687 = T_4681 ? T_4685 : 22'h0;
  assign T_4688 = {T_4264_1_tag,T_4264_1_coh_state};
  assign T_4690 = T_4682 ? T_4688 : 22'h0;
  assign T_4691 = {T_4264_2_tag,T_4264_2_coh_state};
  assign T_4693 = T_4683 ? T_4691 : 22'h0;
  assign T_4694 = {T_4264_3_tag,T_4264_3_coh_state};
  assign T_4696 = T_4684 ? T_4694 : 22'h0;
  assign T_4781 = T_4687 | T_4690;
  assign T_4782 = T_4781 | T_4693;
  assign T_4783 = T_4782 | T_4696;
  assign s2_repl_meta_tag = T_4952;
  assign s2_repl_meta_coh_state = T_4951;
  assign T_4951 = T_4783[1:0];
  assign T_4952 = T_4783[21:2];
  assign T_4954 = s2_hit == 1'h0;
  assign T_4955 = s2_valid_masked & T_4954;
  assign T_4956 = s2_req_cmd == 5'h2;
  assign T_4958 = T_4956 | T_3025;
  assign T_4959 = s2_req_cmd == 5'h0;
  assign T_4961 = T_4959 | T_3027;
  assign T_4963 = T_4961 | T_3019;
  assign T_4967 = T_4963 | T_3023;
  assign T_4968 = T_4958 | T_4967;
  assign T_4976 = T_4968 | T_3024;
  assign T_4977 = T_4955 & T_4976;
  assign T_5062_tag = s2_repl_meta_tag;
  assign T_5062_coh_state = s2_hit_state_state;
  assign T_5146_tag = s2_tag_match ? T_5062_tag : s2_repl_meta_tag;
  assign T_5146_coh_state = s2_tag_match ? T_5062_coh_state : s2_repl_meta_coh_state;
  assign T_5230 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign T_5231 = mshrs_io_req_ready & mshrs_io_req_valid;
  assign T_5235 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign releaseArb_clk = clk;
  assign releaseArb_reset = reset;
  assign releaseArb_io_in_0_valid = wb_io_release_valid;
  assign releaseArb_io_in_0_bits_addr_beat = wb_io_release_bits_addr_beat;
  assign releaseArb_io_in_0_bits_addr_block = wb_io_release_bits_addr_block;
  assign releaseArb_io_in_0_bits_client_xact_id = wb_io_release_bits_client_xact_id;
  assign releaseArb_io_in_0_bits_voluntary = wb_io_release_bits_voluntary;
  assign releaseArb_io_in_0_bits_r_type = wb_io_release_bits_r_type;
  assign releaseArb_io_in_0_bits_data = wb_io_release_bits_data;
  assign releaseArb_io_in_1_valid = prober_io_rep_valid;
  assign releaseArb_io_in_1_bits_addr_beat = prober_io_rep_bits_addr_beat;
  assign releaseArb_io_in_1_bits_addr_block = prober_io_rep_bits_addr_block;
  assign releaseArb_io_in_1_bits_client_xact_id = prober_io_rep_bits_client_xact_id;
  assign releaseArb_io_in_1_bits_voluntary = prober_io_rep_bits_voluntary;
  assign releaseArb_io_in_1_bits_r_type = prober_io_rep_bits_r_type;
  assign releaseArb_io_in_1_bits_data = prober_io_rep_bits_data;
  assign releaseArb_io_out_ready = io_mem_release_ready;
  assign T_5265 = io_mem_probe_valid & T_3103;
  assign T_5268 = prober_io_req_ready & T_3103;
  assign FlowThroughSerializer_1_1_clk = clk;
  assign FlowThroughSerializer_1_1_reset = reset;
  assign FlowThroughSerializer_1_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_1_io_in_bits_manager_id = io_mem_grant_bits_manager_id;
  assign FlowThroughSerializer_1_1_io_out_ready = T_5286;
  assign T_5269 = FlowThroughSerializer_1_1_io_out_ready & FlowThroughSerializer_1_1_io_out_valid;
  assign T_5277_0 = 3'h5;
  assign T_5277_1 = 3'h4;
  assign GEN_86 = {{1'd0}, T_5277_0};
  assign T_5279 = FlowThroughSerializer_1_1_io_out_bits_g_type == GEN_86;
  assign GEN_87 = {{1'd0}, T_5277_1};
  assign T_5280 = FlowThroughSerializer_1_1_io_out_bits_g_type == GEN_87;
  assign T_5281 = T_5279 | T_5280;
  assign T_5282 = FlowThroughSerializer_1_1_io_out_bits_g_type == 4'h0;
  assign T_5283 = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type ? T_5281 : T_5282;
  assign T_5285 = T_5283 == 1'h0;
  assign T_5286 = writeArb_io_in_1_ready | T_5285;
  assign T_5294_0 = 3'h5;
  assign T_5294_1 = 3'h4;
  assign GEN_88 = {{1'd0}, T_5294_0};
  assign T_5296 = FlowThroughSerializer_1_1_io_out_bits_g_type == GEN_88;
  assign GEN_89 = {{1'd0}, T_5294_1};
  assign T_5297 = FlowThroughSerializer_1_1_io_out_bits_g_type == GEN_89;
  assign T_5298 = T_5296 | T_5297;
  assign T_5300 = FlowThroughSerializer_1_1_io_out_bits_is_builtin_type ? T_5298 : T_5282;
  assign T_5301 = FlowThroughSerializer_1_1_io_out_valid & T_5300;
  assign T_5303 = FlowThroughSerializer_1_1_io_out_bits_client_xact_id < 2'h2;
  assign T_5304 = T_5301 & T_5303;
  assign T_5307 = FlowThroughSerializer_1_1_io_out_bits_data;
  assign T_5309 = FlowThroughSerializer_1_1_io_out_valid == 1'h0;
  assign T_5310 = T_5309 | FlowThroughSerializer_1_1_io_out_ready;
  assign wbArb_clk = clk;
  assign wbArb_reset = reset;
  assign wbArb_io_in_0_valid = prober_io_wb_req_valid;
  assign wbArb_io_in_0_bits_addr_beat = prober_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_0_bits_addr_block = prober_io_wb_req_bits_addr_block;
  assign wbArb_io_in_0_bits_client_xact_id = prober_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_0_bits_voluntary = prober_io_wb_req_bits_voluntary;
  assign wbArb_io_in_0_bits_r_type = prober_io_wb_req_bits_r_type;
  assign wbArb_io_in_0_bits_data = prober_io_wb_req_bits_data;
  assign wbArb_io_in_0_bits_way_en = prober_io_wb_req_bits_way_en;
  assign wbArb_io_in_1_valid = mshrs_io_wb_req_valid;
  assign wbArb_io_in_1_bits_addr_beat = mshrs_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_1_bits_addr_block = mshrs_io_wb_req_bits_addr_block;
  assign wbArb_io_in_1_bits_client_xact_id = mshrs_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_1_bits_voluntary = mshrs_io_wb_req_bits_voluntary;
  assign wbArb_io_in_1_bits_r_type = mshrs_io_wb_req_bits_r_type;
  assign wbArb_io_in_1_bits_data = mshrs_io_wb_req_bits_data;
  assign wbArb_io_in_1_bits_way_en = mshrs_io_wb_req_bits_way_en;
  assign wbArb_io_out_ready = wb_io_req_ready;
  assign T_5360 = s3_valid & metaReadArb_io_out_valid;
  assign GEN_69 = T_5360 ? s3_req_addr : s4_req_addr;
  assign GEN_70 = T_5360 ? s3_req_tag : s4_req_tag;
  assign GEN_71 = T_5360 ? s3_req_cmd : s4_req_cmd;
  assign GEN_72 = T_5360 ? s3_req_typ : s4_req_typ;
  assign GEN_73 = T_5360 ? s3_req_phys : s4_req_phys;
  assign GEN_74 = T_5360 ? s3_req_data : s4_req_data;
  assign T_5427 = s2_valid_masked | s2_replay;
  assign T_5430 = T_5427 & T_3208;
  assign T_5431 = s1_addr[31:3];
  assign T_5432 = s2_req_addr[39:3];
  assign GEN_90 = {{8'd0}, T_5431};
  assign T_5433 = GEN_90 == T_5432;
  assign T_5434 = T_5430 & T_5433;
  assign T_5442 = T_5434 & T_3024;
  assign T_5444 = s3_req_addr[39:3];
  assign T_5445 = GEN_90 == T_5444;
  assign T_5446 = s3_valid & T_5445;
  assign T_5447 = s3_req_cmd == 5'h1;
  assign T_5448 = s3_req_cmd == 5'h7;
  assign T_5449 = T_5447 | T_5448;
  assign T_5450 = s3_req_cmd[3];
  assign T_5451 = s3_req_cmd == 5'h4;
  assign T_5452 = T_5450 | T_5451;
  assign T_5453 = T_5449 | T_5452;
  assign T_5454 = T_5446 & T_5453;
  assign T_5456 = s4_req_addr[39:3];
  assign T_5457 = GEN_90 == T_5456;
  assign T_5458 = s4_valid & T_5457;
  assign T_5459 = s4_req_cmd == 5'h1;
  assign T_5460 = s4_req_cmd == 5'h7;
  assign T_5461 = T_5459 | T_5460;
  assign T_5462 = s4_req_cmd[3];
  assign T_5463 = s4_req_cmd == 5'h4;
  assign T_5464 = T_5462 | T_5463;
  assign T_5465 = T_5461 | T_5464;
  assign T_5466 = T_5458 & T_5465;
  assign T_5470 = T_5442 | T_5454;
  assign T_5471 = T_5470 | T_5466;
  assign T_5472 = T_5454 ? s3_req_data : s4_req_data;
  assign T_5473 = T_5442 ? amoalu_io_out : T_5472;
  assign GEN_75 = T_5471 ? T_5473 : s2_store_bypass_data;
  assign GEN_77 = s1_clk_en ? T_5471 : s2_store_bypass;
  assign GEN_78 = s1_clk_en ? GEN_75 : s2_store_bypass_data;
  assign s2_data_word_prebypass = s2_data_muxed >> 7'h0;
  assign s2_data_word = s2_store_bypass ? s2_store_bypass_data : s2_data_word_prebypass;
  assign T_5477 = s2_req_typ[2];
  assign T_5479 = T_5477 == 1'h0;
  assign T_5480 = s2_req_typ[1:0];
  assign T_5481 = dtlb_io_req_valid & dtlb_io_resp_miss;
  assign T_5482 = s1_req_addr[11:6];
  assign T_5483 = T_5482 == prober_io_meta_write_bits_idx;
  assign T_5485 = prober_io_req_ready == 1'h0;
  assign T_5486 = T_5483 & T_5485;
  assign s1_nack = T_5481 | T_5486;
  assign T_5487 = s1_valid | s1_replay;
  assign GEN_79 = T_5487 ? s1_nack : s2_nack_hit;
  assign GEN_80 = s2_nack_hit ? 1'h0 : T_4977;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T_5492 = mshrs_io_req_ready == 1'h0;
  assign s2_nack_miss = T_4954 & T_5492;
  assign T_5493 = s2_nack_hit | s2_nack_victim;
  assign s2_nack = T_5493 | s2_nack_miss;
  assign T_5495 = s2_nack == 1'h0;
  assign T_5496 = s2_valid & T_5495;
  assign T_5498 = T_3218 & s2_hit;
  assign s2_recycle_ecc = T_5498 & T_3204;
  assign GEN_81 = T_5487 ? s2_recycle_ecc : s2_recycle_next;
  assign T_5501 = s2_recycle_ecc | s2_recycle_next;
  assign T_5503 = s2_valid | block_miss;
  assign T_5504 = T_5503 & s2_nack_miss;
  assign GEN_82 = block_miss ? 1'h0 : GEN_33;
  assign cache_resp_valid = T_5863;
  assign cache_resp_bits_addr = s2_req_addr;
  assign cache_resp_bits_tag = s2_req_tag;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign cache_resp_bits_typ = s2_req_typ;
  assign cache_resp_bits_data = T_5933;
  assign cache_resp_bits_replay = s2_replay;
  assign cache_resp_bits_has_data = T_4967;
  assign cache_resp_bits_data_word_bypass = GEN_92;
  assign cache_resp_bits_store_data = s2_req_data;
  assign T_5860 = s2_replay | T_3100;
  assign T_5862 = T_3204 == 1'h0;
  assign T_5863 = T_5860 & T_5862;
  assign T_5873 = s2_req_addr[2];
  assign T_5874 = s2_data_word[63:32];
  assign T_5875 = s2_data_word[31:0];
  assign T_5876 = T_5873 ? T_5874 : T_5875;
  assign T_5882 = T_5480 == 2'h2;
  assign T_5884 = T_5876[31];
  assign T_5885 = T_5479 & T_5884;
  assign T_5889 = T_5885 ? 32'hffffffff : 32'h0;
  assign T_5891 = T_5882 ? T_5889 : T_5874;
  assign T_5892 = {T_5891,T_5876};
  assign T_5893 = s2_req_addr[1];
  assign T_5894 = T_5892[31:16];
  assign T_5895 = T_5892[15:0];
  assign T_5896 = T_5893 ? T_5894 : T_5895;
  assign T_5902 = T_5480 == 2'h1;
  assign T_5904 = T_5896[15];
  assign T_5905 = T_5479 & T_5904;
  assign T_5909 = T_5905 ? 48'hffffffffffff : 48'h0;
  assign T_5910 = T_5892[63:16];
  assign T_5911 = T_5902 ? T_5909 : T_5910;
  assign T_5912 = {T_5911,T_5896};
  assign T_5913 = s2_req_addr[0];
  assign T_5914 = T_5912[15:8];
  assign T_5915 = T_5912[7:0];
  assign T_5916 = T_5913 ? T_5914 : T_5915;
  assign T_5920 = T_3019 ? 8'h0 : T_5916;
  assign T_5922 = T_5480 == 2'h0;
  assign T_5923 = T_5922 | T_3019;
  assign T_5924 = T_5920[7];
  assign T_5925 = T_5479 & T_5924;
  assign T_5929 = T_5925 ? 56'hffffffffffffff : 56'h0;
  assign T_5930 = T_5912[63:8];
  assign T_5931 = T_5923 ? T_5929 : T_5930;
  assign T_5932 = {T_5931,T_5920};
  assign GEN_93 = {{63'd0}, s2_sc_fail};
  assign T_5933 = T_5932 | GEN_93;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign uncache_resp_bits_data_word_bypass = mshrs_io_resp_bits_data_word_bypass;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign T_6289 = T_5487 == 1'h0;
  assign T_6291 = s2_valid & s2_nack;
  assign T_6292_valid = mshrs_io_resp_ready ? uncache_resp_valid : cache_resp_valid;
  assign T_6292_bits_addr = mshrs_io_resp_ready ? uncache_resp_bits_addr : cache_resp_bits_addr;
  assign T_6292_bits_tag = mshrs_io_resp_ready ? uncache_resp_bits_tag : cache_resp_bits_tag;
  assign T_6292_bits_cmd = mshrs_io_resp_ready ? uncache_resp_bits_cmd : cache_resp_bits_cmd;
  assign T_6292_bits_typ = mshrs_io_resp_ready ? uncache_resp_bits_typ : cache_resp_bits_typ;
  assign T_6292_bits_data = mshrs_io_resp_ready ? uncache_resp_bits_data : cache_resp_bits_data;
  assign T_6292_bits_replay = mshrs_io_resp_ready ? uncache_resp_bits_replay : cache_resp_bits_replay;
  assign T_6292_bits_has_data = mshrs_io_resp_ready ? uncache_resp_bits_has_data : cache_resp_bits_has_data;
  assign T_6292_bits_store_data = mshrs_io_resp_ready ? uncache_resp_bits_store_data : cache_resp_bits_store_data;
  assign T_6456 = mshrs_io_fence_rdy & T_2564;
  assign T_6458 = s2_valid == 1'h0;
  assign T_6459 = T_6456 & T_6458;
  assign T_6460 = s1_replay & s1_read;
  assign T_6461 = T_6460 | mshrs_io_replay_next;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_154[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_76 = GEN_155[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_91 = GEN_156[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_92 = GEN_157[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {1{$random}};
  s1_valid = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  s1_req_addr = GEN_95[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {1{$random}};
  s1_req_tag = GEN_96[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  s1_req_cmd = GEN_97[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  s1_req_typ = GEN_98[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  s1_req_phys = GEN_99[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {2{$random}};
  s1_req_data = GEN_100[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  s1_replay = GEN_101[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  s1_clk_en = GEN_102[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  s2_valid = GEN_103[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {2{$random}};
  s2_req_addr = GEN_104[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  s2_req_tag = GEN_105[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  s2_req_cmd = GEN_106[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  s2_req_typ = GEN_107[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  s2_req_phys = GEN_108[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {2{$random}};
  s2_req_data = GEN_109[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2049 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  s3_valid = GEN_111[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {2{$random}};
  s3_req_addr = GEN_112[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  s3_req_tag = GEN_113[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  s3_req_cmd = GEN_114[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  s3_req_typ = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  s3_req_phys = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {2{$random}};
  s3_req_data = GEN_117[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  s3_way = GEN_118[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  s1_recycled = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  s2_tag_match_way = GEN_120[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {1{$random}};
  T_2569_state = GEN_121[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_122 = {1{$random}};
  T_2591_state = GEN_122[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_123 = {1{$random}};
  T_2613_state = GEN_123[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_124 = {1{$random}};
  T_2635_state = GEN_124[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  lrsc_count = GEN_125[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {2{$random}};
  lrsc_addr = GEN_126[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {2{$random}};
  T_3121_0 = GEN_127[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {2{$random}};
  T_3139_0 = GEN_128[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {2{$random}};
  T_3157_0 = GEN_129[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {2{$random}};
  T_3175_0 = GEN_130[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  T_3236 = GEN_131[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  T_3249 = GEN_132[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  T_3253_tag = GEN_133[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  T_3253_coh_state = GEN_134[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  T_3339_tag = GEN_135[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {1{$random}};
  T_3339_coh_state = GEN_136[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  T_3425_tag = GEN_137[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  T_3425_coh_state = GEN_138[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  T_3511_tag = GEN_139[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  T_3511_coh_state = GEN_140[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  s4_valid = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {2{$random}};
  s4_req_addr = GEN_142[39:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  s4_req_tag = GEN_143[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  s4_req_cmd = GEN_144[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  s4_req_typ = GEN_145[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  s4_req_phys = GEN_146[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {2{$random}};
  s4_req_data = GEN_147[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {2{$random}};
  s2_store_bypass_data = GEN_148[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  s2_store_bypass = GEN_149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  s2_nack_hit = GEN_150[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  s2_recycle_next = GEN_151[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  block_miss = GEN_152[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  T_6290 = GEN_153[0:0];
  `endif
  GEN_154 = {1{$random}};
  GEN_155 = {1{$random}};
  GEN_156 = {1{$random}};
  GEN_157 = {2{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_1901;
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_addr <= s2_req_addr;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_addr <= mshrs_io_replay_bits_addr;
        end else begin
          if(prober_io_meta_read_valid) begin
            s1_req_addr <= {{8'd0}, T_2153};
          end else begin
            if(wb_io_meta_read_valid) begin
              s1_req_addr <= {{8'd0}, T_2150};
            end else begin
              if(io_cpu_req_valid) begin
                s1_req_addr <= io_cpu_req_bits_addr;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_tag <= s2_req_tag;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_tag <= mshrs_io_replay_bits_tag;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_tag <= io_cpu_req_bits_tag;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_cmd <= s2_req_cmd;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_cmd <= mshrs_io_replay_bits_cmd;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_cmd <= io_cpu_req_bits_cmd;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_typ <= s2_req_typ;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_typ <= mshrs_io_replay_bits_typ;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_typ <= io_cpu_req_bits_typ;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_phys <= s2_req_phys;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_phys <= mshrs_io_replay_bits_phys;
        end else begin
          if(prober_io_meta_read_valid) begin
            s1_req_phys <= 1'h1;
          end else begin
            if(wb_io_meta_read_valid) begin
              s1_req_phys <= 1'h1;
            end else begin
              if(io_cpu_req_valid) begin
                s1_req_phys <= io_cpu_req_bits_phys;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s2_recycle) begin
        s1_req_data <= s2_req_data;
      end else begin
        if(mshrs_io_replay_valid) begin
          s1_req_data <= mshrs_io_replay_bits_data;
        end else begin
          if(io_cpu_req_valid) begin
            s1_req_data <= io_cpu_req_bits_data;
          end
        end
      end
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T_5235;
    end
    if(1'h0) begin
    end else begin
      s1_clk_en <= metaReadArb_io_out_valid;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_addr <= {{8'd0}, s1_addr};
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_tag <= s1_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_req_phys <= s1_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        if(s1_recycled) begin
          s2_req_data <= s1_req_data;
        end else begin
          if(s1_write) begin
            if(s1_replay) begin
              s2_req_data <= mshrs_io_replay_bits_data;
            end else begin
              s2_req_data <= io_cpu_s1_data;
            end
          end
        end
      end
    end
    if(reset) begin
      T_2049 <= 1'h0;
    end else begin
      T_2049 <= s1_replay;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T_3217;
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_req_addr <= s2_req_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_req_tag <= s2_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_req_cmd <= s2_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_req_typ <= s2_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_req_phys <= s2_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        if(T_3204) begin
          s3_req_data <= s2_data_muxed;
        end else begin
          s3_req_data <= amoalu_io_out;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3227) begin
        s3_way <= s2_tag_match_way;
      end
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else begin
      if(s1_clk_en) begin
        s1_recycled <= s2_recycle;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_tag_match_way <= s1_tag_match_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2569_state <= meta_io_resp_0_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2591_state <= meta_io_resp_1_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2613_state <= meta_io_resp_2_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_2635_state <= meta_io_resp_3_coh_state;
      end
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else begin
      if(io_cpu_invalidate_lr) begin
        lrsc_count <= 5'h0;
      end else begin
        if(T_3101) begin
          if(T_3019) begin
            lrsc_count <= 5'h0;
          end else begin
            if(T_3027) begin
              if(T_3103) begin
                lrsc_count <= 5'h1f;
              end else begin
                if(lrsc_valid) begin
                  lrsc_count <= T_3099;
                end
              end
            end else begin
              if(lrsc_valid) begin
                lrsc_count <= T_3099;
              end
            end
          end
        end else begin
          if(lrsc_valid) begin
            lrsc_count <= T_3099;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3101) begin
        if(T_3027) begin
          lrsc_addr <= T_2522;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3124) begin
        T_3121_0 <= T_3132;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3142) begin
        T_3139_0 <= T_3150;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3160) begin
        T_3157_0 <= T_3168;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3178) begin
        T_3175_0 <= T_3186;
      end
    end
    if(reset) begin
      T_3236 <= 16'h1;
    end else begin
      if(T_3233) begin
        T_3236 <= T_3245;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        T_3249 <= T_3246;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3252) begin
        T_3253_tag <= meta_io_resp_0_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3252) begin
        T_3253_coh_state <= meta_io_resp_0_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3338) begin
        T_3339_tag <= meta_io_resp_1_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3338) begin
        T_3339_coh_state <= meta_io_resp_1_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3424) begin
        T_3425_tag <= meta_io_resp_2_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3424) begin
        T_3425_coh_state <= meta_io_resp_2_coh_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3510) begin
        T_3511_tag <= meta_io_resp_3_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_3510) begin
        T_3511_coh_state <= meta_io_resp_3_coh_state;
      end
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_addr <= s3_req_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_tag <= s3_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_cmd <= s3_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_typ <= s3_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_phys <= s3_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5360) begin
        s4_req_data <= s3_req_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        if(T_5471) begin
          if(T_5442) begin
            s2_store_bypass_data <= amoalu_io_out;
          end else begin
            if(T_5454) begin
              s2_store_bypass_data <= s3_req_data;
            end else begin
              s2_store_bypass_data <= s4_req_data;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_clk_en) begin
        s2_store_bypass <= T_5471;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5487) begin
        s2_nack_hit <= s1_nack;
      end
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else begin
      if(T_5487) begin
        s2_recycle_next <= s2_recycle_ecc;
      end
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T_5504;
    end
    if(1'h0) begin
    end else begin
      T_6290 <= T_6289;
    end
  end
endmodule
module FPUDecoder(
  input   clk,
  input   reset,
  input  [31:0] io_inst,
  output [4:0] io_sigs_cmd,
  output  io_sigs_ldst,
  output  io_sigs_wen,
  output  io_sigs_ren1,
  output  io_sigs_ren2,
  output  io_sigs_ren3,
  output  io_sigs_swap12,
  output  io_sigs_swap23,
  output  io_sigs_single,
  output  io_sigs_fromint,
  output  io_sigs_toint,
  output  io_sigs_fastpipe,
  output  io_sigs_fma,
  output  io_sigs_div,
  output  io_sigs_sqrt,
  output  io_sigs_round,
  output  io_sigs_wflags
);
  wire [31:0] T_20;
  wire  T_22;
  wire [31:0] T_24;
  wire  T_26;
  wire  T_29;
  wire [31:0] T_31;
  wire  T_33;
  wire [31:0] T_35;
  wire  T_37;
  wire  T_40;
  wire [31:0] T_42;
  wire  T_44;
  wire [31:0] T_46;
  wire  T_48;
  wire  T_51;
  wire [31:0] T_53;
  wire  T_55;
  wire  T_58;
  wire [31:0] T_60;
  wire  T_62;
  wire [1:0] T_65;
  wire [1:0] T_66;
  wire [2:0] T_67;
  wire [4:0] decoder_0;
  wire [31:0] T_70;
  wire  T_72;
  wire [31:0] T_74;
  wire  T_76;
  wire [31:0] T_78;
  wire  T_80;
  wire  T_83;
  wire  decoder_2;
  wire [31:0] T_85;
  wire  T_87;
  wire [31:0] T_89;
  wire  T_91;
  wire [31:0] T_93;
  wire  T_95;
  wire  T_98;
  wire  decoder_3;
  wire [31:0] T_100;
  wire  T_102;
  wire [31:0] T_104;
  wire  T_106;
  wire  T_109;
  wire  decoder_4;
  wire [31:0] T_112;
  wire  T_114;
  wire  decoder_6;
  wire [31:0] T_118;
  wire  T_120;
  wire [31:0] T_123;
  wire  T_125;
  wire [31:0] T_127;
  wire  T_129;
  wire  decoder_8;
  wire [31:0] T_133;
  wire  T_135;
  wire  T_140;
  wire  decoder_10;
  wire [31:0] T_144;
  wire  T_146;
  wire [31:0] T_148;
  wire  T_150;
  wire  decoder_11;
  wire [31:0] T_154;
  wire  T_156;
  wire [31:0] T_158;
  wire  T_160;
  wire  T_163;
  wire  decoder_12;
  wire [31:0] T_165;
  wire  T_167;
  wire  T_172;
  wire [31:0] T_175;
  wire  T_177;
  wire [31:0] T_179;
  wire  T_181;
  wire  T_184;
  wire  decoder_15;
  wire [31:0] T_186;
  wire  T_188;
  wire [31:0] T_190;
  wire  T_192;
  wire  T_196;
  wire  decoder_16;
  assign io_sigs_cmd = decoder_0;
  assign io_sigs_ldst = T_44;
  assign io_sigs_wen = decoder_2;
  assign io_sigs_ren1 = decoder_3;
  assign io_sigs_ren2 = decoder_4;
  assign io_sigs_ren3 = T_95;
  assign io_sigs_swap12 = decoder_6;
  assign io_sigs_swap23 = T_120;
  assign io_sigs_single = decoder_8;
  assign io_sigs_fromint = T_135;
  assign io_sigs_toint = decoder_10;
  assign io_sigs_fastpipe = decoder_11;
  assign io_sigs_fma = decoder_12;
  assign io_sigs_div = T_167;
  assign io_sigs_sqrt = T_172;
  assign io_sigs_round = decoder_15;
  assign io_sigs_wflags = decoder_16;
  assign T_20 = io_inst & 32'h4;
  assign T_22 = T_20 == 32'h4;
  assign T_24 = io_inst & 32'h8000010;
  assign T_26 = T_24 == 32'h8000010;
  assign T_29 = T_22 | T_26;
  assign T_31 = io_inst & 32'h8;
  assign T_33 = T_31 == 32'h8;
  assign T_35 = io_inst & 32'h10000010;
  assign T_37 = T_35 == 32'h10000010;
  assign T_40 = T_33 | T_37;
  assign T_42 = io_inst & 32'h40;
  assign T_44 = T_42 == 32'h0;
  assign T_46 = io_inst & 32'h20000000;
  assign T_48 = T_46 == 32'h20000000;
  assign T_51 = T_44 | T_48;
  assign T_53 = io_inst & 32'h40000000;
  assign T_55 = T_53 == 32'h40000000;
  assign T_58 = T_44 | T_55;
  assign T_60 = io_inst & 32'h10;
  assign T_62 = T_60 == 32'h0;
  assign T_65 = {T_40,T_29};
  assign T_66 = {T_62,T_58};
  assign T_67 = {T_66,T_51};
  assign decoder_0 = {T_67,T_65};
  assign T_70 = io_inst & 32'h80000020;
  assign T_72 = T_70 == 32'h0;
  assign T_74 = io_inst & 32'h30;
  assign T_76 = T_74 == 32'h0;
  assign T_78 = io_inst & 32'h10000020;
  assign T_80 = T_78 == 32'h10000000;
  assign T_83 = T_72 | T_76;
  assign decoder_2 = T_83 | T_80;
  assign T_85 = io_inst & 32'h80000004;
  assign T_87 = T_85 == 32'h0;
  assign T_89 = io_inst & 32'h10000004;
  assign T_91 = T_89 == 32'h0;
  assign T_93 = io_inst & 32'h50;
  assign T_95 = T_93 == 32'h40;
  assign T_98 = T_87 | T_91;
  assign decoder_3 = T_98 | T_95;
  assign T_100 = io_inst & 32'h40000004;
  assign T_102 = T_100 == 32'h0;
  assign T_104 = io_inst & 32'h20;
  assign T_106 = T_104 == 32'h20;
  assign T_109 = T_102 | T_106;
  assign decoder_4 = T_109 | T_95;
  assign T_112 = io_inst & 32'h50000010;
  assign T_114 = T_112 == 32'h50000010;
  assign decoder_6 = T_44 | T_114;
  assign T_118 = io_inst & 32'h30000010;
  assign T_120 = T_118 == 32'h10;
  assign T_123 = io_inst & 32'h1040;
  assign T_125 = T_123 == 32'h0;
  assign T_127 = io_inst & 32'h2000040;
  assign T_129 = T_127 == 32'h40;
  assign decoder_8 = T_125 | T_129;
  assign T_133 = io_inst & 32'h90000010;
  assign T_135 = T_133 == 32'h90000010;
  assign T_140 = T_133 == 32'h80000010;
  assign decoder_10 = T_106 | T_140;
  assign T_144 = io_inst & 32'ha0000010;
  assign T_146 = T_144 == 32'h20000010;
  assign T_148 = io_inst & 32'hd0000010;
  assign T_150 = T_148 == 32'h40000010;
  assign decoder_11 = T_146 | T_150;
  assign T_154 = io_inst & 32'h70000004;
  assign T_156 = T_154 == 32'h0;
  assign T_158 = io_inst & 32'h68000004;
  assign T_160 = T_158 == 32'h0;
  assign T_163 = T_156 | T_160;
  assign decoder_12 = T_163 | T_95;
  assign T_165 = io_inst & 32'h58000010;
  assign T_167 = T_165 == 32'h18000010;
  assign T_172 = T_148 == 32'h50000010;
  assign T_175 = io_inst & 32'h20000004;
  assign T_177 = T_175 == 32'h0;
  assign T_179 = io_inst & 32'h40002000;
  assign T_181 = T_179 == 32'h40000000;
  assign T_184 = T_177 | T_95;
  assign decoder_15 = T_184 | T_181;
  assign T_186 = io_inst & 32'h8002000;
  assign T_188 = T_186 == 32'h8000000;
  assign T_190 = io_inst & 32'hc0000004;
  assign T_192 = T_190 == 32'h80000000;
  assign T_196 = T_184 | T_188;
  assign decoder_16 = T_196 | T_192;
endmodule
module MulAddRecFN_preMul(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [1:0] io_roundingMode,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output [2:0] io_toPostMul_highExpA,
  output  io_toPostMul_isNaN_isQuietNaNA,
  output [2:0] io_toPostMul_highExpB,
  output  io_toPostMul_isNaN_isQuietNaNB,
  output  io_toPostMul_signProd,
  output  io_toPostMul_isZeroProd,
  output  io_toPostMul_opSignC,
  output [2:0] io_toPostMul_highExpC,
  output  io_toPostMul_isNaN_isQuietNaNC,
  output  io_toPostMul_isCDominant,
  output  io_toPostMul_CAlignDist_0,
  output [6:0] io_toPostMul_CAlignDist,
  output  io_toPostMul_bit0AlignedNegSigC,
  output [25:0] io_toPostMul_highAlignedNegSigC,
  output [10:0] io_toPostMul_sExpSum,
  output [1:0] io_toPostMul_roundingMode
);
  wire  signA;
  wire [8:0] expA;
  wire [22:0] fractA;
  wire [2:0] T_42;
  wire  isZeroA;
  wire  T_45;
  wire [23:0] sigA;
  wire  signB;
  wire [8:0] expB;
  wire [22:0] fractB;
  wire [2:0] T_46;
  wire  isZeroB;
  wire  T_49;
  wire [23:0] sigB;
  wire  T_50;
  wire  T_51;
  wire  opSignC;
  wire [8:0] expC;
  wire [22:0] fractC;
  wire [2:0] T_52;
  wire  isZeroC;
  wire  T_55;
  wire [23:0] sigC;
  wire  T_56;
  wire  T_57;
  wire  signProd;
  wire  isZeroProd;
  wire  T_58;
  wire  T_60;
  wire [2:0] T_64;
  wire [7:0] T_65;
  wire [10:0] T_66;
  wire [10:0] GEN_0;
  wire [11:0] T_67;
  wire [10:0] T_68;
  wire [11:0] T_70;
  wire [10:0] sExpAlignedProd;
  wire  doSubMags;
  wire [10:0] GEN_1;
  wire [11:0] T_71;
  wire [10:0] sNatCAlignDist;
  wire  T_72;
  wire  CAlignDist_floor;
  wire [9:0] T_73;
  wire  T_75;
  wire  CAlignDist_0;
  wire  T_80;
  wire  T_81;
  wire  isCDominant;
  wire  T_85;
  wire [6:0] T_86;
  wire [6:0] T_88;
  wire [6:0] CAlignDist;
  wire [10:0] sExpSum;
  wire  T_89;
  wire [5:0] T_90;
  wire [64:0] T_92;
  wire [9:0] T_93;
  wire [7:0] T_94;
  wire [3:0] T_99;
  wire [7:0] T_100;
  wire [3:0] T_101;
  wire [7:0] GEN_2;
  wire [7:0] T_102;
  wire [7:0] T_104;
  wire [7:0] T_105;
  wire [5:0] T_109;
  wire [7:0] GEN_3;
  wire [7:0] T_110;
  wire [5:0] T_111;
  wire [7:0] GEN_4;
  wire [7:0] T_112;
  wire [7:0] T_114;
  wire [7:0] T_115;
  wire [6:0] T_119;
  wire [7:0] GEN_5;
  wire [7:0] T_120;
  wire [6:0] T_121;
  wire [7:0] GEN_6;
  wire [7:0] T_122;
  wire [7:0] T_124;
  wire [7:0] T_125;
  wire [1:0] T_126;
  wire  T_127;
  wire  T_128;
  wire [1:0] T_129;
  wire [9:0] T_130;
  wire [23:0] T_132;
  wire [13:0] T_135;
  wire [7:0] T_136;
  wire [3:0] T_141;
  wire [7:0] T_142;
  wire [3:0] T_143;
  wire [7:0] GEN_7;
  wire [7:0] T_144;
  wire [7:0] T_146;
  wire [7:0] T_147;
  wire [5:0] T_151;
  wire [7:0] GEN_8;
  wire [7:0] T_152;
  wire [5:0] T_153;
  wire [7:0] GEN_9;
  wire [7:0] T_154;
  wire [7:0] T_156;
  wire [7:0] T_157;
  wire [6:0] T_161;
  wire [7:0] GEN_10;
  wire [7:0] T_162;
  wire [6:0] T_163;
  wire [7:0] GEN_11;
  wire [7:0] T_164;
  wire [7:0] T_166;
  wire [7:0] T_167;
  wire [5:0] T_168;
  wire [3:0] T_169;
  wire [1:0] T_170;
  wire  T_171;
  wire  T_172;
  wire [1:0] T_173;
  wire [1:0] T_174;
  wire  T_175;
  wire  T_176;
  wire [1:0] T_177;
  wire [3:0] T_178;
  wire [1:0] T_179;
  wire  T_180;
  wire  T_181;
  wire [1:0] T_182;
  wire [5:0] T_183;
  wire [13:0] T_184;
  wire [23:0] CExtraMask;
  wire [23:0] T_185;
  wire [23:0] negSigC;
  wire [49:0] T_189;
  wire [24:0] T_190;
  wire [74:0] T_191;
  wire [74:0] T_192;
  wire [74:0] T_193;
  wire [23:0] T_194;
  wire  T_196;
  wire  T_197;
  wire [74:0] T_198;
  wire [75:0] T_199;
  wire [74:0] alignedNegSigC;
  wire [47:0] T_200;
  wire  T_202;
  wire  T_204;
  wire  T_206;
  wire  T_207;
  wire [25:0] T_208;
  assign io_mulAddA = sigA;
  assign io_mulAddB = sigB;
  assign io_mulAddC = T_200;
  assign io_toPostMul_highExpA = T_42;
  assign io_toPostMul_isNaN_isQuietNaNA = T_202;
  assign io_toPostMul_highExpB = T_46;
  assign io_toPostMul_isNaN_isQuietNaNB = T_204;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_highExpC = T_52;
  assign io_toPostMul_isNaN_isQuietNaNC = T_206;
  assign io_toPostMul_isCDominant = isCDominant;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_bit0AlignedNegSigC = T_207;
  assign io_toPostMul_highAlignedNegSigC = T_208;
  assign io_toPostMul_sExpSum = sExpSum;
  assign io_toPostMul_roundingMode = io_roundingMode;
  assign signA = io_a[32];
  assign expA = io_a[31:23];
  assign fractA = io_a[22:0];
  assign T_42 = expA[8:6];
  assign isZeroA = T_42 == 3'h0;
  assign T_45 = isZeroA == 1'h0;
  assign sigA = {T_45,fractA};
  assign signB = io_b[32];
  assign expB = io_b[31:23];
  assign fractB = io_b[22:0];
  assign T_46 = expB[8:6];
  assign isZeroB = T_46 == 3'h0;
  assign T_49 = isZeroB == 1'h0;
  assign sigB = {T_49,fractB};
  assign T_50 = io_c[32];
  assign T_51 = io_op[0];
  assign opSignC = T_50 ^ T_51;
  assign expC = io_c[31:23];
  assign fractC = io_c[22:0];
  assign T_52 = expC[8:6];
  assign isZeroC = T_52 == 3'h0;
  assign T_55 = isZeroC == 1'h0;
  assign sigC = {T_55,fractC};
  assign T_56 = signA ^ signB;
  assign T_57 = io_op[1];
  assign signProd = T_56 ^ T_57;
  assign isZeroProd = isZeroA | isZeroB;
  assign T_58 = expB[8];
  assign T_60 = T_58 == 1'h0;
  assign T_64 = T_60 ? 3'h7 : 3'h0;
  assign T_65 = expB[7:0];
  assign T_66 = {T_64,T_65};
  assign GEN_0 = {{2'd0}, expA};
  assign T_67 = GEN_0 + T_66;
  assign T_68 = T_67[10:0];
  assign T_70 = T_68 + 11'h1b;
  assign sExpAlignedProd = T_70[10:0];
  assign doSubMags = signProd ^ opSignC;
  assign GEN_1 = {{2'd0}, expC};
  assign T_71 = sExpAlignedProd - GEN_1;
  assign sNatCAlignDist = T_71[10:0];
  assign T_72 = sNatCAlignDist[10];
  assign CAlignDist_floor = isZeroProd | T_72;
  assign T_73 = sNatCAlignDist[9:0];
  assign T_75 = T_73 == 10'h0;
  assign CAlignDist_0 = CAlignDist_floor | T_75;
  assign T_80 = T_73 < 10'h19;
  assign T_81 = CAlignDist_floor | T_80;
  assign isCDominant = T_55 & T_81;
  assign T_85 = T_73 < 10'h4a;
  assign T_86 = sNatCAlignDist[6:0];
  assign T_88 = T_85 ? T_86 : 7'h4a;
  assign CAlignDist = CAlignDist_floor ? 7'h0 : T_88;
  assign sExpSum = CAlignDist_floor ? {{2'd0}, expC} : sExpAlignedProd;
  assign T_89 = CAlignDist[6];
  assign T_90 = CAlignDist[5:0];
  assign T_92 = $signed(65'sh10000000000000000) >>> T_90;
  assign T_93 = T_92[63:54];
  assign T_94 = T_93[7:0];
  assign T_99 = T_94[7:4];
  assign T_100 = {{4'd0}, T_99};
  assign T_101 = T_94[3:0];
  assign GEN_2 = {{4'd0}, T_101};
  assign T_102 = GEN_2 << 4;
  assign T_104 = T_102 & 8'hf0;
  assign T_105 = T_100 | T_104;
  assign T_109 = T_105[7:2];
  assign GEN_3 = {{2'd0}, T_109};
  assign T_110 = GEN_3 & 8'h33;
  assign T_111 = T_105[5:0];
  assign GEN_4 = {{2'd0}, T_111};
  assign T_112 = GEN_4 << 2;
  assign T_114 = T_112 & 8'hcc;
  assign T_115 = T_110 | T_114;
  assign T_119 = T_115[7:1];
  assign GEN_5 = {{1'd0}, T_119};
  assign T_120 = GEN_5 & 8'h55;
  assign T_121 = T_115[6:0];
  assign GEN_6 = {{1'd0}, T_121};
  assign T_122 = GEN_6 << 1;
  assign T_124 = T_122 & 8'haa;
  assign T_125 = T_120 | T_124;
  assign T_126 = T_93[9:8];
  assign T_127 = T_126[0];
  assign T_128 = T_126[1];
  assign T_129 = {T_127,T_128};
  assign T_130 = {T_125,T_129};
  assign T_132 = {T_130,14'h3fff};
  assign T_135 = T_92[13:0];
  assign T_136 = T_135[7:0];
  assign T_141 = T_136[7:4];
  assign T_142 = {{4'd0}, T_141};
  assign T_143 = T_136[3:0];
  assign GEN_7 = {{4'd0}, T_143};
  assign T_144 = GEN_7 << 4;
  assign T_146 = T_144 & 8'hf0;
  assign T_147 = T_142 | T_146;
  assign T_151 = T_147[7:2];
  assign GEN_8 = {{2'd0}, T_151};
  assign T_152 = GEN_8 & 8'h33;
  assign T_153 = T_147[5:0];
  assign GEN_9 = {{2'd0}, T_153};
  assign T_154 = GEN_9 << 2;
  assign T_156 = T_154 & 8'hcc;
  assign T_157 = T_152 | T_156;
  assign T_161 = T_157[7:1];
  assign GEN_10 = {{1'd0}, T_161};
  assign T_162 = GEN_10 & 8'h55;
  assign T_163 = T_157[6:0];
  assign GEN_11 = {{1'd0}, T_163};
  assign T_164 = GEN_11 << 1;
  assign T_166 = T_164 & 8'haa;
  assign T_167 = T_162 | T_166;
  assign T_168 = T_135[13:8];
  assign T_169 = T_168[3:0];
  assign T_170 = T_169[1:0];
  assign T_171 = T_170[0];
  assign T_172 = T_170[1];
  assign T_173 = {T_171,T_172};
  assign T_174 = T_169[3:2];
  assign T_175 = T_174[0];
  assign T_176 = T_174[1];
  assign T_177 = {T_175,T_176};
  assign T_178 = {T_173,T_177};
  assign T_179 = T_168[5:4];
  assign T_180 = T_179[0];
  assign T_181 = T_179[1];
  assign T_182 = {T_180,T_181};
  assign T_183 = {T_178,T_182};
  assign T_184 = {T_167,T_183};
  assign CExtraMask = T_89 ? T_132 : {{10'd0}, T_184};
  assign T_185 = ~ sigC;
  assign negSigC = doSubMags ? T_185 : sigC;
  assign T_189 = doSubMags ? 50'h3ffffffffffff : 50'h0;
  assign T_190 = {doSubMags,negSigC};
  assign T_191 = {T_190,T_189};
  assign T_192 = $signed(T_191);
  assign T_193 = $signed(T_192) >>> CAlignDist;
  assign T_194 = sigC & CExtraMask;
  assign T_196 = T_194 != 24'h0;
  assign T_197 = T_196 ^ doSubMags;
  assign T_198 = $unsigned(T_193);
  assign T_199 = {T_198,T_197};
  assign alignedNegSigC = T_199[74:0];
  assign T_200 = alignedNegSigC[48:1];
  assign T_202 = fractA[22];
  assign T_204 = fractB[22];
  assign T_206 = fractC[22];
  assign T_207 = alignedNegSigC[0];
  assign T_208 = alignedNegSigC[74:49];
endmodule
module MulAddRecFN_postMul(
  input   clk,
  input   reset,
  input  [2:0] io_fromPreMul_highExpA,
  input   io_fromPreMul_isNaN_isQuietNaNA,
  input  [2:0] io_fromPreMul_highExpB,
  input   io_fromPreMul_isNaN_isQuietNaNB,
  input   io_fromPreMul_signProd,
  input   io_fromPreMul_isZeroProd,
  input   io_fromPreMul_opSignC,
  input  [2:0] io_fromPreMul_highExpC,
  input   io_fromPreMul_isNaN_isQuietNaNC,
  input   io_fromPreMul_isCDominant,
  input   io_fromPreMul_CAlignDist_0,
  input  [6:0] io_fromPreMul_CAlignDist,
  input   io_fromPreMul_bit0AlignedNegSigC,
  input  [25:0] io_fromPreMul_highAlignedNegSigC,
  input  [10:0] io_fromPreMul_sExpSum,
  input  [1:0] io_fromPreMul_roundingMode,
  input  [48:0] io_mulAddResult,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  isZeroA;
  wire [1:0] T_38;
  wire  isSpecialA;
  wire  T_40;
  wire  T_42;
  wire  isInfA;
  wire  isNaNA;
  wire  T_45;
  wire  isSigNaNA;
  wire  isZeroB;
  wire [1:0] T_47;
  wire  isSpecialB;
  wire  T_49;
  wire  T_51;
  wire  isInfB;
  wire  isNaNB;
  wire  T_54;
  wire  isSigNaNB;
  wire  isZeroC;
  wire [1:0] T_56;
  wire  isSpecialC;
  wire  T_58;
  wire  T_60;
  wire  isInfC;
  wire  isNaNC;
  wire  T_63;
  wire  isSigNaNC;
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  doSubMags;
  wire  T_70;
  wire [26:0] T_72;
  wire [25:0] T_73;
  wire [25:0] T_74;
  wire [47:0] T_75;
  wire [73:0] T_76;
  wire [74:0] sigSum;
  wire [49:0] T_78;
  wire [50:0] GEN_0;
  wire [50:0] T_81;
  wire [50:0] T_82;
  wire [49:0] T_84;
  wire [17:0] T_85;
  wire [31:0] T_86;
  wire  T_88;
  wire [1:0] T_89;
  wire [15:0] T_90;
  wire  T_92;
  wire  T_93;
  wire [7:0] T_94;
  wire [7:0] T_95;
  wire  T_97;
  wire [3:0] T_98;
  wire [3:0] T_99;
  wire  T_101;
  wire  T_102;
  wire  T_104;
  wire  T_106;
  wire [1:0] T_108;
  wire [1:0] T_109;
  wire  T_110;
  wire  T_112;
  wire  T_114;
  wire [1:0] T_116;
  wire [1:0] T_117;
  wire [1:0] T_118;
  wire [2:0] T_119;
  wire [3:0] T_120;
  wire [3:0] T_121;
  wire  T_123;
  wire  T_124;
  wire  T_126;
  wire  T_128;
  wire [1:0] T_130;
  wire [1:0] T_131;
  wire  T_132;
  wire  T_134;
  wire  T_136;
  wire [1:0] T_138;
  wire [1:0] T_139;
  wire [1:0] T_140;
  wire [2:0] T_141;
  wire [2:0] T_142;
  wire [3:0] T_143;
  wire [3:0] T_145;
  wire [4:0] T_146;
  wire [15:0] T_147;
  wire [15:0] T_148;
  wire  T_150;
  wire [7:0] T_151;
  wire [7:0] T_152;
  wire  T_154;
  wire [3:0] T_155;
  wire [3:0] T_156;
  wire  T_158;
  wire  T_159;
  wire  T_161;
  wire  T_163;
  wire [1:0] T_165;
  wire [1:0] T_166;
  wire  T_167;
  wire  T_169;
  wire  T_171;
  wire [1:0] T_173;
  wire [1:0] T_174;
  wire [1:0] T_175;
  wire [2:0] T_176;
  wire [3:0] T_177;
  wire [3:0] T_178;
  wire  T_180;
  wire  T_181;
  wire  T_183;
  wire  T_185;
  wire [1:0] T_187;
  wire [1:0] T_188;
  wire  T_189;
  wire  T_191;
  wire  T_193;
  wire [1:0] T_195;
  wire [1:0] T_196;
  wire [1:0] T_197;
  wire [2:0] T_198;
  wire [2:0] T_199;
  wire [3:0] T_200;
  wire [7:0] T_201;
  wire [7:0] T_202;
  wire  T_204;
  wire [3:0] T_205;
  wire [3:0] T_206;
  wire  T_208;
  wire  T_209;
  wire  T_211;
  wire  T_213;
  wire [1:0] T_215;
  wire [1:0] T_216;
  wire  T_217;
  wire  T_219;
  wire  T_221;
  wire [1:0] T_223;
  wire [1:0] T_224;
  wire [1:0] T_225;
  wire [2:0] T_226;
  wire [3:0] T_227;
  wire [3:0] T_228;
  wire  T_230;
  wire  T_231;
  wire  T_233;
  wire  T_235;
  wire [1:0] T_237;
  wire [1:0] T_238;
  wire  T_239;
  wire  T_241;
  wire  T_243;
  wire [1:0] T_245;
  wire [1:0] T_246;
  wire [1:0] T_247;
  wire [2:0] T_248;
  wire [2:0] T_249;
  wire [3:0] T_250;
  wire [3:0] T_251;
  wire [4:0] T_252;
  wire [4:0] T_253;
  wire [5:0] T_254;
  wire [6:0] GEN_2;
  wire [7:0] T_255;
  wire [6:0] estNormPos_dist;
  wire [15:0] T_256;
  wire  T_258;
  wire [17:0] T_259;
  wire  T_261;
  wire [1:0] firstReduceSigSum;
  wire [74:0] complSigSum;
  wire [15:0] T_262;
  wire  T_264;
  wire [17:0] T_265;
  wire  T_267;
  wire [1:0] firstReduceComplSigSum;
  wire  T_268;
  wire [7:0] T_270;
  wire [6:0] T_271;
  wire [4:0] T_272;
  wire [6:0] CDom_estNormDist;
  wire  T_274;
  wire  T_275;
  wire  T_277;
  wire  T_278;
  wire [40:0] T_279;
  wire  T_281;
  wire [41:0] T_282;
  wire [41:0] T_284;
  wire  T_288;
  wire [40:0] T_289;
  wire  T_290;
  wire [41:0] T_291;
  wire [41:0] T_293;
  wire [41:0] T_294;
  wire  T_298;
  wire [40:0] T_299;
  wire  T_301;
  wire [41:0] T_302;
  wire [41:0] T_304;
  wire [41:0] T_305;
  wire  T_307;
  wire [40:0] T_308;
  wire  T_309;
  wire [41:0] T_310;
  wire [41:0] T_312;
  wire [41:0] CDom_firstNormAbsSigSum;
  wire [32:0] T_313;
  wire  T_316;
  wire  T_318;
  wire [33:0] T_319;
  wire [41:0] T_320;
  wire  T_321;
  wire  T_322;
  wire [25:0] T_323;
  wire [15:0] T_327;
  wire [41:0] T_328;
  wire [41:0] T_329;
  wire [9:0] T_331;
  wire [31:0] T_335;
  wire [41:0] T_336;
  wire [41:0] T_337;
  wire [41:0] notCDom_pos_firstNormAbsSigSum;
  wire [31:0] T_338;
  wire [32:0] T_340;
  wire [41:0] T_341;
  wire [26:0] T_344;
  wire [42:0] GEN_3;
  wire [42:0] T_345;
  wire [42:0] T_346;
  wire [10:0] T_348;
  wire [42:0] GEN_4;
  wire [42:0] T_349;
  wire [42:0] T_350;
  wire [42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire  notCDom_signSigSum;
  wire  T_352;
  wire  T_353;
  wire  doNegSignSum;
  wire [6:0] estNormDist;
  wire [42:0] T_355;
  wire [41:0] T_356;
  wire [42:0] cFirstNormAbsSigSum;
  wire  T_358;
  wire  T_360;
  wire  T_361;
  wire  doIncrSig;
  wire [3:0] estNormDist_5;
  wire [3:0] normTo2ShiftDist;
  wire [16:0] T_363;
  wire [14:0] T_364;
  wire [7:0] T_365;
  wire [3:0] T_370;
  wire [7:0] T_371;
  wire [3:0] T_372;
  wire [7:0] GEN_5;
  wire [7:0] T_373;
  wire [7:0] T_375;
  wire [7:0] T_376;
  wire [5:0] T_380;
  wire [7:0] GEN_6;
  wire [7:0] T_381;
  wire [5:0] T_382;
  wire [7:0] GEN_7;
  wire [7:0] T_383;
  wire [7:0] T_385;
  wire [7:0] T_386;
  wire [6:0] T_390;
  wire [7:0] GEN_8;
  wire [7:0] T_391;
  wire [6:0] T_392;
  wire [7:0] GEN_9;
  wire [7:0] T_393;
  wire [7:0] T_395;
  wire [7:0] T_396;
  wire [6:0] T_397;
  wire [3:0] T_398;
  wire [1:0] T_399;
  wire  T_400;
  wire  T_401;
  wire [1:0] T_402;
  wire [1:0] T_403;
  wire  T_404;
  wire  T_405;
  wire [1:0] T_406;
  wire [3:0] T_407;
  wire [2:0] T_408;
  wire [1:0] T_409;
  wire  T_410;
  wire  T_411;
  wire [1:0] T_412;
  wire  T_413;
  wire [2:0] T_414;
  wire [6:0] T_415;
  wire [14:0] T_416;
  wire [15:0] absSigSumExtraMask;
  wire [41:0] T_418;
  wire [41:0] T_419;
  wire [15:0] T_420;
  wire [15:0] T_421;
  wire [15:0] T_422;
  wire  T_424;
  wire [15:0] T_426;
  wire  T_428;
  wire  T_429;
  wire [42:0] T_430;
  wire [27:0] sigX3;
  wire [1:0] T_431;
  wire  sigX3Shift1;
  wire [10:0] GEN_10;
  wire [11:0] T_433;
  wire [10:0] sExpX3;
  wire [2:0] T_434;
  wire  isZeroY;
  wire  T_436;
  wire  signY;
  wire [9:0] sExpX3_13;
  wire  T_437;
  wire [26:0] T_441;
  wire [9:0] T_442;
  wire  T_443;
  wire [8:0] T_444;
  wire  T_445;
  wire [7:0] T_446;
  wire  T_447;
  wire [6:0] T_448;
  wire  T_449;
  wire [5:0] T_450;
  wire [64:0] T_453;
  wire [20:0] T_454;
  wire [15:0] T_455;
  wire [7:0] T_460;
  wire [15:0] T_461;
  wire [7:0] T_462;
  wire [15:0] GEN_11;
  wire [15:0] T_463;
  wire [15:0] T_465;
  wire [15:0] T_466;
  wire [11:0] T_470;
  wire [15:0] GEN_12;
  wire [15:0] T_471;
  wire [11:0] T_472;
  wire [15:0] GEN_13;
  wire [15:0] T_473;
  wire [15:0] T_475;
  wire [15:0] T_476;
  wire [13:0] T_480;
  wire [15:0] GEN_14;
  wire [15:0] T_481;
  wire [13:0] T_482;
  wire [15:0] GEN_15;
  wire [15:0] T_483;
  wire [15:0] T_485;
  wire [15:0] T_486;
  wire [14:0] T_490;
  wire [15:0] GEN_16;
  wire [15:0] T_491;
  wire [14:0] T_492;
  wire [15:0] GEN_17;
  wire [15:0] T_493;
  wire [15:0] T_495;
  wire [15:0] T_496;
  wire [4:0] T_497;
  wire [3:0] T_498;
  wire [1:0] T_499;
  wire  T_500;
  wire  T_501;
  wire [1:0] T_502;
  wire [1:0] T_503;
  wire  T_504;
  wire  T_505;
  wire [1:0] T_506;
  wire [3:0] T_507;
  wire  T_508;
  wire [4:0] T_509;
  wire [20:0] T_510;
  wire [20:0] T_511;
  wire [20:0] T_512;
  wire [20:0] T_513;
  wire [24:0] T_515;
  wire [3:0] T_520;
  wire [1:0] T_521;
  wire  T_522;
  wire  T_523;
  wire [1:0] T_524;
  wire [1:0] T_525;
  wire  T_526;
  wire  T_527;
  wire [1:0] T_528;
  wire [3:0] T_529;
  wire [3:0] T_531;
  wire [24:0] T_532;
  wire [24:0] T_534;
  wire [24:0] T_536;
  wire  T_537;
  wire [24:0] GEN_18;
  wire [24:0] T_538;
  wire [26:0] T_540;
  wire [26:0] roundMask;
  wire [25:0] T_541;
  wire [25:0] T_542;
  wire [26:0] GEN_19;
  wire [26:0] roundPosMask;
  wire [27:0] GEN_20;
  wire [27:0] T_543;
  wire  roundPosBit;
  wire [27:0] GEN_21;
  wire [27:0] T_546;
  wire  anyRoundExtra;
  wire [27:0] T_548;
  wire [27:0] T_550;
  wire  allRoundExtra;
  wire  anyRound;
  wire  allRound;
  wire  roundDirectUp;
  wire  T_553;
  wire  T_554;
  wire  T_555;
  wire  T_556;
  wire  T_559;
  wire  T_560;
  wire  T_561;
  wire  T_562;
  wire  T_563;
  wire  T_564;
  wire  T_565;
  wire  T_566;
  wire  T_567;
  wire  roundUp;
  wire  T_571;
  wire  T_572;
  wire  T_573;
  wire  T_574;
  wire  T_576;
  wire  T_577;
  wire  roundEven;
  wire  T_579;
  wire  roundInexact;
  wire [27:0] GEN_23;
  wire [27:0] T_580;
  wire [25:0] T_581;
  wire [26:0] T_583;
  wire [25:0] T_584;
  wire  T_586;
  wire  T_588;
  wire  T_589;
  wire [26:0] T_590;
  wire [27:0] GEN_24;
  wire [27:0] T_591;
  wire [25:0] T_592;
  wire [25:0] T_594;
  wire [25:0] T_596;
  wire [25:0] T_597;
  wire [25:0] T_600;
  wire [25:0] T_602;
  wire [25:0] sigY3;
  wire  T_603;
  wire [11:0] T_605;
  wire [10:0] T_606;
  wire [10:0] T_608;
  wire  T_609;
  wire [10:0] T_611;
  wire [10:0] T_612;
  wire [1:0] T_613;
  wire  T_615;
  wire [11:0] T_617;
  wire [10:0] T_618;
  wire [10:0] T_620;
  wire [10:0] sExpY;
  wire [8:0] expY;
  wire [22:0] T_621;
  wire [22:0] T_622;
  wire [22:0] fractY;
  wire [2:0] T_623;
  wire  overflowY;
  wire  T_626;
  wire  T_627;
  wire  T_630;
  wire  T_631;
  wire  totalUnderflowY;
  wire [7:0] T_635;
  wire [9:0] GEN_25;
  wire  T_636;
  wire  T_637;
  wire  underflowY;
  wire  T_638;
  wire  T_640;
  wire  T_641;
  wire  roundMagUp;
  wire  overflowY_roundMagUp;
  wire  mulSpecial;
  wire  addSpecial;
  wire  notSpecial_addZeros;
  wire  T_643;
  wire  T_645;
  wire  commonCase;
  wire  T_646;
  wire  T_647;
  wire  T_648;
  wire  T_650;
  wire  T_652;
  wire  T_653;
  wire  T_654;
  wire  T_655;
  wire  T_656;
  wire  T_657;
  wire  notSigNaN_invalid;
  wire  T_658;
  wire  T_659;
  wire  invalid;
  wire  overflow;
  wire  underflow;
  wire  T_660;
  wire  inexact;
  wire  T_661;
  wire  notSpecial_isZeroOut;
  wire  T_662;
  wire  pegMinFiniteMagOut;
  wire  T_664;
  wire  pegMaxFiniteMagOut;
  wire  T_666;
  wire  T_667;
  wire  notNaN_isInfOut;
  wire  T_668;
  wire  T_669;
  wire  isNaNOut;
  wire  T_672;
  wire  T_674;
  wire  T_675;
  wire  T_676;
  wire  T_677;
  wire  T_679;
  wire  T_680;
  wire  T_681;
  wire  T_682;
  wire  T_685;
  wire  T_686;
  wire  T_687;
  wire  uncommonCaseSignOut;
  wire  T_689;
  wire  T_690;
  wire  T_691;
  wire  signOut;
  wire [8:0] T_694;
  wire [8:0] T_695;
  wire [8:0] T_696;
  wire [8:0] T_700;
  wire [8:0] T_701;
  wire [8:0] T_702;
  wire [8:0] T_705;
  wire [8:0] T_706;
  wire [8:0] T_707;
  wire [8:0] T_710;
  wire [8:0] T_711;
  wire [8:0] T_712;
  wire [8:0] T_715;
  wire [8:0] T_716;
  wire [8:0] T_719;
  wire [8:0] T_720;
  wire [8:0] T_723;
  wire [8:0] T_724;
  wire [8:0] T_727;
  wire [8:0] expOut;
  wire  T_728;
  wire  T_729;
  wire [22:0] T_733;
  wire [22:0] T_734;
  wire [22:0] T_738;
  wire [22:0] fractOut;
  wire [9:0] T_739;
  wire [32:0] T_740;
  wire [1:0] T_742;
  wire [1:0] T_743;
  wire [2:0] T_744;
  wire [4:0] T_745;
  assign io_out = T_740;
  assign io_exceptionFlags = T_745;
  assign isZeroA = io_fromPreMul_highExpA == 3'h0;
  assign T_38 = io_fromPreMul_highExpA[2:1];
  assign isSpecialA = T_38 == 2'h3;
  assign T_40 = io_fromPreMul_highExpA[0];
  assign T_42 = T_40 == 1'h0;
  assign isInfA = isSpecialA & T_42;
  assign isNaNA = isSpecialA & T_40;
  assign T_45 = io_fromPreMul_isNaN_isQuietNaNA == 1'h0;
  assign isSigNaNA = isNaNA & T_45;
  assign isZeroB = io_fromPreMul_highExpB == 3'h0;
  assign T_47 = io_fromPreMul_highExpB[2:1];
  assign isSpecialB = T_47 == 2'h3;
  assign T_49 = io_fromPreMul_highExpB[0];
  assign T_51 = T_49 == 1'h0;
  assign isInfB = isSpecialB & T_51;
  assign isNaNB = isSpecialB & T_49;
  assign T_54 = io_fromPreMul_isNaN_isQuietNaNB == 1'h0;
  assign isSigNaNB = isNaNB & T_54;
  assign isZeroC = io_fromPreMul_highExpC == 3'h0;
  assign T_56 = io_fromPreMul_highExpC[2:1];
  assign isSpecialC = T_56 == 2'h3;
  assign T_58 = io_fromPreMul_highExpC[0];
  assign T_60 = T_58 == 1'h0;
  assign isInfC = isSpecialC & T_60;
  assign isNaNC = isSpecialC & T_58;
  assign T_63 = io_fromPreMul_isNaN_isQuietNaNC == 1'h0;
  assign isSigNaNC = isNaNC & T_63;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T_70 = io_mulAddResult[48];
  assign T_72 = io_fromPreMul_highAlignedNegSigC + 26'h1;
  assign T_73 = T_72[25:0];
  assign T_74 = T_70 ? T_73 : io_fromPreMul_highAlignedNegSigC;
  assign T_75 = io_mulAddResult[47:0];
  assign T_76 = {T_74,T_75};
  assign sigSum = {T_76,io_fromPreMul_bit0AlignedNegSigC};
  assign T_78 = sigSum[50:1];
  assign GEN_0 = {{1'd0}, T_78};
  assign T_81 = GEN_0 << 1;
  assign T_82 = GEN_0 ^ T_81;
  assign T_84 = T_82[49:0];
  assign T_85 = T_84[49:32];
  assign T_86 = T_84[31:0];
  assign T_88 = T_85 != 18'h0;
  assign T_89 = T_85[17:16];
  assign T_90 = T_85[15:0];
  assign T_92 = T_89 != 2'h0;
  assign T_93 = T_89[1];
  assign T_94 = T_90[15:8];
  assign T_95 = T_90[7:0];
  assign T_97 = T_94 != 8'h0;
  assign T_98 = T_94[7:4];
  assign T_99 = T_94[3:0];
  assign T_101 = T_98 != 4'h0;
  assign T_102 = T_98[3];
  assign T_104 = T_98[2];
  assign T_106 = T_98[1];
  assign T_108 = T_104 ? 2'h2 : {{1'd0}, T_106};
  assign T_109 = T_102 ? 2'h3 : T_108;
  assign T_110 = T_99[3];
  assign T_112 = T_99[2];
  assign T_114 = T_99[1];
  assign T_116 = T_112 ? 2'h2 : {{1'd0}, T_114};
  assign T_117 = T_110 ? 2'h3 : T_116;
  assign T_118 = T_101 ? T_109 : T_117;
  assign T_119 = {T_101,T_118};
  assign T_120 = T_95[7:4];
  assign T_121 = T_95[3:0];
  assign T_123 = T_120 != 4'h0;
  assign T_124 = T_120[3];
  assign T_126 = T_120[2];
  assign T_128 = T_120[1];
  assign T_130 = T_126 ? 2'h2 : {{1'd0}, T_128};
  assign T_131 = T_124 ? 2'h3 : T_130;
  assign T_132 = T_121[3];
  assign T_134 = T_121[2];
  assign T_136 = T_121[1];
  assign T_138 = T_134 ? 2'h2 : {{1'd0}, T_136};
  assign T_139 = T_132 ? 2'h3 : T_138;
  assign T_140 = T_123 ? T_131 : T_139;
  assign T_141 = {T_123,T_140};
  assign T_142 = T_97 ? T_119 : T_141;
  assign T_143 = {T_97,T_142};
  assign T_145 = T_92 ? {{3'd0}, T_93} : T_143;
  assign T_146 = {T_92,T_145};
  assign T_147 = T_86[31:16];
  assign T_148 = T_86[15:0];
  assign T_150 = T_147 != 16'h0;
  assign T_151 = T_147[15:8];
  assign T_152 = T_147[7:0];
  assign T_154 = T_151 != 8'h0;
  assign T_155 = T_151[7:4];
  assign T_156 = T_151[3:0];
  assign T_158 = T_155 != 4'h0;
  assign T_159 = T_155[3];
  assign T_161 = T_155[2];
  assign T_163 = T_155[1];
  assign T_165 = T_161 ? 2'h2 : {{1'd0}, T_163};
  assign T_166 = T_159 ? 2'h3 : T_165;
  assign T_167 = T_156[3];
  assign T_169 = T_156[2];
  assign T_171 = T_156[1];
  assign T_173 = T_169 ? 2'h2 : {{1'd0}, T_171};
  assign T_174 = T_167 ? 2'h3 : T_173;
  assign T_175 = T_158 ? T_166 : T_174;
  assign T_176 = {T_158,T_175};
  assign T_177 = T_152[7:4];
  assign T_178 = T_152[3:0];
  assign T_180 = T_177 != 4'h0;
  assign T_181 = T_177[3];
  assign T_183 = T_177[2];
  assign T_185 = T_177[1];
  assign T_187 = T_183 ? 2'h2 : {{1'd0}, T_185};
  assign T_188 = T_181 ? 2'h3 : T_187;
  assign T_189 = T_178[3];
  assign T_191 = T_178[2];
  assign T_193 = T_178[1];
  assign T_195 = T_191 ? 2'h2 : {{1'd0}, T_193};
  assign T_196 = T_189 ? 2'h3 : T_195;
  assign T_197 = T_180 ? T_188 : T_196;
  assign T_198 = {T_180,T_197};
  assign T_199 = T_154 ? T_176 : T_198;
  assign T_200 = {T_154,T_199};
  assign T_201 = T_148[15:8];
  assign T_202 = T_148[7:0];
  assign T_204 = T_201 != 8'h0;
  assign T_205 = T_201[7:4];
  assign T_206 = T_201[3:0];
  assign T_208 = T_205 != 4'h0;
  assign T_209 = T_205[3];
  assign T_211 = T_205[2];
  assign T_213 = T_205[1];
  assign T_215 = T_211 ? 2'h2 : {{1'd0}, T_213};
  assign T_216 = T_209 ? 2'h3 : T_215;
  assign T_217 = T_206[3];
  assign T_219 = T_206[2];
  assign T_221 = T_206[1];
  assign T_223 = T_219 ? 2'h2 : {{1'd0}, T_221};
  assign T_224 = T_217 ? 2'h3 : T_223;
  assign T_225 = T_208 ? T_216 : T_224;
  assign T_226 = {T_208,T_225};
  assign T_227 = T_202[7:4];
  assign T_228 = T_202[3:0];
  assign T_230 = T_227 != 4'h0;
  assign T_231 = T_227[3];
  assign T_233 = T_227[2];
  assign T_235 = T_227[1];
  assign T_237 = T_233 ? 2'h2 : {{1'd0}, T_235};
  assign T_238 = T_231 ? 2'h3 : T_237;
  assign T_239 = T_228[3];
  assign T_241 = T_228[2];
  assign T_243 = T_228[1];
  assign T_245 = T_241 ? 2'h2 : {{1'd0}, T_243};
  assign T_246 = T_239 ? 2'h3 : T_245;
  assign T_247 = T_230 ? T_238 : T_246;
  assign T_248 = {T_230,T_247};
  assign T_249 = T_204 ? T_226 : T_248;
  assign T_250 = {T_204,T_249};
  assign T_251 = T_150 ? T_200 : T_250;
  assign T_252 = {T_150,T_251};
  assign T_253 = T_88 ? T_146 : T_252;
  assign T_254 = {T_88,T_253};
  assign GEN_2 = {{1'd0}, T_254};
  assign T_255 = 7'h49 - GEN_2;
  assign estNormPos_dist = T_255[6:0];
  assign T_256 = sigSum[33:18];
  assign T_258 = T_256 != 16'h0;
  assign T_259 = sigSum[17:0];
  assign T_261 = T_259 != 18'h0;
  assign firstReduceSigSum = {T_258,T_261};
  assign complSigSum = ~ sigSum;
  assign T_262 = complSigSum[33:18];
  assign T_264 = T_262 != 16'h0;
  assign T_265 = complSigSum[17:0];
  assign T_267 = T_265 != 18'h0;
  assign firstReduceComplSigSum = {T_264,T_267};
  assign T_268 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign T_270 = io_fromPreMul_CAlignDist - 7'h1;
  assign T_271 = T_270[6:0];
  assign T_272 = T_271[4:0];
  assign CDom_estNormDist = T_268 ? io_fromPreMul_CAlignDist : {{2'd0}, T_272};
  assign T_274 = doSubMags == 1'h0;
  assign T_275 = CDom_estNormDist[4];
  assign T_277 = T_275 == 1'h0;
  assign T_278 = T_274 & T_277;
  assign T_279 = sigSum[74:34];
  assign T_281 = firstReduceSigSum != 2'h0;
  assign T_282 = {T_279,T_281};
  assign T_284 = T_278 ? T_282 : 42'h0;
  assign T_288 = T_274 & T_275;
  assign T_289 = sigSum[58:18];
  assign T_290 = firstReduceSigSum[0];
  assign T_291 = {T_289,T_290};
  assign T_293 = T_288 ? T_291 : 42'h0;
  assign T_294 = T_284 | T_293;
  assign T_298 = doSubMags & T_277;
  assign T_299 = complSigSum[74:34];
  assign T_301 = firstReduceComplSigSum != 2'h0;
  assign T_302 = {T_299,T_301};
  assign T_304 = T_298 ? T_302 : 42'h0;
  assign T_305 = T_294 | T_304;
  assign T_307 = doSubMags & T_275;
  assign T_308 = complSigSum[58:18];
  assign T_309 = firstReduceComplSigSum[0];
  assign T_310 = {T_308,T_309};
  assign T_312 = T_307 ? T_310 : 42'h0;
  assign CDom_firstNormAbsSigSum = T_305 | T_312;
  assign T_313 = sigSum[50:18];
  assign T_316 = T_309 == 1'h0;
  assign T_318 = doSubMags ? T_316 : T_290;
  assign T_319 = {T_313,T_318};
  assign T_320 = sigSum[42:1];
  assign T_321 = estNormPos_dist[5];
  assign T_322 = estNormPos_dist[4];
  assign T_323 = sigSum[26:1];
  assign T_327 = doSubMags ? 16'hffff : 16'h0;
  assign T_328 = {T_323,T_327};
  assign T_329 = T_322 ? T_328 : T_320;
  assign T_331 = sigSum[10:1];
  assign T_335 = doSubMags ? 32'hffffffff : 32'h0;
  assign T_336 = {T_331,T_335};
  assign T_337 = T_322 ? {{8'd0}, T_319} : T_336;
  assign notCDom_pos_firstNormAbsSigSum = T_321 ? T_329 : T_337;
  assign T_338 = complSigSum[49:18];
  assign T_340 = {T_338,T_309};
  assign T_341 = complSigSum[42:1];
  assign T_344 = complSigSum[27:1];
  assign GEN_3 = {{16'd0}, T_344};
  assign T_345 = GEN_3 << 16;
  assign T_346 = T_322 ? T_345 : {{1'd0}, T_341};
  assign T_348 = complSigSum[11:1];
  assign GEN_4 = {{32'd0}, T_348};
  assign T_349 = GEN_4 << 32;
  assign T_350 = T_322 ? {{10'd0}, T_340} : T_349;
  assign notCDom_neg_cFirstNormAbsSigSum = T_321 ? T_346 : T_350;
  assign notCDom_signSigSum = sigSum[51];
  assign T_352 = isZeroC == 1'h0;
  assign T_353 = doSubMags & T_352;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T_353 : notCDom_signSigSum;
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : estNormPos_dist;
  assign T_355 = io_fromPreMul_isCDominant ? {{1'd0}, CDom_firstNormAbsSigSum} : notCDom_neg_cFirstNormAbsSigSum;
  assign T_356 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T_355 : {{1'd0}, T_356};
  assign T_358 = io_fromPreMul_isCDominant == 1'h0;
  assign T_360 = notCDom_signSigSum == 1'h0;
  assign T_361 = T_358 & T_360;
  assign doIncrSig = T_361 & doSubMags;
  assign estNormDist_5 = estNormDist[3:0];
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign T_363 = $signed(17'sh10000) >>> normTo2ShiftDist;
  assign T_364 = T_363[15:1];
  assign T_365 = T_364[7:0];
  assign T_370 = T_365[7:4];
  assign T_371 = {{4'd0}, T_370};
  assign T_372 = T_365[3:0];
  assign GEN_5 = {{4'd0}, T_372};
  assign T_373 = GEN_5 << 4;
  assign T_375 = T_373 & 8'hf0;
  assign T_376 = T_371 | T_375;
  assign T_380 = T_376[7:2];
  assign GEN_6 = {{2'd0}, T_380};
  assign T_381 = GEN_6 & 8'h33;
  assign T_382 = T_376[5:0];
  assign GEN_7 = {{2'd0}, T_382};
  assign T_383 = GEN_7 << 2;
  assign T_385 = T_383 & 8'hcc;
  assign T_386 = T_381 | T_385;
  assign T_390 = T_386[7:1];
  assign GEN_8 = {{1'd0}, T_390};
  assign T_391 = GEN_8 & 8'h55;
  assign T_392 = T_386[6:0];
  assign GEN_9 = {{1'd0}, T_392};
  assign T_393 = GEN_9 << 1;
  assign T_395 = T_393 & 8'haa;
  assign T_396 = T_391 | T_395;
  assign T_397 = T_364[14:8];
  assign T_398 = T_397[3:0];
  assign T_399 = T_398[1:0];
  assign T_400 = T_399[0];
  assign T_401 = T_399[1];
  assign T_402 = {T_400,T_401};
  assign T_403 = T_398[3:2];
  assign T_404 = T_403[0];
  assign T_405 = T_403[1];
  assign T_406 = {T_404,T_405};
  assign T_407 = {T_402,T_406};
  assign T_408 = T_397[6:4];
  assign T_409 = T_408[1:0];
  assign T_410 = T_409[0];
  assign T_411 = T_409[1];
  assign T_412 = {T_410,T_411};
  assign T_413 = T_408[2];
  assign T_414 = {T_412,T_413};
  assign T_415 = {T_407,T_414};
  assign T_416 = {T_396,T_415};
  assign absSigSumExtraMask = {T_416,1'h1};
  assign T_418 = cFirstNormAbsSigSum[42:1];
  assign T_419 = T_418 >> normTo2ShiftDist;
  assign T_420 = cFirstNormAbsSigSum[15:0];
  assign T_421 = ~ T_420;
  assign T_422 = T_421 & absSigSumExtraMask;
  assign T_424 = T_422 == 16'h0;
  assign T_426 = T_420 & absSigSumExtraMask;
  assign T_428 = T_426 != 16'h0;
  assign T_429 = doIncrSig ? T_424 : T_428;
  assign T_430 = {T_419,T_429};
  assign sigX3 = T_430[27:0];
  assign T_431 = sigX3[27:26];
  assign sigX3Shift1 = T_431 == 2'h0;
  assign GEN_10 = {{4'd0}, estNormDist};
  assign T_433 = io_fromPreMul_sExpSum - GEN_10;
  assign sExpX3 = T_433[10:0];
  assign T_434 = sigX3[27:25];
  assign isZeroY = T_434 == 3'h0;
  assign T_436 = io_fromPreMul_signProd ^ doNegSignSum;
  assign signY = isZeroY ? roundingMode_min : T_436;
  assign sExpX3_13 = sExpX3[9:0];
  assign T_437 = sExpX3[10];
  assign T_441 = T_437 ? 27'h7ffffff : 27'h0;
  assign T_442 = ~ sExpX3_13;
  assign T_443 = T_442[9];
  assign T_444 = T_442[8:0];
  assign T_445 = T_444[8];
  assign T_446 = T_444[7:0];
  assign T_447 = T_446[7];
  assign T_448 = T_446[6:0];
  assign T_449 = T_448[6];
  assign T_450 = T_448[5:0];
  assign T_453 = $signed(65'sh10000000000000000) >>> T_450;
  assign T_454 = T_453[63:43];
  assign T_455 = T_454[15:0];
  assign T_460 = T_455[15:8];
  assign T_461 = {{8'd0}, T_460};
  assign T_462 = T_455[7:0];
  assign GEN_11 = {{8'd0}, T_462};
  assign T_463 = GEN_11 << 8;
  assign T_465 = T_463 & 16'hff00;
  assign T_466 = T_461 | T_465;
  assign T_470 = T_466[15:4];
  assign GEN_12 = {{4'd0}, T_470};
  assign T_471 = GEN_12 & 16'hf0f;
  assign T_472 = T_466[11:0];
  assign GEN_13 = {{4'd0}, T_472};
  assign T_473 = GEN_13 << 4;
  assign T_475 = T_473 & 16'hf0f0;
  assign T_476 = T_471 | T_475;
  assign T_480 = T_476[15:2];
  assign GEN_14 = {{2'd0}, T_480};
  assign T_481 = GEN_14 & 16'h3333;
  assign T_482 = T_476[13:0];
  assign GEN_15 = {{2'd0}, T_482};
  assign T_483 = GEN_15 << 2;
  assign T_485 = T_483 & 16'hcccc;
  assign T_486 = T_481 | T_485;
  assign T_490 = T_486[15:1];
  assign GEN_16 = {{1'd0}, T_490};
  assign T_491 = GEN_16 & 16'h5555;
  assign T_492 = T_486[14:0];
  assign GEN_17 = {{1'd0}, T_492};
  assign T_493 = GEN_17 << 1;
  assign T_495 = T_493 & 16'haaaa;
  assign T_496 = T_491 | T_495;
  assign T_497 = T_454[20:16];
  assign T_498 = T_497[3:0];
  assign T_499 = T_498[1:0];
  assign T_500 = T_499[0];
  assign T_501 = T_499[1];
  assign T_502 = {T_500,T_501};
  assign T_503 = T_498[3:2];
  assign T_504 = T_503[0];
  assign T_505 = T_503[1];
  assign T_506 = {T_504,T_505};
  assign T_507 = {T_502,T_506};
  assign T_508 = T_497[4];
  assign T_509 = {T_507,T_508};
  assign T_510 = {T_496,T_509};
  assign T_511 = ~ T_510;
  assign T_512 = T_449 ? 21'h0 : T_511;
  assign T_513 = ~ T_512;
  assign T_515 = {T_513,4'hf};
  assign T_520 = T_453[3:0];
  assign T_521 = T_520[1:0];
  assign T_522 = T_521[0];
  assign T_523 = T_521[1];
  assign T_524 = {T_522,T_523};
  assign T_525 = T_520[3:2];
  assign T_526 = T_525[0];
  assign T_527 = T_525[1];
  assign T_528 = {T_526,T_527};
  assign T_529 = {T_524,T_528};
  assign T_531 = T_449 ? T_529 : 4'h0;
  assign T_532 = T_447 ? T_515 : {{21'd0}, T_531};
  assign T_534 = T_445 ? T_532 : 25'h0;
  assign T_536 = T_443 ? T_534 : 25'h0;
  assign T_537 = sigX3[26];
  assign GEN_18 = {{24'd0}, T_537};
  assign T_538 = T_536 | GEN_18;
  assign T_540 = {T_538,2'h3};
  assign roundMask = T_441 | T_540;
  assign T_541 = roundMask[26:1];
  assign T_542 = ~ T_541;
  assign GEN_19 = {{1'd0}, T_542};
  assign roundPosMask = GEN_19 & roundMask;
  assign GEN_20 = {{1'd0}, roundPosMask};
  assign T_543 = sigX3 & GEN_20;
  assign roundPosBit = T_543 != 28'h0;
  assign GEN_21 = {{2'd0}, T_541};
  assign T_546 = sigX3 & GEN_21;
  assign anyRoundExtra = T_546 != 28'h0;
  assign T_548 = ~ sigX3;
  assign T_550 = T_548 & GEN_21;
  assign allRoundExtra = T_550 == 28'h0;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign allRound = roundPosBit & allRoundExtra;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign T_553 = doIncrSig == 1'h0;
  assign T_554 = T_553 & roundingMode_nearest_even;
  assign T_555 = T_554 & roundPosBit;
  assign T_556 = T_555 & anyRoundExtra;
  assign T_559 = T_553 & roundDirectUp;
  assign T_560 = T_559 & anyRound;
  assign T_561 = T_556 | T_560;
  assign T_562 = doIncrSig & allRound;
  assign T_563 = T_561 | T_562;
  assign T_564 = doIncrSig & roundingMode_nearest_even;
  assign T_565 = T_564 & roundPosBit;
  assign T_566 = T_563 | T_565;
  assign T_567 = doIncrSig & roundDirectUp;
  assign roundUp = T_566 | T_567;
  assign T_571 = roundPosBit == 1'h0;
  assign T_572 = roundingMode_nearest_even & T_571;
  assign T_573 = T_572 & allRoundExtra;
  assign T_574 = roundingMode_nearest_even & roundPosBit;
  assign T_576 = anyRoundExtra == 1'h0;
  assign T_577 = T_574 & T_576;
  assign roundEven = doIncrSig ? T_573 : T_577;
  assign T_579 = allRound == 1'h0;
  assign roundInexact = doIncrSig ? T_579 : anyRound;
  assign GEN_23 = {{1'd0}, roundMask};
  assign T_580 = sigX3 | GEN_23;
  assign T_581 = T_580[27:2];
  assign T_583 = T_581 + 26'h1;
  assign T_584 = T_583[25:0];
  assign T_586 = roundUp == 1'h0;
  assign T_588 = roundEven == 1'h0;
  assign T_589 = T_586 & T_588;
  assign T_590 = ~ roundMask;
  assign GEN_24 = {{1'd0}, T_590};
  assign T_591 = sigX3 & GEN_24;
  assign T_592 = T_591[27:2];
  assign T_594 = T_589 ? T_592 : 26'h0;
  assign T_596 = roundUp ? T_584 : 26'h0;
  assign T_597 = T_594 | T_596;
  assign T_600 = T_584 & T_542;
  assign T_602 = roundEven ? T_600 : 26'h0;
  assign sigY3 = T_597 | T_602;
  assign T_603 = sigY3[25];
  assign T_605 = sExpX3 + 11'h1;
  assign T_606 = T_605[10:0];
  assign T_608 = T_603 ? T_606 : 11'h0;
  assign T_609 = sigY3[24];
  assign T_611 = T_609 ? sExpX3 : 11'h0;
  assign T_612 = T_608 | T_611;
  assign T_613 = sigY3[25:24];
  assign T_615 = T_613 == 2'h0;
  assign T_617 = sExpX3 - 11'h1;
  assign T_618 = T_617[10:0];
  assign T_620 = T_615 ? T_618 : 11'h0;
  assign sExpY = T_612 | T_620;
  assign expY = sExpY[8:0];
  assign T_621 = sigY3[22:0];
  assign T_622 = sigY3[23:1];
  assign fractY = sigX3Shift1 ? T_621 : T_622;
  assign T_623 = sExpY[9:7];
  assign overflowY = T_623 == 3'h3;
  assign T_626 = isZeroY == 1'h0;
  assign T_627 = sExpY[9];
  assign T_630 = expY < 9'h6b;
  assign T_631 = T_627 | T_630;
  assign totalUnderflowY = T_626 & T_631;
  assign T_635 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign GEN_25 = {{2'd0}, T_635};
  assign T_636 = sExpX3_13 <= GEN_25;
  assign T_637 = T_437 | T_636;
  assign underflowY = roundInexact & T_637;
  assign T_638 = roundingMode_min & signY;
  assign T_640 = signY == 1'h0;
  assign T_641 = roundingMode_max & T_640;
  assign roundMagUp = T_638 | T_641;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign mulSpecial = isSpecialA | isSpecialB;
  assign addSpecial = mulSpecial | isSpecialC;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign T_643 = addSpecial == 1'h0;
  assign T_645 = notSpecial_addZeros == 1'h0;
  assign commonCase = T_643 & T_645;
  assign T_646 = isInfA & isZeroB;
  assign T_647 = isZeroA & isInfB;
  assign T_648 = T_646 | T_647;
  assign T_650 = isNaNA == 1'h0;
  assign T_652 = isNaNB == 1'h0;
  assign T_653 = T_650 & T_652;
  assign T_654 = isInfA | isInfB;
  assign T_655 = T_653 & T_654;
  assign T_656 = T_655 & isInfC;
  assign T_657 = T_656 & doSubMags;
  assign notSigNaN_invalid = T_648 | T_657;
  assign T_658 = isSigNaNA | isSigNaNB;
  assign T_659 = T_658 | isSigNaNC;
  assign invalid = T_659 | notSigNaN_invalid;
  assign overflow = commonCase & overflowY;
  assign underflow = commonCase & underflowY;
  assign T_660 = commonCase & roundInexact;
  assign inexact = overflow | T_660;
  assign T_661 = notSpecial_addZeros | isZeroY;
  assign notSpecial_isZeroOut = T_661 | totalUnderflowY;
  assign T_662 = commonCase & totalUnderflowY;
  assign pegMinFiniteMagOut = T_662 & roundMagUp;
  assign T_664 = overflowY_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = overflow & T_664;
  assign T_666 = T_654 | isInfC;
  assign T_667 = overflow & overflowY_roundMagUp;
  assign notNaN_isInfOut = T_666 | T_667;
  assign T_668 = isNaNA | isNaNB;
  assign T_669 = T_668 | isNaNC;
  assign isNaNOut = T_669 | notSigNaN_invalid;
  assign T_672 = T_274 & io_fromPreMul_opSignC;
  assign T_674 = isSpecialC == 1'h0;
  assign T_675 = mulSpecial & T_674;
  assign T_676 = T_675 & io_fromPreMul_signProd;
  assign T_677 = T_672 | T_676;
  assign T_679 = mulSpecial == 1'h0;
  assign T_680 = T_679 & isSpecialC;
  assign T_681 = T_680 & io_fromPreMul_opSignC;
  assign T_682 = T_677 | T_681;
  assign T_685 = T_679 & notSpecial_addZeros;
  assign T_686 = T_685 & doSubMags;
  assign T_687 = T_686 & roundingMode_min;
  assign uncommonCaseSignOut = T_682 | T_687;
  assign T_689 = isNaNOut == 1'h0;
  assign T_690 = T_689 & uncommonCaseSignOut;
  assign T_691 = commonCase & signY;
  assign signOut = T_690 | T_691;
  assign T_694 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign T_695 = ~ T_694;
  assign T_696 = expY & T_695;
  assign T_700 = pegMinFiniteMagOut ? 9'h194 : 9'h0;
  assign T_701 = ~ T_700;
  assign T_702 = T_696 & T_701;
  assign T_705 = pegMaxFiniteMagOut ? 9'h80 : 9'h0;
  assign T_706 = ~ T_705;
  assign T_707 = T_702 & T_706;
  assign T_710 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T_711 = ~ T_710;
  assign T_712 = T_707 & T_711;
  assign T_715 = pegMinFiniteMagOut ? 9'h6b : 9'h0;
  assign T_716 = T_712 | T_715;
  assign T_719 = pegMaxFiniteMagOut ? 9'h17f : 9'h0;
  assign T_720 = T_716 | T_719;
  assign T_723 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign T_724 = T_720 | T_723;
  assign T_727 = isNaNOut ? 9'h1c0 : 9'h0;
  assign expOut = T_724 | T_727;
  assign T_728 = totalUnderflowY & roundMagUp;
  assign T_729 = T_728 | isNaNOut;
  assign T_733 = isNaNOut ? 23'h400000 : 23'h0;
  assign T_734 = T_729 ? T_733 : fractY;
  assign T_738 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0;
  assign fractOut = T_734 | T_738;
  assign T_739 = {signOut,expOut};
  assign T_740 = {T_739,fractOut};
  assign T_742 = {underflow,inexact};
  assign T_743 = {invalid,1'h0};
  assign T_744 = {T_743,overflow};
  assign T_745 = {T_744,T_742};
endmodule
module MulAddRecFN(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  mulAddRecFN_preMul_clk;
  wire  mulAddRecFN_preMul_reset;
  wire [1:0] mulAddRecFN_preMul_io_op;
  wire [32:0] mulAddRecFN_preMul_io_a;
  wire [32:0] mulAddRecFN_preMul_io_b;
  wire [32:0] mulAddRecFN_preMul_io_c;
  wire [1:0] mulAddRecFN_preMul_io_roundingMode;
  wire [23:0] mulAddRecFN_preMul_io_mulAddA;
  wire [23:0] mulAddRecFN_preMul_io_mulAddB;
  wire [47:0] mulAddRecFN_preMul_io_mulAddC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_preMul_io_toPostMul_signProd;
  wire  mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire  mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire  mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire [6:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire  mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire [25:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire [10:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire [1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire  mulAddRecFN_postMul_clk;
  wire  mulAddRecFN_postMul_reset;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpA;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpB;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_postMul_io_fromPreMul_signProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_isZeroProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_opSignC;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isCDominant;
  wire  mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0;
  wire [6:0] mulAddRecFN_postMul_io_fromPreMul_CAlignDist;
  wire  mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC;
  wire [25:0] mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC;
  wire [10:0] mulAddRecFN_postMul_io_fromPreMul_sExpSum;
  wire [1:0] mulAddRecFN_postMul_io_fromPreMul_roundingMode;
  wire [48:0] mulAddRecFN_postMul_io_mulAddResult;
  wire [32:0] mulAddRecFN_postMul_io_out;
  wire [4:0] mulAddRecFN_postMul_io_exceptionFlags;
  wire [47:0] T_7;
  wire [48:0] T_9;
  wire [48:0] GEN_0;
  wire [49:0] T_10;
  wire [48:0] T_11;
  MulAddRecFN_preMul mulAddRecFN_preMul (
    .clk(mulAddRecFN_preMul_clk),
    .reset(mulAddRecFN_preMul_reset),
    .io_op(mulAddRecFN_preMul_io_op),
    .io_a(mulAddRecFN_preMul_io_a),
    .io_b(mulAddRecFN_preMul_io_b),
    .io_c(mulAddRecFN_preMul_io_c),
    .io_roundingMode(mulAddRecFN_preMul_io_roundingMode),
    .io_mulAddA(mulAddRecFN_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFN_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFN_preMul_io_mulAddC),
    .io_toPostMul_highExpA(mulAddRecFN_preMul_io_toPostMul_highExpA),
    .io_toPostMul_isNaN_isQuietNaNA(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA),
    .io_toPostMul_highExpB(mulAddRecFN_preMul_io_toPostMul_highExpB),
    .io_toPostMul_isNaN_isQuietNaNB(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB),
    .io_toPostMul_signProd(mulAddRecFN_preMul_io_toPostMul_signProd),
    .io_toPostMul_isZeroProd(mulAddRecFN_preMul_io_toPostMul_isZeroProd),
    .io_toPostMul_opSignC(mulAddRecFN_preMul_io_toPostMul_opSignC),
    .io_toPostMul_highExpC(mulAddRecFN_preMul_io_toPostMul_highExpC),
    .io_toPostMul_isNaN_isQuietNaNC(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC),
    .io_toPostMul_isCDominant(mulAddRecFN_preMul_io_toPostMul_isCDominant),
    .io_toPostMul_CAlignDist_0(mulAddRecFN_preMul_io_toPostMul_CAlignDist_0),
    .io_toPostMul_CAlignDist(mulAddRecFN_preMul_io_toPostMul_CAlignDist),
    .io_toPostMul_bit0AlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC),
    .io_toPostMul_highAlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC),
    .io_toPostMul_sExpSum(mulAddRecFN_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_roundingMode(mulAddRecFN_preMul_io_toPostMul_roundingMode)
  );
  MulAddRecFN_postMul mulAddRecFN_postMul (
    .clk(mulAddRecFN_postMul_clk),
    .reset(mulAddRecFN_postMul_reset),
    .io_fromPreMul_highExpA(mulAddRecFN_postMul_io_fromPreMul_highExpA),
    .io_fromPreMul_isNaN_isQuietNaNA(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA),
    .io_fromPreMul_highExpB(mulAddRecFN_postMul_io_fromPreMul_highExpB),
    .io_fromPreMul_isNaN_isQuietNaNB(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB),
    .io_fromPreMul_signProd(mulAddRecFN_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isZeroProd(mulAddRecFN_postMul_io_fromPreMul_isZeroProd),
    .io_fromPreMul_opSignC(mulAddRecFN_postMul_io_fromPreMul_opSignC),
    .io_fromPreMul_highExpC(mulAddRecFN_postMul_io_fromPreMul_highExpC),
    .io_fromPreMul_isNaN_isQuietNaNC(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC),
    .io_fromPreMul_isCDominant(mulAddRecFN_postMul_io_fromPreMul_isCDominant),
    .io_fromPreMul_CAlignDist_0(mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0),
    .io_fromPreMul_CAlignDist(mulAddRecFN_postMul_io_fromPreMul_CAlignDist),
    .io_fromPreMul_bit0AlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC),
    .io_fromPreMul_highAlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC),
    .io_fromPreMul_sExpSum(mulAddRecFN_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_roundingMode(mulAddRecFN_postMul_io_fromPreMul_roundingMode),
    .io_mulAddResult(mulAddRecFN_postMul_io_mulAddResult),
    .io_out(mulAddRecFN_postMul_io_out),
    .io_exceptionFlags(mulAddRecFN_postMul_io_exceptionFlags)
  );
  assign io_out = mulAddRecFN_postMul_io_out;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign mulAddRecFN_preMul_clk = clk;
  assign mulAddRecFN_preMul_reset = reset;
  assign mulAddRecFN_preMul_io_op = io_op;
  assign mulAddRecFN_preMul_io_a = io_a;
  assign mulAddRecFN_preMul_io_b = io_b;
  assign mulAddRecFN_preMul_io_c = io_c;
  assign mulAddRecFN_preMul_io_roundingMode = io_roundingMode;
  assign mulAddRecFN_postMul_clk = clk;
  assign mulAddRecFN_postMul_reset = reset;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpA = mulAddRecFN_preMul_io_toPostMul_highExpA;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpB = mulAddRecFN_preMul_io_toPostMul_highExpB;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  assign mulAddRecFN_postMul_io_fromPreMul_signProd = mulAddRecFN_preMul_io_toPostMul_signProd;
  assign mulAddRecFN_postMul_io_fromPreMul_isZeroProd = mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  assign mulAddRecFN_postMul_io_fromPreMul_opSignC = mulAddRecFN_preMul_io_toPostMul_opSignC;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpC = mulAddRecFN_preMul_io_toPostMul_highExpC;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  assign mulAddRecFN_postMul_io_fromPreMul_isCDominant = mulAddRecFN_preMul_io_toPostMul_isCDominant;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0 = mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist = mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  assign mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_sExpSum = mulAddRecFN_preMul_io_toPostMul_sExpSum;
  assign mulAddRecFN_postMul_io_fromPreMul_roundingMode = mulAddRecFN_preMul_io_toPostMul_roundingMode;
  assign mulAddRecFN_postMul_io_mulAddResult = T_11;
  assign T_7 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign T_9 = {1'h0,mulAddRecFN_preMul_io_mulAddC};
  assign GEN_0 = {{1'd0}, T_7};
  assign T_10 = GEN_0 + T_9;
  assign T_11 = T_10[48:0];
endmodule
module FPUFMAPipe(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [32:0] GEN_26;
  wire [32:0] zero;
  reg  valid;
  reg [31:0] GEN_27;
  reg [4:0] in_cmd;
  reg [31:0] GEN_28;
  reg  in_ldst;
  reg [31:0] GEN_29;
  reg  in_wen;
  reg [31:0] GEN_30;
  reg  in_ren1;
  reg [31:0] GEN_31;
  reg  in_ren2;
  reg [31:0] GEN_32;
  reg  in_ren3;
  reg [31:0] GEN_33;
  reg  in_swap12;
  reg [31:0] GEN_34;
  reg  in_swap23;
  reg [31:0] GEN_35;
  reg  in_single;
  reg [31:0] GEN_36;
  reg  in_fromint;
  reg [31:0] GEN_37;
  reg  in_toint;
  reg [31:0] GEN_38;
  reg  in_fastpipe;
  reg [31:0] GEN_39;
  reg  in_fma;
  reg [31:0] GEN_40;
  reg  in_div;
  reg [31:0] GEN_41;
  reg  in_sqrt;
  reg [31:0] GEN_42;
  reg  in_round;
  reg [31:0] GEN_43;
  reg  in_wflags;
  reg [31:0] GEN_44;
  reg [2:0] in_rm;
  reg [31:0] GEN_45;
  reg [1:0] in_typ;
  reg [31:0] GEN_46;
  reg [64:0] in_in1;
  reg [95:0] GEN_47;
  reg [64:0] in_in2;
  reg [95:0] GEN_48;
  reg [64:0] in_in3;
  reg [95:0] GEN_49;
  wire  T_179;
  wire  T_180;
  wire  T_181;
  wire  T_182;
  wire [1:0] T_183;
  wire [64:0] GEN_0;
  wire  T_186;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  fma_clk;
  wire  fma_reset;
  wire [1:0] fma_io_op;
  wire [32:0] fma_io_a;
  wire [32:0] fma_io_b;
  wire [32:0] fma_io_c;
  wire [1:0] fma_io_roundingMode;
  wire [32:0] fma_io_out;
  wire [4:0] fma_io_exceptionFlags;
  wire [64:0] res_data;
  wire [4:0] res_exc;
  wire [64:0] T_193;
  reg  T_196;
  reg [31:0] GEN_50;
  reg [64:0] T_197_data;
  reg [95:0] GEN_51;
  reg [4:0] T_197_exc;
  reg [31:0] GEN_52;
  wire [64:0] GEN_24;
  wire [4:0] GEN_25;
  wire  T_208_valid;
  wire [64:0] T_208_bits_data;
  wire [4:0] T_208_bits_exc;
  MulAddRecFN fma (
    .clk(fma_clk),
    .reset(fma_reset),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags)
  );
  assign io_out_valid = T_208_valid;
  assign io_out_bits_data = T_208_bits_data;
  assign io_out_bits_exc = T_208_bits_exc;
  assign T_131 = io_in_bits_in1[32];
  assign T_132 = io_in_bits_in2[32];
  assign T_133 = T_131 ^ T_132;
  assign GEN_26 = {{32'd0}, T_133};
  assign zero = GEN_26 << 32;
  assign T_179 = io_in_bits_cmd[1];
  assign T_180 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T_181 = T_179 & T_180;
  assign T_182 = io_in_bits_cmd[0];
  assign T_183 = {T_181,T_182};
  assign GEN_0 = io_in_bits_swap23 ? 65'h80000000 : io_in_bits_in2;
  assign T_186 = T_180 == 1'h0;
  assign GEN_1 = T_186 ? {{32'd0}, zero} : io_in_bits_in3;
  assign GEN_2 = io_in_valid ? {{3'd0}, T_183} : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_0 : in_in2;
  assign GEN_23 = io_in_valid ? GEN_1 : in_in3;
  assign fma_clk = clk;
  assign fma_reset = reset;
  assign fma_io_op = in_cmd[1:0];
  assign fma_io_a = in_in1[32:0];
  assign fma_io_b = in_in2[32:0];
  assign fma_io_c = in_in3[32:0];
  assign fma_io_roundingMode = in_rm[1:0];
  assign res_data = T_193;
  assign res_exc = fma_io_exceptionFlags;
  assign T_193 = {32'hffffffff,fma_io_out};
  assign GEN_24 = valid ? res_data : T_197_data;
  assign GEN_25 = valid ? res_exc : T_197_exc;
  assign T_208_valid = T_196;
  assign T_208_bits_data = T_197_data;
  assign T_208_bits_exc = T_197_exc;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  valid = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  in_cmd = GEN_28[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  in_ldst = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  in_wen = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  in_ren1 = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  in_ren2 = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  in_ren3 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  in_swap12 = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  in_swap23 = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  in_single = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  in_fromint = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  in_toint = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  in_fastpipe = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  in_fma = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  in_div = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  in_sqrt = GEN_42[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  in_round = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  in_wflags = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  in_rm = GEN_45[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  in_typ = GEN_46[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {3{$random}};
  in_in1 = GEN_47[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {3{$random}};
  in_in2 = GEN_48[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {3{$random}};
  in_in3 = GEN_49[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  T_196 = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {3{$random}};
  T_197_data = GEN_51[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  T_197_exc = GEN_52[4:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_cmd <= {{3'd0}, T_183};
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ldst <= io_in_bits_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wen <= io_in_bits_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren1 <= io_in_bits_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren2 <= io_in_bits_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren3 <= io_in_bits_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap12 <= io_in_bits_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap23 <= io_in_bits_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_single <= io_in_bits_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fromint <= io_in_bits_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_toint <= io_in_bits_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fastpipe <= io_in_bits_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fma <= io_in_bits_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_div <= io_in_bits_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_sqrt <= io_in_bits_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_round <= io_in_bits_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wflags <= io_in_bits_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_rm <= io_in_bits_rm;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_typ <= io_in_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_in1 <= io_in_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(io_in_bits_swap23) begin
          in_in2 <= 65'h80000000;
        end else begin
          in_in2 <= io_in_bits_in2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(T_186) begin
          in_in3 <= {{32'd0}, zero};
        end else begin
          in_in3 <= io_in_bits_in3;
        end
      end
    end
    if(reset) begin
      T_196 <= 1'h0;
    end else begin
      T_196 <= valid;
    end
    if(1'h0) begin
    end else begin
      if(valid) begin
        T_197_data <= res_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(valid) begin
        T_197_exc <= res_exc;
      end
    end
  end
endmodule
module CompareRecFN(
  input   clk,
  input   reset,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input   io_signaling,
  output  io_lt,
  output  io_eq,
  output  io_gt,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_7;
  wire [2:0] T_8;
  wire  T_10;
  wire [1:0] T_11;
  wire  T_13;
  wire  rawA_sign;
  wire  rawA_isNaN;
  wire  rawA_isInf;
  wire  rawA_isZero;
  wire [12:0] rawA_sExp;
  wire [55:0] rawA_sig;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_32;
  wire  T_33;
  wire [12:0] T_34;
  wire  T_37;
  wire [51:0] T_38;
  wire [53:0] T_40;
  wire [1:0] T_41;
  wire [55:0] T_42;
  wire [11:0] T_43;
  wire [2:0] T_44;
  wire  T_46;
  wire [1:0] T_47;
  wire  T_49;
  wire  rawB_sign;
  wire  rawB_isNaN;
  wire  rawB_isInf;
  wire  rawB_isZero;
  wire [12:0] rawB_sExp;
  wire [55:0] rawB_sig;
  wire  T_63;
  wire  T_64;
  wire  T_65;
  wire  T_68;
  wire  T_69;
  wire [12:0] T_70;
  wire  T_73;
  wire [51:0] T_74;
  wire [53:0] T_76;
  wire [1:0] T_77;
  wire [55:0] T_78;
  wire  T_80;
  wire  T_82;
  wire  ordered;
  wire  bothInfs;
  wire  bothZeros;
  wire  eqExps;
  wire  T_83;
  wire  T_84;
  wire  T_85;
  wire  common_ltMags;
  wire  T_86;
  wire  common_eqMags;
  wire  T_88;
  wire  T_90;
  wire  T_91;
  wire  T_93;
  wire  T_95;
  wire  T_96;
  wire  T_98;
  wire  T_99;
  wire  T_102;
  wire  T_103;
  wire  T_104;
  wire  T_105;
  wire  ordered_lt;
  wire  T_106;
  wire  T_107;
  wire  T_108;
  wire  ordered_eq;
  wire  T_109;
  wire  T_111;
  wire  T_112;
  wire  T_113;
  wire  T_115;
  wire  T_116;
  wire  T_117;
  wire  T_119;
  wire  T_120;
  wire  invalid;
  wire  T_121;
  wire  T_122;
  wire  T_124;
  wire  T_125;
  wire  T_127;
  wire  T_128;
  wire [4:0] T_130;
  assign io_lt = T_121;
  assign io_eq = T_122;
  assign io_gt = T_128;
  assign io_exceptionFlags = T_130;
  assign T_7 = io_a[63:52];
  assign T_8 = T_7[11:9];
  assign T_10 = T_8 == 3'h0;
  assign T_11 = T_7[11:10];
  assign T_13 = T_11 == 2'h3;
  assign rawA_sign = T_27;
  assign rawA_isNaN = T_29;
  assign rawA_isInf = T_33;
  assign rawA_isZero = T_10;
  assign rawA_sExp = T_34;
  assign rawA_sig = T_42;
  assign T_27 = io_a[64];
  assign T_28 = T_7[9];
  assign T_29 = T_13 & T_28;
  assign T_32 = T_28 == 1'h0;
  assign T_33 = T_13 & T_32;
  assign T_34 = {1'b0,$signed(T_7)};
  assign T_37 = T_10 == 1'h0;
  assign T_38 = io_a[51:0];
  assign T_40 = {T_38,2'h0};
  assign T_41 = {1'h0,T_37};
  assign T_42 = {T_41,T_40};
  assign T_43 = io_b[63:52];
  assign T_44 = T_43[11:9];
  assign T_46 = T_44 == 3'h0;
  assign T_47 = T_43[11:10];
  assign T_49 = T_47 == 2'h3;
  assign rawB_sign = T_63;
  assign rawB_isNaN = T_65;
  assign rawB_isInf = T_69;
  assign rawB_isZero = T_46;
  assign rawB_sExp = T_70;
  assign rawB_sig = T_78;
  assign T_63 = io_b[64];
  assign T_64 = T_43[9];
  assign T_65 = T_49 & T_64;
  assign T_68 = T_64 == 1'h0;
  assign T_69 = T_49 & T_68;
  assign T_70 = {1'b0,$signed(T_43)};
  assign T_73 = T_46 == 1'h0;
  assign T_74 = io_b[51:0];
  assign T_76 = {T_74,2'h0};
  assign T_77 = {1'h0,T_73};
  assign T_78 = {T_77,T_76};
  assign T_80 = rawA_isNaN == 1'h0;
  assign T_82 = rawB_isNaN == 1'h0;
  assign ordered = T_80 & T_82;
  assign bothInfs = rawA_isInf & rawB_isInf;
  assign bothZeros = rawA_isZero & rawB_isZero;
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp);
  assign T_83 = $signed(rawA_sExp) < $signed(rawB_sExp);
  assign T_84 = rawA_sig < rawB_sig;
  assign T_85 = eqExps & T_84;
  assign common_ltMags = T_83 | T_85;
  assign T_86 = rawA_sig == rawB_sig;
  assign common_eqMags = eqExps & T_86;
  assign T_88 = bothZeros == 1'h0;
  assign T_90 = rawB_sign == 1'h0;
  assign T_91 = rawA_sign & T_90;
  assign T_93 = bothInfs == 1'h0;
  assign T_95 = common_ltMags == 1'h0;
  assign T_96 = rawA_sign & T_95;
  assign T_98 = common_eqMags == 1'h0;
  assign T_99 = T_96 & T_98;
  assign T_102 = T_90 & common_ltMags;
  assign T_103 = T_99 | T_102;
  assign T_104 = T_93 & T_103;
  assign T_105 = T_91 | T_104;
  assign ordered_lt = T_88 & T_105;
  assign T_106 = rawA_sign == rawB_sign;
  assign T_107 = bothInfs | common_eqMags;
  assign T_108 = T_106 & T_107;
  assign ordered_eq = bothZeros | T_108;
  assign T_109 = rawA_sig[53];
  assign T_111 = T_109 == 1'h0;
  assign T_112 = rawA_isNaN & T_111;
  assign T_113 = rawB_sig[53];
  assign T_115 = T_113 == 1'h0;
  assign T_116 = rawB_isNaN & T_115;
  assign T_117 = T_112 | T_116;
  assign T_119 = ordered == 1'h0;
  assign T_120 = io_signaling & T_119;
  assign invalid = T_117 | T_120;
  assign T_121 = ordered & ordered_lt;
  assign T_122 = ordered & ordered_eq;
  assign T_124 = ordered_lt == 1'h0;
  assign T_125 = ordered & T_124;
  assign T_127 = ordered_eq == 1'h0;
  assign T_128 = T_125 & T_127;
  assign T_130 = {invalid,4'h0};
endmodule
module RecFNToIN(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  input   io_signedOut,
  output [31:0] io_out,
  output [2:0] io_intExceptionFlags
);
  wire  sign;
  wire [11:0] exp;
  wire [51:0] fract;
  wire [2:0] T_5;
  wire  isZero;
  wire [1:0] T_7;
  wire  isSpecial;
  wire  T_9;
  wire  isNaN;
  wire  notSpecial_magGeOne;
  wire [52:0] T_10;
  wire [4:0] T_11;
  wire [4:0] T_13;
  wire [83:0] GEN_0;
  wire [83:0] shiftedSig;
  wire [31:0] unroundedInt;
  wire [1:0] T_14;
  wire [50:0] T_15;
  wire  T_17;
  wire [2:0] roundBits;
  wire [1:0] T_18;
  wire  T_20;
  wire  T_22;
  wire  roundInexact;
  wire [1:0] T_23;
  wire [1:0] T_24;
  wire  T_26;
  wire [1:0] T_28;
  wire  T_30;
  wire  T_31;
  wire [10:0] T_32;
  wire [10:0] T_33;
  wire  T_35;
  wire  T_40;
  wire  roundIncr_nearestEven;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire  T_45;
  wire  T_46;
  wire  T_47;
  wire  T_49;
  wire  T_50;
  wire  T_51;
  wire  roundIncr;
  wire [31:0] T_52;
  wire [31:0] complUnroundedInt;
  wire  T_53;
  wire [32:0] T_55;
  wire [31:0] T_56;
  wire [31:0] roundedInt;
  wire [29:0] T_57;
  wire [29:0] T_58;
  wire  T_60;
  wire  roundCarryBut2;
  wire  T_62;
  wire  T_64;
  wire [30:0] T_67;
  wire  T_69;
  wire  T_70;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire  T_77;
  wire  T_78;
  wire  T_79;
  wire  T_80;
  wire  overflow_signed;
  wire  T_84;
  wire  T_87;
  wire  T_88;
  wire  T_89;
  wire  T_90;
  wire  T_91;
  wire  overflow_unsigned;
  wire  overflow;
  wire  T_93;
  wire  excSign;
  wire  T_94;
  wire [31:0] T_98;
  wire  T_100;
  wire  T_101;
  wire [30:0] T_104;
  wire [31:0] GEN_1;
  wire [31:0] T_105;
  wire  T_107;
  wire  T_110;
  wire [31:0] T_113;
  wire [31:0] excValue;
  wire  T_115;
  wire  T_116;
  wire  T_118;
  wire  inexact;
  wire  T_119;
  wire [31:0] T_120;
  wire [1:0] T_121;
  wire [2:0] T_122;
  assign io_out = T_120;
  assign io_intExceptionFlags = T_122;
  assign sign = io_in[64];
  assign exp = io_in[63:52];
  assign fract = io_in[51:0];
  assign T_5 = exp[11:9];
  assign isZero = T_5 == 3'h0;
  assign T_7 = exp[11:10];
  assign isSpecial = T_7 == 2'h3;
  assign T_9 = exp[9];
  assign isNaN = isSpecial & T_9;
  assign notSpecial_magGeOne = exp[11];
  assign T_10 = {notSpecial_magGeOne,fract};
  assign T_11 = exp[4:0];
  assign T_13 = notSpecial_magGeOne ? T_11 : 5'h0;
  assign GEN_0 = {{31'd0}, T_10};
  assign shiftedSig = GEN_0 << T_13;
  assign unroundedInt = shiftedSig[83:52];
  assign T_14 = shiftedSig[52:51];
  assign T_15 = shiftedSig[50:0];
  assign T_17 = T_15 != 51'h0;
  assign roundBits = {T_14,T_17};
  assign T_18 = roundBits[1:0];
  assign T_20 = T_18 != 2'h0;
  assign T_22 = isZero == 1'h0;
  assign roundInexact = notSpecial_magGeOne ? T_20 : T_22;
  assign T_23 = roundBits[2:1];
  assign T_24 = ~ T_23;
  assign T_26 = T_24 == 2'h0;
  assign T_28 = ~ T_18;
  assign T_30 = T_28 == 2'h0;
  assign T_31 = T_26 | T_30;
  assign T_32 = exp[10:0];
  assign T_33 = ~ T_32;
  assign T_35 = T_33 == 11'h0;
  assign T_40 = T_35 ? T_20 : 1'h0;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T_31 : T_40;
  assign T_41 = io_roundingMode == 2'h0;
  assign T_42 = T_41 & roundIncr_nearestEven;
  assign T_43 = io_roundingMode == 2'h2;
  assign T_44 = sign & roundInexact;
  assign T_45 = T_43 & T_44;
  assign T_46 = T_42 | T_45;
  assign T_47 = io_roundingMode == 2'h3;
  assign T_49 = sign == 1'h0;
  assign T_50 = T_49 & roundInexact;
  assign T_51 = T_47 & T_50;
  assign roundIncr = T_46 | T_51;
  assign T_52 = ~ unroundedInt;
  assign complUnroundedInt = sign ? T_52 : unroundedInt;
  assign T_53 = roundIncr ^ sign;
  assign T_55 = complUnroundedInt + 32'h1;
  assign T_56 = T_55[31:0];
  assign roundedInt = T_53 ? T_56 : complUnroundedInt;
  assign T_57 = unroundedInt[29:0];
  assign T_58 = ~ T_57;
  assign T_60 = T_58 == 30'h0;
  assign roundCarryBut2 = T_60 & roundIncr;
  assign T_62 = T_32 >= 11'h20;
  assign T_64 = T_32 == 11'h1f;
  assign T_67 = unroundedInt[30:0];
  assign T_69 = T_67 != 31'h0;
  assign T_70 = T_49 | T_69;
  assign T_71 = T_70 | roundIncr;
  assign T_72 = T_64 & T_71;
  assign T_73 = T_62 | T_72;
  assign T_77 = T_32 == 11'h1e;
  assign T_78 = T_49 & T_77;
  assign T_79 = T_78 & roundCarryBut2;
  assign T_80 = T_73 | T_79;
  assign overflow_signed = notSpecial_magGeOne ? T_80 : 1'h0;
  assign T_84 = sign | T_62;
  assign T_87 = unroundedInt[30];
  assign T_88 = T_64 & T_87;
  assign T_89 = T_88 & roundCarryBut2;
  assign T_90 = T_84 | T_89;
  assign T_91 = sign & roundIncr;
  assign overflow_unsigned = notSpecial_magGeOne ? T_90 : T_91;
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign T_93 = isNaN == 1'h0;
  assign excSign = sign & T_93;
  assign T_94 = io_signedOut & excSign;
  assign T_98 = T_94 ? 32'h80000000 : 32'h0;
  assign T_100 = excSign == 1'h0;
  assign T_101 = io_signedOut & T_100;
  assign T_104 = T_101 ? 31'h7fffffff : 31'h0;
  assign GEN_1 = {{1'd0}, T_104};
  assign T_105 = T_98 | GEN_1;
  assign T_107 = io_signedOut == 1'h0;
  assign T_110 = T_107 & T_100;
  assign T_113 = T_110 ? 32'hffffffff : 32'h0;
  assign excValue = T_105 | T_113;
  assign T_115 = isSpecial == 1'h0;
  assign T_116 = roundInexact & T_115;
  assign T_118 = overflow == 1'h0;
  assign inexact = T_116 & T_118;
  assign T_119 = isSpecial | overflow;
  assign T_120 = T_119 ? excValue : roundedInt;
  assign T_121 = {isSpecial,overflow};
  assign T_122 = {T_121,inexact};
endmodule
module RecFNToIN_1(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  input   io_signedOut,
  output [63:0] io_out,
  output [2:0] io_intExceptionFlags
);
  wire  sign;
  wire [11:0] exp;
  wire [51:0] fract;
  wire [2:0] T_5;
  wire  isZero;
  wire [1:0] T_7;
  wire  isSpecial;
  wire  T_9;
  wire  isNaN;
  wire  notSpecial_magGeOne;
  wire [52:0] T_10;
  wire [5:0] T_11;
  wire [5:0] T_13;
  wire [115:0] GEN_0;
  wire [115:0] shiftedSig;
  wire [63:0] unroundedInt;
  wire [1:0] T_14;
  wire [50:0] T_15;
  wire  T_17;
  wire [2:0] roundBits;
  wire [1:0] T_18;
  wire  T_20;
  wire  T_22;
  wire  roundInexact;
  wire [1:0] T_23;
  wire [1:0] T_24;
  wire  T_26;
  wire [1:0] T_28;
  wire  T_30;
  wire  T_31;
  wire [10:0] T_32;
  wire [10:0] T_33;
  wire  T_35;
  wire  T_40;
  wire  roundIncr_nearestEven;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire  T_45;
  wire  T_46;
  wire  T_47;
  wire  T_49;
  wire  T_50;
  wire  T_51;
  wire  roundIncr;
  wire [63:0] T_52;
  wire [63:0] complUnroundedInt;
  wire  T_53;
  wire [64:0] T_55;
  wire [63:0] T_56;
  wire [63:0] roundedInt;
  wire [61:0] T_57;
  wire [61:0] T_58;
  wire  T_60;
  wire  roundCarryBut2;
  wire  T_62;
  wire  T_64;
  wire [62:0] T_67;
  wire  T_69;
  wire  T_70;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire  T_77;
  wire  T_78;
  wire  T_79;
  wire  T_80;
  wire  overflow_signed;
  wire  T_84;
  wire  T_87;
  wire  T_88;
  wire  T_89;
  wire  T_90;
  wire  T_91;
  wire  overflow_unsigned;
  wire  overflow;
  wire  T_93;
  wire  excSign;
  wire  T_94;
  wire [63:0] T_98;
  wire  T_100;
  wire  T_101;
  wire [62:0] T_104;
  wire [63:0] GEN_1;
  wire [63:0] T_105;
  wire  T_107;
  wire  T_110;
  wire [63:0] T_113;
  wire [63:0] excValue;
  wire  T_115;
  wire  T_116;
  wire  T_118;
  wire  inexact;
  wire  T_119;
  wire [63:0] T_120;
  wire [1:0] T_121;
  wire [2:0] T_122;
  assign io_out = T_120;
  assign io_intExceptionFlags = T_122;
  assign sign = io_in[64];
  assign exp = io_in[63:52];
  assign fract = io_in[51:0];
  assign T_5 = exp[11:9];
  assign isZero = T_5 == 3'h0;
  assign T_7 = exp[11:10];
  assign isSpecial = T_7 == 2'h3;
  assign T_9 = exp[9];
  assign isNaN = isSpecial & T_9;
  assign notSpecial_magGeOne = exp[11];
  assign T_10 = {notSpecial_magGeOne,fract};
  assign T_11 = exp[5:0];
  assign T_13 = notSpecial_magGeOne ? T_11 : 6'h0;
  assign GEN_0 = {{63'd0}, T_10};
  assign shiftedSig = GEN_0 << T_13;
  assign unroundedInt = shiftedSig[115:52];
  assign T_14 = shiftedSig[52:51];
  assign T_15 = shiftedSig[50:0];
  assign T_17 = T_15 != 51'h0;
  assign roundBits = {T_14,T_17};
  assign T_18 = roundBits[1:0];
  assign T_20 = T_18 != 2'h0;
  assign T_22 = isZero == 1'h0;
  assign roundInexact = notSpecial_magGeOne ? T_20 : T_22;
  assign T_23 = roundBits[2:1];
  assign T_24 = ~ T_23;
  assign T_26 = T_24 == 2'h0;
  assign T_28 = ~ T_18;
  assign T_30 = T_28 == 2'h0;
  assign T_31 = T_26 | T_30;
  assign T_32 = exp[10:0];
  assign T_33 = ~ T_32;
  assign T_35 = T_33 == 11'h0;
  assign T_40 = T_35 ? T_20 : 1'h0;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T_31 : T_40;
  assign T_41 = io_roundingMode == 2'h0;
  assign T_42 = T_41 & roundIncr_nearestEven;
  assign T_43 = io_roundingMode == 2'h2;
  assign T_44 = sign & roundInexact;
  assign T_45 = T_43 & T_44;
  assign T_46 = T_42 | T_45;
  assign T_47 = io_roundingMode == 2'h3;
  assign T_49 = sign == 1'h0;
  assign T_50 = T_49 & roundInexact;
  assign T_51 = T_47 & T_50;
  assign roundIncr = T_46 | T_51;
  assign T_52 = ~ unroundedInt;
  assign complUnroundedInt = sign ? T_52 : unroundedInt;
  assign T_53 = roundIncr ^ sign;
  assign T_55 = complUnroundedInt + 64'h1;
  assign T_56 = T_55[63:0];
  assign roundedInt = T_53 ? T_56 : complUnroundedInt;
  assign T_57 = unroundedInt[61:0];
  assign T_58 = ~ T_57;
  assign T_60 = T_58 == 62'h0;
  assign roundCarryBut2 = T_60 & roundIncr;
  assign T_62 = T_32 >= 11'h40;
  assign T_64 = T_32 == 11'h3f;
  assign T_67 = unroundedInt[62:0];
  assign T_69 = T_67 != 63'h0;
  assign T_70 = T_49 | T_69;
  assign T_71 = T_70 | roundIncr;
  assign T_72 = T_64 & T_71;
  assign T_73 = T_62 | T_72;
  assign T_77 = T_32 == 11'h3e;
  assign T_78 = T_49 & T_77;
  assign T_79 = T_78 & roundCarryBut2;
  assign T_80 = T_73 | T_79;
  assign overflow_signed = notSpecial_magGeOne ? T_80 : 1'h0;
  assign T_84 = sign | T_62;
  assign T_87 = unroundedInt[62];
  assign T_88 = T_64 & T_87;
  assign T_89 = T_88 & roundCarryBut2;
  assign T_90 = T_84 | T_89;
  assign T_91 = sign & roundIncr;
  assign overflow_unsigned = notSpecial_magGeOne ? T_90 : T_91;
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign T_93 = isNaN == 1'h0;
  assign excSign = sign & T_93;
  assign T_94 = io_signedOut & excSign;
  assign T_98 = T_94 ? 64'h8000000000000000 : 64'h0;
  assign T_100 = excSign == 1'h0;
  assign T_101 = io_signedOut & T_100;
  assign T_104 = T_101 ? 63'h7fffffffffffffff : 63'h0;
  assign GEN_1 = {{1'd0}, T_104};
  assign T_105 = T_98 | GEN_1;
  assign T_107 = io_signedOut == 1'h0;
  assign T_110 = T_107 & T_100;
  assign T_113 = T_110 ? 64'hffffffffffffffff : 64'h0;
  assign excValue = T_105 | T_113;
  assign T_115 = isSpecial == 1'h0;
  assign T_116 = roundInexact & T_115;
  assign T_118 = overflow == 1'h0;
  assign inexact = T_116 & T_118;
  assign T_119 = isSpecial | overflow;
  assign T_120 = T_119 ? excValue : roundedInt;
  assign T_121 = {isSpecial,overflow};
  assign T_122 = {T_121,inexact};
endmodule
module FPToInt(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [4:0] io_as_double_cmd,
  output  io_as_double_ldst,
  output  io_as_double_wen,
  output  io_as_double_ren1,
  output  io_as_double_ren2,
  output  io_as_double_ren3,
  output  io_as_double_swap12,
  output  io_as_double_swap23,
  output  io_as_double_single,
  output  io_as_double_fromint,
  output  io_as_double_toint,
  output  io_as_double_fastpipe,
  output  io_as_double_fma,
  output  io_as_double_div,
  output  io_as_double_sqrt,
  output  io_as_double_round,
  output  io_as_double_wflags,
  output [2:0] io_as_double_rm,
  output [1:0] io_as_double_typ,
  output [64:0] io_as_double_in1,
  output [64:0] io_as_double_in2,
  output [64:0] io_as_double_in3,
  output  io_out_valid,
  output  io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0] io_out_bits_exc
);
  reg [4:0] in_cmd;
  reg [31:0] GEN_30;
  reg  in_ldst;
  reg [31:0] GEN_31;
  reg  in_wen;
  reg [31:0] GEN_32;
  reg  in_ren1;
  reg [31:0] GEN_33;
  reg  in_ren2;
  reg [31:0] GEN_34;
  reg  in_ren3;
  reg [31:0] GEN_37;
  reg  in_swap12;
  reg [31:0] GEN_38;
  reg  in_swap23;
  reg [31:0] GEN_39;
  reg  in_single;
  reg [31:0] GEN_40;
  reg  in_fromint;
  reg [31:0] GEN_41;
  reg  in_toint;
  reg [31:0] GEN_47;
  reg  in_fastpipe;
  reg [31:0] GEN_48;
  reg  in_fma;
  reg [31:0] GEN_49;
  reg  in_div;
  reg [31:0] GEN_50;
  reg  in_sqrt;
  reg [31:0] GEN_51;
  reg  in_round;
  reg [31:0] GEN_52;
  reg  in_wflags;
  reg [31:0] GEN_53;
  reg [2:0] in_rm;
  reg [31:0] GEN_54;
  reg [1:0] in_typ;
  reg [31:0] GEN_55;
  reg [64:0] in_in1;
  reg [95:0] GEN_56;
  reg [64:0] in_in2;
  reg [95:0] GEN_57;
  reg [64:0] in_in3;
  reg [95:0] GEN_58;
  reg  valid;
  reg [31:0] GEN_59;
  wire  T_228;
  wire  T_229;
  wire [4:0] T_232;
  wire  T_233;
  wire  T_235;
  wire  T_236;
  wire  T_237;
  wire [22:0] T_238;
  wire [8:0] T_239;
  wire [75:0] GEN_42;
  wire [75:0] T_240;
  wire [51:0] T_241;
  wire [2:0] T_242;
  wire [11:0] GEN_43;
  wire [12:0] T_244;
  wire [11:0] T_245;
  wire [12:0] T_247;
  wire [11:0] T_248;
  wire  T_250;
  wire  T_252;
  wire  T_253;
  wire [8:0] T_254;
  wire [11:0] T_255;
  wire [11:0] T_257;
  wire [12:0] T_258;
  wire [64:0] T_259;
  wire  T_260;
  wire [22:0] T_261;
  wire [8:0] T_262;
  wire [75:0] GEN_44;
  wire [75:0] T_263;
  wire [51:0] T_264;
  wire [2:0] T_265;
  wire [11:0] GEN_45;
  wire [12:0] T_267;
  wire [11:0] T_268;
  wire [12:0] T_270;
  wire [11:0] T_271;
  wire  T_273;
  wire  T_275;
  wire  T_276;
  wire [8:0] T_277;
  wire [11:0] T_278;
  wire [11:0] T_280;
  wire [12:0] T_281;
  wire [64:0] T_282;
  wire [64:0] GEN_0;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  T_283;
  wire [8:0] T_284;
  wire [22:0] T_285;
  wire [6:0] T_286;
  wire  T_288;
  wire [2:0] T_289;
  wire  T_291;
  wire [1:0] T_292;
  wire  T_294;
  wire  T_295;
  wire  T_296;
  wire  T_301;
  wire  T_302;
  wire  T_305;
  wire  T_306;
  wire  T_309;
  wire  T_310;
  wire  T_311;
  wire [4:0] T_313;
  wire [5:0] T_314;
  wire [4:0] T_315;
  wire [23:0] T_317;
  wire [23:0] T_318;
  wire [22:0] T_319;
  wire [7:0] T_320;
  wire [8:0] T_322;
  wire [7:0] T_323;
  wire [7:0] T_327;
  wire [7:0] T_328;
  wire  T_329;
  wire [22:0] T_331;
  wire [22:0] T_332;
  wire [8:0] T_333;
  wire [31:0] T_334;
  wire  T_335;
  wire [31:0] T_339;
  wire [63:0] unrec_s;
  wire  T_340;
  wire [11:0] T_341;
  wire [51:0] T_342;
  wire [9:0] T_343;
  wire  T_345;
  wire [2:0] T_346;
  wire  T_348;
  wire [1:0] T_349;
  wire  T_351;
  wire  T_352;
  wire  T_353;
  wire  T_358;
  wire  T_359;
  wire  T_362;
  wire  T_363;
  wire  T_366;
  wire  T_367;
  wire  T_368;
  wire [5:0] T_370;
  wire [6:0] T_371;
  wire [5:0] T_372;
  wire [52:0] T_374;
  wire [52:0] T_375;
  wire [51:0] T_376;
  wire [10:0] T_377;
  wire [11:0] T_379;
  wire [10:0] T_380;
  wire [10:0] T_384;
  wire [10:0] T_385;
  wire  T_386;
  wire [51:0] T_388;
  wire [51:0] T_389;
  wire [11:0] T_390;
  wire [63:0] T_391;
  wire [63:0] unrec_mem;
  wire [1:0] T_396;
  wire  T_398;
  wire  T_405;
  wire  T_406;
  wire  T_407;
  wire  T_412;
  wire  T_414;
  wire  T_415;
  wire  T_417;
  wire  T_420;
  wire  T_421;
  wire [2:0] T_422;
  wire  T_424;
  wire  T_425;
  wire  T_427;
  wire  T_428;
  wire  T_430;
  wire  T_432;
  wire  T_433;
  wire  T_436;
  wire  T_439;
  wire  T_442;
  wire  T_443;
  wire  T_444;
  wire  T_445;
  wire  T_446;
  wire [1:0] T_447;
  wire [1:0] T_448;
  wire [2:0] T_449;
  wire [4:0] T_450;
  wire [1:0] T_451;
  wire [1:0] T_452;
  wire [2:0] T_453;
  wire [4:0] T_454;
  wire [9:0] classify_s;
  wire [1:0] T_459;
  wire  T_461;
  wire  T_468;
  wire  T_469;
  wire  T_470;
  wire  T_475;
  wire  T_477;
  wire  T_478;
  wire  T_480;
  wire  T_483;
  wire  T_484;
  wire [2:0] T_485;
  wire  T_487;
  wire  T_488;
  wire  T_490;
  wire  T_491;
  wire  T_493;
  wire  T_495;
  wire  T_496;
  wire  T_499;
  wire  T_502;
  wire  T_505;
  wire  T_506;
  wire  T_507;
  wire  T_508;
  wire  T_509;
  wire [1:0] T_510;
  wire [1:0] T_511;
  wire [2:0] T_512;
  wire [4:0] T_513;
  wire [1:0] T_514;
  wire [1:0] T_515;
  wire [2:0] T_516;
  wire [4:0] T_517;
  wire [9:0] T_518;
  wire [9:0] classify_out;
  wire  dcmp_clk;
  wire  dcmp_reset;
  wire [64:0] dcmp_io_a;
  wire [64:0] dcmp_io_b;
  wire  dcmp_io_signaling;
  wire  dcmp_io_lt;
  wire  dcmp_io_eq;
  wire  dcmp_io_gt;
  wire [4:0] dcmp_io_exceptionFlags;
  wire [2:0] T_520;
  wire [1:0] T_521;
  wire [2:0] GEN_46;
  wire [2:0] T_522;
  wire  dcmp_out;
  wire  T_524;
  wire [63:0] T_525;
  wire [4:0] T_529;
  wire  T_530;
  wire [63:0] GEN_24;
  wire [4:0] GEN_25;
  wire  T_534;
  wire  RecFNToIN_2_clk;
  wire  RecFNToIN_2_reset;
  wire [64:0] RecFNToIN_2_io_in;
  wire [1:0] RecFNToIN_2_io_roundingMode;
  wire  RecFNToIN_2_io_signedOut;
  wire [31:0] RecFNToIN_2_io_out;
  wire [2:0] RecFNToIN_2_io_intExceptionFlags;
  wire  T_535;
  wire  T_536;
  wire  T_537;
  wire  T_539;
  wire  T_540;
  wire [31:0] T_544;
  wire [63:0] T_545;
  wire [1:0] T_546;
  wire  T_548;
  wire  T_550;
  wire [3:0] T_551;
  wire [4:0] T_552;
  wire [63:0] GEN_26;
  wire [4:0] GEN_27;
  wire  RecFNToIN_1_1_clk;
  wire  RecFNToIN_1_1_reset;
  wire [64:0] RecFNToIN_1_1_io_in;
  wire [1:0] RecFNToIN_1_1_io_roundingMode;
  wire  RecFNToIN_1_1_io_signedOut;
  wire [63:0] RecFNToIN_1_1_io_out;
  wire [2:0] RecFNToIN_1_1_io_intExceptionFlags;
  wire [1:0] T_558;
  wire  T_560;
  wire  T_562;
  wire [3:0] T_563;
  wire [4:0] T_564;
  wire [63:0] GEN_28;
  wire [4:0] GEN_29;
  wire [63:0] GEN_35;
  wire [4:0] GEN_36;
  CompareRecFN dcmp (
    .clk(dcmp_clk),
    .reset(dcmp_reset),
    .io_a(dcmp_io_a),
    .io_b(dcmp_io_b),
    .io_signaling(dcmp_io_signaling),
    .io_lt(dcmp_io_lt),
    .io_eq(dcmp_io_eq),
    .io_gt(dcmp_io_gt),
    .io_exceptionFlags(dcmp_io_exceptionFlags)
  );
  RecFNToIN RecFNToIN_2 (
    .clk(RecFNToIN_2_clk),
    .reset(RecFNToIN_2_reset),
    .io_in(RecFNToIN_2_io_in),
    .io_roundingMode(RecFNToIN_2_io_roundingMode),
    .io_signedOut(RecFNToIN_2_io_signedOut),
    .io_out(RecFNToIN_2_io_out),
    .io_intExceptionFlags(RecFNToIN_2_io_intExceptionFlags)
  );
  RecFNToIN_1 RecFNToIN_1_1 (
    .clk(RecFNToIN_1_1_clk),
    .reset(RecFNToIN_1_1_reset),
    .io_in(RecFNToIN_1_1_io_in),
    .io_roundingMode(RecFNToIN_1_1_io_roundingMode),
    .io_signedOut(RecFNToIN_1_1_io_signedOut),
    .io_out(RecFNToIN_1_1_io_out),
    .io_intExceptionFlags(RecFNToIN_1_1_io_intExceptionFlags)
  );
  assign io_as_double_cmd = in_cmd;
  assign io_as_double_ldst = in_ldst;
  assign io_as_double_wen = in_wen;
  assign io_as_double_ren1 = in_ren1;
  assign io_as_double_ren2 = in_ren2;
  assign io_as_double_ren3 = in_ren3;
  assign io_as_double_swap12 = in_swap12;
  assign io_as_double_swap23 = in_swap23;
  assign io_as_double_single = in_single;
  assign io_as_double_fromint = in_fromint;
  assign io_as_double_toint = in_toint;
  assign io_as_double_fastpipe = in_fastpipe;
  assign io_as_double_fma = in_fma;
  assign io_as_double_div = in_div;
  assign io_as_double_sqrt = in_sqrt;
  assign io_as_double_round = in_round;
  assign io_as_double_wflags = in_wflags;
  assign io_as_double_rm = in_rm;
  assign io_as_double_typ = in_typ;
  assign io_as_double_in1 = in_in1;
  assign io_as_double_in2 = in_in2;
  assign io_as_double_in3 = in_in3;
  assign io_out_valid = valid;
  assign io_out_bits_lt = dcmp_io_lt;
  assign io_out_bits_store = unrec_mem;
  assign io_out_bits_toint = GEN_35;
  assign io_out_bits_exc = GEN_36;
  assign T_228 = io_in_bits_ldst == 1'h0;
  assign T_229 = io_in_bits_single & T_228;
  assign T_232 = io_in_bits_cmd & 5'hc;
  assign T_233 = 5'hc == T_232;
  assign T_235 = T_233 == 1'h0;
  assign T_236 = T_229 & T_235;
  assign T_237 = io_in_bits_in1[32];
  assign T_238 = io_in_bits_in1[22:0];
  assign T_239 = io_in_bits_in1[31:23];
  assign GEN_42 = {{53'd0}, T_238};
  assign T_240 = GEN_42 << 53;
  assign T_241 = T_240[75:24];
  assign T_242 = T_239[8:6];
  assign GEN_43 = {{3'd0}, T_239};
  assign T_244 = GEN_43 + 12'h800;
  assign T_245 = T_244[11:0];
  assign T_247 = T_245 - 12'h100;
  assign T_248 = T_247[11:0];
  assign T_250 = T_242 == 3'h0;
  assign T_252 = T_242 >= 3'h6;
  assign T_253 = T_250 | T_252;
  assign T_254 = T_248[8:0];
  assign T_255 = {T_242,T_254};
  assign T_257 = T_253 ? T_255 : T_248;
  assign T_258 = {T_237,T_257};
  assign T_259 = {T_258,T_241};
  assign T_260 = io_in_bits_in2[32];
  assign T_261 = io_in_bits_in2[22:0];
  assign T_262 = io_in_bits_in2[31:23];
  assign GEN_44 = {{53'd0}, T_261};
  assign T_263 = GEN_44 << 53;
  assign T_264 = T_263[75:24];
  assign T_265 = T_262[8:6];
  assign GEN_45 = {{3'd0}, T_262};
  assign T_267 = GEN_45 + 12'h800;
  assign T_268 = T_267[11:0];
  assign T_270 = T_268 - 12'h100;
  assign T_271 = T_270[11:0];
  assign T_273 = T_265 == 3'h0;
  assign T_275 = T_265 >= 3'h6;
  assign T_276 = T_273 | T_275;
  assign T_277 = T_271[8:0];
  assign T_278 = {T_265,T_277};
  assign T_280 = T_276 ? T_278 : T_271;
  assign T_281 = {T_260,T_280};
  assign T_282 = {T_281,T_264};
  assign GEN_0 = T_236 ? T_259 : io_in_bits_in1;
  assign GEN_1 = T_236 ? T_282 : io_in_bits_in2;
  assign GEN_2 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? GEN_0 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_1 : in_in2;
  assign GEN_23 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T_283 = in_in1[32];
  assign T_284 = in_in1[31:23];
  assign T_285 = in_in1[22:0];
  assign T_286 = T_284[6:0];
  assign T_288 = T_286 < 7'h2;
  assign T_289 = T_284[8:6];
  assign T_291 = T_289 == 3'h1;
  assign T_292 = T_284[8:7];
  assign T_294 = T_292 == 2'h1;
  assign T_295 = T_294 & T_288;
  assign T_296 = T_291 | T_295;
  assign T_301 = T_288 == 1'h0;
  assign T_302 = T_294 & T_301;
  assign T_305 = T_292 == 2'h2;
  assign T_306 = T_302 | T_305;
  assign T_309 = T_292 == 2'h3;
  assign T_310 = T_284[6];
  assign T_311 = T_309 & T_310;
  assign T_313 = T_284[4:0];
  assign T_314 = 5'h2 - T_313;
  assign T_315 = T_314[4:0];
  assign T_317 = {1'h1,T_285};
  assign T_318 = T_317 >> T_315;
  assign T_319 = T_318[22:0];
  assign T_320 = T_284[7:0];
  assign T_322 = T_320 - 8'h81;
  assign T_323 = T_322[7:0];
  assign T_327 = T_309 ? 8'hff : 8'h0;
  assign T_328 = T_306 ? T_323 : T_327;
  assign T_329 = T_306 | T_311;
  assign T_331 = T_296 ? T_319 : 23'h0;
  assign T_332 = T_329 ? T_285 : T_331;
  assign T_333 = {T_283,T_328};
  assign T_334 = {T_333,T_332};
  assign T_335 = T_334[31];
  assign T_339 = T_335 ? 32'hffffffff : 32'h0;
  assign unrec_s = {T_339,T_334};
  assign T_340 = in_in1[64];
  assign T_341 = in_in1[63:52];
  assign T_342 = in_in1[51:0];
  assign T_343 = T_341[9:0];
  assign T_345 = T_343 < 10'h2;
  assign T_346 = T_341[11:9];
  assign T_348 = T_346 == 3'h1;
  assign T_349 = T_341[11:10];
  assign T_351 = T_349 == 2'h1;
  assign T_352 = T_351 & T_345;
  assign T_353 = T_348 | T_352;
  assign T_358 = T_345 == 1'h0;
  assign T_359 = T_351 & T_358;
  assign T_362 = T_349 == 2'h2;
  assign T_363 = T_359 | T_362;
  assign T_366 = T_349 == 2'h3;
  assign T_367 = T_341[9];
  assign T_368 = T_366 & T_367;
  assign T_370 = T_341[5:0];
  assign T_371 = 6'h2 - T_370;
  assign T_372 = T_371[5:0];
  assign T_374 = {1'h1,T_342};
  assign T_375 = T_374 >> T_372;
  assign T_376 = T_375[51:0];
  assign T_377 = T_341[10:0];
  assign T_379 = T_377 - 11'h401;
  assign T_380 = T_379[10:0];
  assign T_384 = T_366 ? 11'h7ff : 11'h0;
  assign T_385 = T_363 ? T_380 : T_384;
  assign T_386 = T_363 | T_368;
  assign T_388 = T_353 ? T_376 : 52'h0;
  assign T_389 = T_386 ? T_342 : T_388;
  assign T_390 = {T_340,T_385};
  assign T_391 = {T_390,T_389};
  assign unrec_mem = in_single ? unrec_s : T_391;
  assign T_396 = T_289[2:1];
  assign T_398 = T_396 == 2'h3;
  assign T_405 = T_396 == 2'h1;
  assign T_406 = T_405 & T_288;
  assign T_407 = T_291 | T_406;
  assign T_412 = T_405 & T_301;
  assign T_414 = T_396 == 2'h2;
  assign T_415 = T_412 | T_414;
  assign T_417 = T_289 == 3'h0;
  assign T_420 = T_310 == 1'h0;
  assign T_421 = T_398 & T_420;
  assign T_422 = ~ T_289;
  assign T_424 = T_422 == 3'h0;
  assign T_425 = T_285[22];
  assign T_427 = T_425 == 1'h0;
  assign T_428 = T_424 & T_427;
  assign T_430 = T_424 & T_425;
  assign T_432 = T_283 == 1'h0;
  assign T_433 = T_421 & T_432;
  assign T_436 = T_415 & T_432;
  assign T_439 = T_407 & T_432;
  assign T_442 = T_417 & T_432;
  assign T_443 = T_417 & T_283;
  assign T_444 = T_407 & T_283;
  assign T_445 = T_415 & T_283;
  assign T_446 = T_421 & T_283;
  assign T_447 = {T_445,T_446};
  assign T_448 = {T_442,T_443};
  assign T_449 = {T_448,T_444};
  assign T_450 = {T_449,T_447};
  assign T_451 = {T_436,T_439};
  assign T_452 = {T_430,T_428};
  assign T_453 = {T_452,T_433};
  assign T_454 = {T_453,T_451};
  assign classify_s = {T_454,T_450};
  assign T_459 = T_346[2:1];
  assign T_461 = T_459 == 2'h3;
  assign T_468 = T_459 == 2'h1;
  assign T_469 = T_468 & T_345;
  assign T_470 = T_348 | T_469;
  assign T_475 = T_468 & T_358;
  assign T_477 = T_459 == 2'h2;
  assign T_478 = T_475 | T_477;
  assign T_480 = T_346 == 3'h0;
  assign T_483 = T_367 == 1'h0;
  assign T_484 = T_461 & T_483;
  assign T_485 = ~ T_346;
  assign T_487 = T_485 == 3'h0;
  assign T_488 = T_342[51];
  assign T_490 = T_488 == 1'h0;
  assign T_491 = T_487 & T_490;
  assign T_493 = T_487 & T_488;
  assign T_495 = T_340 == 1'h0;
  assign T_496 = T_484 & T_495;
  assign T_499 = T_478 & T_495;
  assign T_502 = T_470 & T_495;
  assign T_505 = T_480 & T_495;
  assign T_506 = T_480 & T_340;
  assign T_507 = T_470 & T_340;
  assign T_508 = T_478 & T_340;
  assign T_509 = T_484 & T_340;
  assign T_510 = {T_508,T_509};
  assign T_511 = {T_505,T_506};
  assign T_512 = {T_511,T_507};
  assign T_513 = {T_512,T_510};
  assign T_514 = {T_499,T_502};
  assign T_515 = {T_493,T_491};
  assign T_516 = {T_515,T_496};
  assign T_517 = {T_516,T_514};
  assign T_518 = {T_517,T_513};
  assign classify_out = in_single ? classify_s : T_518;
  assign dcmp_clk = clk;
  assign dcmp_reset = reset;
  assign dcmp_io_a = in_in1;
  assign dcmp_io_b = in_in2;
  assign dcmp_io_signaling = 1'h1;
  assign T_520 = ~ in_rm;
  assign T_521 = {dcmp_io_lt,dcmp_io_eq};
  assign GEN_46 = {{1'd0}, T_521};
  assign T_522 = T_520 & GEN_46;
  assign dcmp_out = T_522 != 3'h0;
  assign T_524 = in_rm[0];
  assign T_525 = T_524 ? {{54'd0}, classify_out} : unrec_mem;
  assign T_529 = in_cmd & 5'hc;
  assign T_530 = 5'h4 == T_529;
  assign GEN_24 = T_530 ? {{63'd0}, dcmp_out} : T_525;
  assign GEN_25 = T_530 ? dcmp_io_exceptionFlags : 5'h0;
  assign T_534 = 5'h8 == T_529;
  assign RecFNToIN_2_clk = clk;
  assign RecFNToIN_2_reset = reset;
  assign RecFNToIN_2_io_in = in_in1;
  assign RecFNToIN_2_io_roundingMode = in_rm[1:0];
  assign RecFNToIN_2_io_signedOut = T_536;
  assign T_535 = in_typ[0];
  assign T_536 = ~ T_535;
  assign T_537 = in_typ[1];
  assign T_539 = T_537 == 1'h0;
  assign T_540 = RecFNToIN_2_io_out[31];
  assign T_544 = T_540 ? 32'hffffffff : 32'h0;
  assign T_545 = {T_544,RecFNToIN_2_io_out};
  assign T_546 = RecFNToIN_2_io_intExceptionFlags[2:1];
  assign T_548 = T_546 != 2'h0;
  assign T_550 = RecFNToIN_2_io_intExceptionFlags[0];
  assign T_551 = {T_548,3'h0};
  assign T_552 = {T_551,T_550};
  assign GEN_26 = T_539 ? T_545 : GEN_24;
  assign GEN_27 = T_539 ? T_552 : GEN_25;
  assign RecFNToIN_1_1_clk = clk;
  assign RecFNToIN_1_1_reset = reset;
  assign RecFNToIN_1_1_io_in = in_in1;
  assign RecFNToIN_1_1_io_roundingMode = in_rm[1:0];
  assign RecFNToIN_1_1_io_signedOut = T_536;
  assign T_558 = RecFNToIN_1_1_io_intExceptionFlags[2:1];
  assign T_560 = T_558 != 2'h0;
  assign T_562 = RecFNToIN_1_1_io_intExceptionFlags[0];
  assign T_563 = {T_560,3'h0};
  assign T_564 = {T_563,T_562};
  assign GEN_28 = T_537 ? RecFNToIN_1_1_io_out : GEN_26;
  assign GEN_29 = T_537 ? T_564 : GEN_27;
  assign GEN_35 = T_534 ? GEN_28 : GEN_24;
  assign GEN_36 = T_534 ? GEN_29 : GEN_25;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  in_cmd = GEN_30[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  in_ldst = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  in_wen = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  in_ren1 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  in_ren2 = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  in_ren3 = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  in_swap12 = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  in_swap23 = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  in_single = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  in_fromint = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  in_toint = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  in_fastpipe = GEN_48[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  in_fma = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  in_div = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  in_sqrt = GEN_51[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  in_round = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  in_wflags = GEN_53[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  in_rm = GEN_54[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  in_typ = GEN_55[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {3{$random}};
  in_in1 = GEN_56[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {3{$random}};
  in_in2 = GEN_57[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {3{$random}};
  in_in3 = GEN_58[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  valid = GEN_59[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_cmd <= io_in_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ldst <= io_in_bits_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wen <= io_in_bits_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren1 <= io_in_bits_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren2 <= io_in_bits_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren3 <= io_in_bits_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap12 <= io_in_bits_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap23 <= io_in_bits_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_single <= io_in_bits_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fromint <= io_in_bits_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_toint <= io_in_bits_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fastpipe <= io_in_bits_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fma <= io_in_bits_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_div <= io_in_bits_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_sqrt <= io_in_bits_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_round <= io_in_bits_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wflags <= io_in_bits_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_rm <= io_in_bits_rm;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_typ <= io_in_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(T_236) begin
          in_in1 <= T_259;
        end else begin
          in_in1 <= io_in_bits_in1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(T_236) begin
          in_in2 <= T_282;
        end else begin
          in_in2 <= io_in_bits_in2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_in3 <= io_in_bits_in3;
      end
    end
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
  end
endmodule
module INToRecFN(
  input   clk,
  input   reset,
  input   io_signedIn,
  input  [63:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  T_5;
  wire  sign;
  wire [64:0] T_7;
  wire [63:0] T_8;
  wire [63:0] absIn;
  wire [31:0] T_10;
  wire [31:0] T_11;
  wire  T_13;
  wire [15:0] T_14;
  wire [15:0] T_15;
  wire  T_17;
  wire [7:0] T_18;
  wire [7:0] T_19;
  wire  T_21;
  wire [3:0] T_22;
  wire [3:0] T_23;
  wire  T_25;
  wire  T_26;
  wire  T_28;
  wire  T_30;
  wire [1:0] T_32;
  wire [1:0] T_33;
  wire  T_34;
  wire  T_36;
  wire  T_38;
  wire [1:0] T_40;
  wire [1:0] T_41;
  wire [1:0] T_42;
  wire [2:0] T_43;
  wire [3:0] T_44;
  wire [3:0] T_45;
  wire  T_47;
  wire  T_48;
  wire  T_50;
  wire  T_52;
  wire [1:0] T_54;
  wire [1:0] T_55;
  wire  T_56;
  wire  T_58;
  wire  T_60;
  wire [1:0] T_62;
  wire [1:0] T_63;
  wire [1:0] T_64;
  wire [2:0] T_65;
  wire [2:0] T_66;
  wire [3:0] T_67;
  wire [7:0] T_68;
  wire [7:0] T_69;
  wire  T_71;
  wire [3:0] T_72;
  wire [3:0] T_73;
  wire  T_75;
  wire  T_76;
  wire  T_78;
  wire  T_80;
  wire [1:0] T_82;
  wire [1:0] T_83;
  wire  T_84;
  wire  T_86;
  wire  T_88;
  wire [1:0] T_90;
  wire [1:0] T_91;
  wire [1:0] T_92;
  wire [2:0] T_93;
  wire [3:0] T_94;
  wire [3:0] T_95;
  wire  T_97;
  wire  T_98;
  wire  T_100;
  wire  T_102;
  wire [1:0] T_104;
  wire [1:0] T_105;
  wire  T_106;
  wire  T_108;
  wire  T_110;
  wire [1:0] T_112;
  wire [1:0] T_113;
  wire [1:0] T_114;
  wire [2:0] T_115;
  wire [2:0] T_116;
  wire [3:0] T_117;
  wire [3:0] T_118;
  wire [4:0] T_119;
  wire [15:0] T_120;
  wire [15:0] T_121;
  wire  T_123;
  wire [7:0] T_124;
  wire [7:0] T_125;
  wire  T_127;
  wire [3:0] T_128;
  wire [3:0] T_129;
  wire  T_131;
  wire  T_132;
  wire  T_134;
  wire  T_136;
  wire [1:0] T_138;
  wire [1:0] T_139;
  wire  T_140;
  wire  T_142;
  wire  T_144;
  wire [1:0] T_146;
  wire [1:0] T_147;
  wire [1:0] T_148;
  wire [2:0] T_149;
  wire [3:0] T_150;
  wire [3:0] T_151;
  wire  T_153;
  wire  T_154;
  wire  T_156;
  wire  T_158;
  wire [1:0] T_160;
  wire [1:0] T_161;
  wire  T_162;
  wire  T_164;
  wire  T_166;
  wire [1:0] T_168;
  wire [1:0] T_169;
  wire [1:0] T_170;
  wire [2:0] T_171;
  wire [2:0] T_172;
  wire [3:0] T_173;
  wire [7:0] T_174;
  wire [7:0] T_175;
  wire  T_177;
  wire [3:0] T_178;
  wire [3:0] T_179;
  wire  T_181;
  wire  T_182;
  wire  T_184;
  wire  T_186;
  wire [1:0] T_188;
  wire [1:0] T_189;
  wire  T_190;
  wire  T_192;
  wire  T_194;
  wire [1:0] T_196;
  wire [1:0] T_197;
  wire [1:0] T_198;
  wire [2:0] T_199;
  wire [3:0] T_200;
  wire [3:0] T_201;
  wire  T_203;
  wire  T_204;
  wire  T_206;
  wire  T_208;
  wire [1:0] T_210;
  wire [1:0] T_211;
  wire  T_212;
  wire  T_214;
  wire  T_216;
  wire [1:0] T_218;
  wire [1:0] T_219;
  wire [1:0] T_220;
  wire [2:0] T_221;
  wire [2:0] T_222;
  wire [3:0] T_223;
  wire [3:0] T_224;
  wire [4:0] T_225;
  wire [4:0] T_226;
  wire [5:0] T_227;
  wire [5:0] normCount;
  wire [126:0] GEN_0;
  wire [126:0] T_228;
  wire [63:0] normAbsIn;
  wire [1:0] T_230;
  wire [38:0] T_231;
  wire  T_233;
  wire [2:0] roundBits;
  wire [1:0] T_234;
  wire  roundInexact;
  wire  T_236;
  wire [1:0] T_237;
  wire [1:0] T_238;
  wire  T_240;
  wire [1:0] T_242;
  wire  T_244;
  wire  T_245;
  wire  T_247;
  wire  T_248;
  wire  T_249;
  wire  T_251;
  wire  T_252;
  wire  T_253;
  wire  T_255;
  wire  T_256;
  wire  T_258;
  wire  round;
  wire [23:0] T_260;
  wire [24:0] unroundedNorm;
  wire [25:0] T_263;
  wire [24:0] T_264;
  wire [24:0] roundedNorm;
  wire [5:0] T_265;
  wire [6:0] unroundedExp;
  wire [7:0] T_268;
  wire  T_269;
  wire [7:0] GEN_1;
  wire [8:0] T_270;
  wire [7:0] roundedExp;
  wire  T_271;
  wire [8:0] expOut;
  wire [22:0] T_275;
  wire [9:0] T_276;
  wire [32:0] T_277;
  wire [1:0] T_280;
  wire [4:0] T_282;
  assign io_out = T_277;
  assign io_exceptionFlags = T_282;
  assign T_5 = io_in[63];
  assign sign = io_signedIn & T_5;
  assign T_7 = 64'h0 - io_in;
  assign T_8 = T_7[63:0];
  assign absIn = sign ? T_8 : io_in;
  assign T_10 = absIn[63:32];
  assign T_11 = absIn[31:0];
  assign T_13 = T_10 != 32'h0;
  assign T_14 = T_10[31:16];
  assign T_15 = T_10[15:0];
  assign T_17 = T_14 != 16'h0;
  assign T_18 = T_14[15:8];
  assign T_19 = T_14[7:0];
  assign T_21 = T_18 != 8'h0;
  assign T_22 = T_18[7:4];
  assign T_23 = T_18[3:0];
  assign T_25 = T_22 != 4'h0;
  assign T_26 = T_22[3];
  assign T_28 = T_22[2];
  assign T_30 = T_22[1];
  assign T_32 = T_28 ? 2'h2 : {{1'd0}, T_30};
  assign T_33 = T_26 ? 2'h3 : T_32;
  assign T_34 = T_23[3];
  assign T_36 = T_23[2];
  assign T_38 = T_23[1];
  assign T_40 = T_36 ? 2'h2 : {{1'd0}, T_38};
  assign T_41 = T_34 ? 2'h3 : T_40;
  assign T_42 = T_25 ? T_33 : T_41;
  assign T_43 = {T_25,T_42};
  assign T_44 = T_19[7:4];
  assign T_45 = T_19[3:0];
  assign T_47 = T_44 != 4'h0;
  assign T_48 = T_44[3];
  assign T_50 = T_44[2];
  assign T_52 = T_44[1];
  assign T_54 = T_50 ? 2'h2 : {{1'd0}, T_52};
  assign T_55 = T_48 ? 2'h3 : T_54;
  assign T_56 = T_45[3];
  assign T_58 = T_45[2];
  assign T_60 = T_45[1];
  assign T_62 = T_58 ? 2'h2 : {{1'd0}, T_60};
  assign T_63 = T_56 ? 2'h3 : T_62;
  assign T_64 = T_47 ? T_55 : T_63;
  assign T_65 = {T_47,T_64};
  assign T_66 = T_21 ? T_43 : T_65;
  assign T_67 = {T_21,T_66};
  assign T_68 = T_15[15:8];
  assign T_69 = T_15[7:0];
  assign T_71 = T_68 != 8'h0;
  assign T_72 = T_68[7:4];
  assign T_73 = T_68[3:0];
  assign T_75 = T_72 != 4'h0;
  assign T_76 = T_72[3];
  assign T_78 = T_72[2];
  assign T_80 = T_72[1];
  assign T_82 = T_78 ? 2'h2 : {{1'd0}, T_80};
  assign T_83 = T_76 ? 2'h3 : T_82;
  assign T_84 = T_73[3];
  assign T_86 = T_73[2];
  assign T_88 = T_73[1];
  assign T_90 = T_86 ? 2'h2 : {{1'd0}, T_88};
  assign T_91 = T_84 ? 2'h3 : T_90;
  assign T_92 = T_75 ? T_83 : T_91;
  assign T_93 = {T_75,T_92};
  assign T_94 = T_69[7:4];
  assign T_95 = T_69[3:0];
  assign T_97 = T_94 != 4'h0;
  assign T_98 = T_94[3];
  assign T_100 = T_94[2];
  assign T_102 = T_94[1];
  assign T_104 = T_100 ? 2'h2 : {{1'd0}, T_102};
  assign T_105 = T_98 ? 2'h3 : T_104;
  assign T_106 = T_95[3];
  assign T_108 = T_95[2];
  assign T_110 = T_95[1];
  assign T_112 = T_108 ? 2'h2 : {{1'd0}, T_110};
  assign T_113 = T_106 ? 2'h3 : T_112;
  assign T_114 = T_97 ? T_105 : T_113;
  assign T_115 = {T_97,T_114};
  assign T_116 = T_71 ? T_93 : T_115;
  assign T_117 = {T_71,T_116};
  assign T_118 = T_17 ? T_67 : T_117;
  assign T_119 = {T_17,T_118};
  assign T_120 = T_11[31:16];
  assign T_121 = T_11[15:0];
  assign T_123 = T_120 != 16'h0;
  assign T_124 = T_120[15:8];
  assign T_125 = T_120[7:0];
  assign T_127 = T_124 != 8'h0;
  assign T_128 = T_124[7:4];
  assign T_129 = T_124[3:0];
  assign T_131 = T_128 != 4'h0;
  assign T_132 = T_128[3];
  assign T_134 = T_128[2];
  assign T_136 = T_128[1];
  assign T_138 = T_134 ? 2'h2 : {{1'd0}, T_136};
  assign T_139 = T_132 ? 2'h3 : T_138;
  assign T_140 = T_129[3];
  assign T_142 = T_129[2];
  assign T_144 = T_129[1];
  assign T_146 = T_142 ? 2'h2 : {{1'd0}, T_144};
  assign T_147 = T_140 ? 2'h3 : T_146;
  assign T_148 = T_131 ? T_139 : T_147;
  assign T_149 = {T_131,T_148};
  assign T_150 = T_125[7:4];
  assign T_151 = T_125[3:0];
  assign T_153 = T_150 != 4'h0;
  assign T_154 = T_150[3];
  assign T_156 = T_150[2];
  assign T_158 = T_150[1];
  assign T_160 = T_156 ? 2'h2 : {{1'd0}, T_158};
  assign T_161 = T_154 ? 2'h3 : T_160;
  assign T_162 = T_151[3];
  assign T_164 = T_151[2];
  assign T_166 = T_151[1];
  assign T_168 = T_164 ? 2'h2 : {{1'd0}, T_166};
  assign T_169 = T_162 ? 2'h3 : T_168;
  assign T_170 = T_153 ? T_161 : T_169;
  assign T_171 = {T_153,T_170};
  assign T_172 = T_127 ? T_149 : T_171;
  assign T_173 = {T_127,T_172};
  assign T_174 = T_121[15:8];
  assign T_175 = T_121[7:0];
  assign T_177 = T_174 != 8'h0;
  assign T_178 = T_174[7:4];
  assign T_179 = T_174[3:0];
  assign T_181 = T_178 != 4'h0;
  assign T_182 = T_178[3];
  assign T_184 = T_178[2];
  assign T_186 = T_178[1];
  assign T_188 = T_184 ? 2'h2 : {{1'd0}, T_186};
  assign T_189 = T_182 ? 2'h3 : T_188;
  assign T_190 = T_179[3];
  assign T_192 = T_179[2];
  assign T_194 = T_179[1];
  assign T_196 = T_192 ? 2'h2 : {{1'd0}, T_194};
  assign T_197 = T_190 ? 2'h3 : T_196;
  assign T_198 = T_181 ? T_189 : T_197;
  assign T_199 = {T_181,T_198};
  assign T_200 = T_175[7:4];
  assign T_201 = T_175[3:0];
  assign T_203 = T_200 != 4'h0;
  assign T_204 = T_200[3];
  assign T_206 = T_200[2];
  assign T_208 = T_200[1];
  assign T_210 = T_206 ? 2'h2 : {{1'd0}, T_208};
  assign T_211 = T_204 ? 2'h3 : T_210;
  assign T_212 = T_201[3];
  assign T_214 = T_201[2];
  assign T_216 = T_201[1];
  assign T_218 = T_214 ? 2'h2 : {{1'd0}, T_216};
  assign T_219 = T_212 ? 2'h3 : T_218;
  assign T_220 = T_203 ? T_211 : T_219;
  assign T_221 = {T_203,T_220};
  assign T_222 = T_177 ? T_199 : T_221;
  assign T_223 = {T_177,T_222};
  assign T_224 = T_123 ? T_173 : T_223;
  assign T_225 = {T_123,T_224};
  assign T_226 = T_13 ? T_119 : T_225;
  assign T_227 = {T_13,T_226};
  assign normCount = ~ T_227;
  assign GEN_0 = {{63'd0}, absIn};
  assign T_228 = GEN_0 << normCount;
  assign normAbsIn = T_228[63:0];
  assign T_230 = normAbsIn[40:39];
  assign T_231 = normAbsIn[38:0];
  assign T_233 = T_231 != 39'h0;
  assign roundBits = {T_230,T_233};
  assign T_234 = roundBits[1:0];
  assign roundInexact = T_234 != 2'h0;
  assign T_236 = io_roundingMode == 2'h0;
  assign T_237 = roundBits[2:1];
  assign T_238 = ~ T_237;
  assign T_240 = T_238 == 2'h0;
  assign T_242 = ~ T_234;
  assign T_244 = T_242 == 2'h0;
  assign T_245 = T_240 | T_244;
  assign T_247 = T_236 ? T_245 : 1'h0;
  assign T_248 = io_roundingMode == 2'h2;
  assign T_249 = sign & roundInexact;
  assign T_251 = T_248 ? T_249 : 1'h0;
  assign T_252 = T_247 | T_251;
  assign T_253 = io_roundingMode == 2'h3;
  assign T_255 = sign == 1'h0;
  assign T_256 = T_255 & roundInexact;
  assign T_258 = T_253 ? T_256 : 1'h0;
  assign round = T_252 | T_258;
  assign T_260 = normAbsIn[63:40];
  assign unroundedNorm = {1'h0,T_260};
  assign T_263 = unroundedNorm + 25'h1;
  assign T_264 = T_263[24:0];
  assign roundedNorm = round ? T_264 : unroundedNorm;
  assign T_265 = ~ normCount;
  assign unroundedExp = {1'h0,T_265};
  assign T_268 = {1'h0,unroundedExp};
  assign T_269 = roundedNorm[24];
  assign GEN_1 = {{7'd0}, T_269};
  assign T_270 = T_268 + GEN_1;
  assign roundedExp = T_270[7:0];
  assign T_271 = normAbsIn[63];
  assign expOut = {T_271,roundedExp};
  assign T_275 = roundedNorm[22:0];
  assign T_276 = {sign,expOut};
  assign T_277 = {T_276,T_275};
  assign T_280 = {1'h0,roundInexact};
  assign T_282 = {3'h0,T_280};
endmodule
module INToRecFN_1(
  input   clk,
  input   reset,
  input   io_signedIn,
  input  [63:0] io_in,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  T_5;
  wire  sign;
  wire [64:0] T_7;
  wire [63:0] T_8;
  wire [63:0] absIn;
  wire [31:0] T_10;
  wire [31:0] T_11;
  wire  T_13;
  wire [15:0] T_14;
  wire [15:0] T_15;
  wire  T_17;
  wire [7:0] T_18;
  wire [7:0] T_19;
  wire  T_21;
  wire [3:0] T_22;
  wire [3:0] T_23;
  wire  T_25;
  wire  T_26;
  wire  T_28;
  wire  T_30;
  wire [1:0] T_32;
  wire [1:0] T_33;
  wire  T_34;
  wire  T_36;
  wire  T_38;
  wire [1:0] T_40;
  wire [1:0] T_41;
  wire [1:0] T_42;
  wire [2:0] T_43;
  wire [3:0] T_44;
  wire [3:0] T_45;
  wire  T_47;
  wire  T_48;
  wire  T_50;
  wire  T_52;
  wire [1:0] T_54;
  wire [1:0] T_55;
  wire  T_56;
  wire  T_58;
  wire  T_60;
  wire [1:0] T_62;
  wire [1:0] T_63;
  wire [1:0] T_64;
  wire [2:0] T_65;
  wire [2:0] T_66;
  wire [3:0] T_67;
  wire [7:0] T_68;
  wire [7:0] T_69;
  wire  T_71;
  wire [3:0] T_72;
  wire [3:0] T_73;
  wire  T_75;
  wire  T_76;
  wire  T_78;
  wire  T_80;
  wire [1:0] T_82;
  wire [1:0] T_83;
  wire  T_84;
  wire  T_86;
  wire  T_88;
  wire [1:0] T_90;
  wire [1:0] T_91;
  wire [1:0] T_92;
  wire [2:0] T_93;
  wire [3:0] T_94;
  wire [3:0] T_95;
  wire  T_97;
  wire  T_98;
  wire  T_100;
  wire  T_102;
  wire [1:0] T_104;
  wire [1:0] T_105;
  wire  T_106;
  wire  T_108;
  wire  T_110;
  wire [1:0] T_112;
  wire [1:0] T_113;
  wire [1:0] T_114;
  wire [2:0] T_115;
  wire [2:0] T_116;
  wire [3:0] T_117;
  wire [3:0] T_118;
  wire [4:0] T_119;
  wire [15:0] T_120;
  wire [15:0] T_121;
  wire  T_123;
  wire [7:0] T_124;
  wire [7:0] T_125;
  wire  T_127;
  wire [3:0] T_128;
  wire [3:0] T_129;
  wire  T_131;
  wire  T_132;
  wire  T_134;
  wire  T_136;
  wire [1:0] T_138;
  wire [1:0] T_139;
  wire  T_140;
  wire  T_142;
  wire  T_144;
  wire [1:0] T_146;
  wire [1:0] T_147;
  wire [1:0] T_148;
  wire [2:0] T_149;
  wire [3:0] T_150;
  wire [3:0] T_151;
  wire  T_153;
  wire  T_154;
  wire  T_156;
  wire  T_158;
  wire [1:0] T_160;
  wire [1:0] T_161;
  wire  T_162;
  wire  T_164;
  wire  T_166;
  wire [1:0] T_168;
  wire [1:0] T_169;
  wire [1:0] T_170;
  wire [2:0] T_171;
  wire [2:0] T_172;
  wire [3:0] T_173;
  wire [7:0] T_174;
  wire [7:0] T_175;
  wire  T_177;
  wire [3:0] T_178;
  wire [3:0] T_179;
  wire  T_181;
  wire  T_182;
  wire  T_184;
  wire  T_186;
  wire [1:0] T_188;
  wire [1:0] T_189;
  wire  T_190;
  wire  T_192;
  wire  T_194;
  wire [1:0] T_196;
  wire [1:0] T_197;
  wire [1:0] T_198;
  wire [2:0] T_199;
  wire [3:0] T_200;
  wire [3:0] T_201;
  wire  T_203;
  wire  T_204;
  wire  T_206;
  wire  T_208;
  wire [1:0] T_210;
  wire [1:0] T_211;
  wire  T_212;
  wire  T_214;
  wire  T_216;
  wire [1:0] T_218;
  wire [1:0] T_219;
  wire [1:0] T_220;
  wire [2:0] T_221;
  wire [2:0] T_222;
  wire [3:0] T_223;
  wire [3:0] T_224;
  wire [4:0] T_225;
  wire [4:0] T_226;
  wire [5:0] T_227;
  wire [5:0] normCount;
  wire [126:0] GEN_0;
  wire [126:0] T_228;
  wire [63:0] normAbsIn;
  wire [1:0] T_230;
  wire [9:0] T_231;
  wire  T_233;
  wire [2:0] roundBits;
  wire [1:0] T_234;
  wire  roundInexact;
  wire  T_236;
  wire [1:0] T_237;
  wire [1:0] T_238;
  wire  T_240;
  wire [1:0] T_242;
  wire  T_244;
  wire  T_245;
  wire  T_247;
  wire  T_248;
  wire  T_249;
  wire  T_251;
  wire  T_252;
  wire  T_253;
  wire  T_255;
  wire  T_256;
  wire  T_258;
  wire  round;
  wire [52:0] T_260;
  wire [53:0] unroundedNorm;
  wire [54:0] T_263;
  wire [53:0] T_264;
  wire [53:0] roundedNorm;
  wire [5:0] T_265;
  wire [9:0] unroundedExp;
  wire [10:0] T_268;
  wire  T_269;
  wire [10:0] GEN_1;
  wire [11:0] T_270;
  wire [10:0] roundedExp;
  wire  T_271;
  wire [11:0] expOut;
  wire [51:0] T_275;
  wire [12:0] T_276;
  wire [64:0] T_277;
  wire [1:0] T_280;
  wire [4:0] T_282;
  assign io_out = T_277;
  assign io_exceptionFlags = T_282;
  assign T_5 = io_in[63];
  assign sign = io_signedIn & T_5;
  assign T_7 = 64'h0 - io_in;
  assign T_8 = T_7[63:0];
  assign absIn = sign ? T_8 : io_in;
  assign T_10 = absIn[63:32];
  assign T_11 = absIn[31:0];
  assign T_13 = T_10 != 32'h0;
  assign T_14 = T_10[31:16];
  assign T_15 = T_10[15:0];
  assign T_17 = T_14 != 16'h0;
  assign T_18 = T_14[15:8];
  assign T_19 = T_14[7:0];
  assign T_21 = T_18 != 8'h0;
  assign T_22 = T_18[7:4];
  assign T_23 = T_18[3:0];
  assign T_25 = T_22 != 4'h0;
  assign T_26 = T_22[3];
  assign T_28 = T_22[2];
  assign T_30 = T_22[1];
  assign T_32 = T_28 ? 2'h2 : {{1'd0}, T_30};
  assign T_33 = T_26 ? 2'h3 : T_32;
  assign T_34 = T_23[3];
  assign T_36 = T_23[2];
  assign T_38 = T_23[1];
  assign T_40 = T_36 ? 2'h2 : {{1'd0}, T_38};
  assign T_41 = T_34 ? 2'h3 : T_40;
  assign T_42 = T_25 ? T_33 : T_41;
  assign T_43 = {T_25,T_42};
  assign T_44 = T_19[7:4];
  assign T_45 = T_19[3:0];
  assign T_47 = T_44 != 4'h0;
  assign T_48 = T_44[3];
  assign T_50 = T_44[2];
  assign T_52 = T_44[1];
  assign T_54 = T_50 ? 2'h2 : {{1'd0}, T_52};
  assign T_55 = T_48 ? 2'h3 : T_54;
  assign T_56 = T_45[3];
  assign T_58 = T_45[2];
  assign T_60 = T_45[1];
  assign T_62 = T_58 ? 2'h2 : {{1'd0}, T_60};
  assign T_63 = T_56 ? 2'h3 : T_62;
  assign T_64 = T_47 ? T_55 : T_63;
  assign T_65 = {T_47,T_64};
  assign T_66 = T_21 ? T_43 : T_65;
  assign T_67 = {T_21,T_66};
  assign T_68 = T_15[15:8];
  assign T_69 = T_15[7:0];
  assign T_71 = T_68 != 8'h0;
  assign T_72 = T_68[7:4];
  assign T_73 = T_68[3:0];
  assign T_75 = T_72 != 4'h0;
  assign T_76 = T_72[3];
  assign T_78 = T_72[2];
  assign T_80 = T_72[1];
  assign T_82 = T_78 ? 2'h2 : {{1'd0}, T_80};
  assign T_83 = T_76 ? 2'h3 : T_82;
  assign T_84 = T_73[3];
  assign T_86 = T_73[2];
  assign T_88 = T_73[1];
  assign T_90 = T_86 ? 2'h2 : {{1'd0}, T_88};
  assign T_91 = T_84 ? 2'h3 : T_90;
  assign T_92 = T_75 ? T_83 : T_91;
  assign T_93 = {T_75,T_92};
  assign T_94 = T_69[7:4];
  assign T_95 = T_69[3:0];
  assign T_97 = T_94 != 4'h0;
  assign T_98 = T_94[3];
  assign T_100 = T_94[2];
  assign T_102 = T_94[1];
  assign T_104 = T_100 ? 2'h2 : {{1'd0}, T_102};
  assign T_105 = T_98 ? 2'h3 : T_104;
  assign T_106 = T_95[3];
  assign T_108 = T_95[2];
  assign T_110 = T_95[1];
  assign T_112 = T_108 ? 2'h2 : {{1'd0}, T_110};
  assign T_113 = T_106 ? 2'h3 : T_112;
  assign T_114 = T_97 ? T_105 : T_113;
  assign T_115 = {T_97,T_114};
  assign T_116 = T_71 ? T_93 : T_115;
  assign T_117 = {T_71,T_116};
  assign T_118 = T_17 ? T_67 : T_117;
  assign T_119 = {T_17,T_118};
  assign T_120 = T_11[31:16];
  assign T_121 = T_11[15:0];
  assign T_123 = T_120 != 16'h0;
  assign T_124 = T_120[15:8];
  assign T_125 = T_120[7:0];
  assign T_127 = T_124 != 8'h0;
  assign T_128 = T_124[7:4];
  assign T_129 = T_124[3:0];
  assign T_131 = T_128 != 4'h0;
  assign T_132 = T_128[3];
  assign T_134 = T_128[2];
  assign T_136 = T_128[1];
  assign T_138 = T_134 ? 2'h2 : {{1'd0}, T_136};
  assign T_139 = T_132 ? 2'h3 : T_138;
  assign T_140 = T_129[3];
  assign T_142 = T_129[2];
  assign T_144 = T_129[1];
  assign T_146 = T_142 ? 2'h2 : {{1'd0}, T_144};
  assign T_147 = T_140 ? 2'h3 : T_146;
  assign T_148 = T_131 ? T_139 : T_147;
  assign T_149 = {T_131,T_148};
  assign T_150 = T_125[7:4];
  assign T_151 = T_125[3:0];
  assign T_153 = T_150 != 4'h0;
  assign T_154 = T_150[3];
  assign T_156 = T_150[2];
  assign T_158 = T_150[1];
  assign T_160 = T_156 ? 2'h2 : {{1'd0}, T_158};
  assign T_161 = T_154 ? 2'h3 : T_160;
  assign T_162 = T_151[3];
  assign T_164 = T_151[2];
  assign T_166 = T_151[1];
  assign T_168 = T_164 ? 2'h2 : {{1'd0}, T_166};
  assign T_169 = T_162 ? 2'h3 : T_168;
  assign T_170 = T_153 ? T_161 : T_169;
  assign T_171 = {T_153,T_170};
  assign T_172 = T_127 ? T_149 : T_171;
  assign T_173 = {T_127,T_172};
  assign T_174 = T_121[15:8];
  assign T_175 = T_121[7:0];
  assign T_177 = T_174 != 8'h0;
  assign T_178 = T_174[7:4];
  assign T_179 = T_174[3:0];
  assign T_181 = T_178 != 4'h0;
  assign T_182 = T_178[3];
  assign T_184 = T_178[2];
  assign T_186 = T_178[1];
  assign T_188 = T_184 ? 2'h2 : {{1'd0}, T_186};
  assign T_189 = T_182 ? 2'h3 : T_188;
  assign T_190 = T_179[3];
  assign T_192 = T_179[2];
  assign T_194 = T_179[1];
  assign T_196 = T_192 ? 2'h2 : {{1'd0}, T_194};
  assign T_197 = T_190 ? 2'h3 : T_196;
  assign T_198 = T_181 ? T_189 : T_197;
  assign T_199 = {T_181,T_198};
  assign T_200 = T_175[7:4];
  assign T_201 = T_175[3:0];
  assign T_203 = T_200 != 4'h0;
  assign T_204 = T_200[3];
  assign T_206 = T_200[2];
  assign T_208 = T_200[1];
  assign T_210 = T_206 ? 2'h2 : {{1'd0}, T_208};
  assign T_211 = T_204 ? 2'h3 : T_210;
  assign T_212 = T_201[3];
  assign T_214 = T_201[2];
  assign T_216 = T_201[1];
  assign T_218 = T_214 ? 2'h2 : {{1'd0}, T_216};
  assign T_219 = T_212 ? 2'h3 : T_218;
  assign T_220 = T_203 ? T_211 : T_219;
  assign T_221 = {T_203,T_220};
  assign T_222 = T_177 ? T_199 : T_221;
  assign T_223 = {T_177,T_222};
  assign T_224 = T_123 ? T_173 : T_223;
  assign T_225 = {T_123,T_224};
  assign T_226 = T_13 ? T_119 : T_225;
  assign T_227 = {T_13,T_226};
  assign normCount = ~ T_227;
  assign GEN_0 = {{63'd0}, absIn};
  assign T_228 = GEN_0 << normCount;
  assign normAbsIn = T_228[63:0];
  assign T_230 = normAbsIn[11:10];
  assign T_231 = normAbsIn[9:0];
  assign T_233 = T_231 != 10'h0;
  assign roundBits = {T_230,T_233};
  assign T_234 = roundBits[1:0];
  assign roundInexact = T_234 != 2'h0;
  assign T_236 = io_roundingMode == 2'h0;
  assign T_237 = roundBits[2:1];
  assign T_238 = ~ T_237;
  assign T_240 = T_238 == 2'h0;
  assign T_242 = ~ T_234;
  assign T_244 = T_242 == 2'h0;
  assign T_245 = T_240 | T_244;
  assign T_247 = T_236 ? T_245 : 1'h0;
  assign T_248 = io_roundingMode == 2'h2;
  assign T_249 = sign & roundInexact;
  assign T_251 = T_248 ? T_249 : 1'h0;
  assign T_252 = T_247 | T_251;
  assign T_253 = io_roundingMode == 2'h3;
  assign T_255 = sign == 1'h0;
  assign T_256 = T_255 & roundInexact;
  assign T_258 = T_253 ? T_256 : 1'h0;
  assign round = T_252 | T_258;
  assign T_260 = normAbsIn[63:11];
  assign unroundedNorm = {1'h0,T_260};
  assign T_263 = unroundedNorm + 54'h1;
  assign T_264 = T_263[53:0];
  assign roundedNorm = round ? T_264 : unroundedNorm;
  assign T_265 = ~ normCount;
  assign unroundedExp = {4'h0,T_265};
  assign T_268 = {1'h0,unroundedExp};
  assign T_269 = roundedNorm[53];
  assign GEN_1 = {{10'd0}, T_269};
  assign T_270 = T_268 + GEN_1;
  assign roundedExp = T_270[10:0];
  assign T_271 = normAbsIn[63];
  assign expOut = {T_271,roundedExp};
  assign T_275 = roundedNorm[51:0];
  assign T_276 = {sign,expOut};
  assign T_277 = {T_276,T_275};
  assign T_280 = {1'h0,roundInexact};
  assign T_282 = {3'h0,T_280};
endmodule
module IntToFP(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  reg  T_132;
  reg [31:0] GEN_26;
  reg [4:0] T_133_cmd;
  reg [31:0] GEN_27;
  reg  T_133_ldst;
  reg [31:0] GEN_28;
  reg  T_133_wen;
  reg [31:0] GEN_29;
  reg  T_133_ren1;
  reg [31:0] GEN_30;
  reg  T_133_ren2;
  reg [31:0] GEN_33;
  reg  T_133_ren3;
  reg [31:0] GEN_34;
  reg  T_133_swap12;
  reg [31:0] GEN_35;
  reg  T_133_swap23;
  reg [31:0] GEN_36;
  reg  T_133_single;
  reg [31:0] GEN_37;
  reg  T_133_fromint;
  reg [31:0] GEN_56;
  reg  T_133_toint;
  reg [31:0] GEN_57;
  reg  T_133_fastpipe;
  reg [31:0] GEN_58;
  reg  T_133_fma;
  reg [31:0] GEN_59;
  reg  T_133_div;
  reg [31:0] GEN_60;
  reg  T_133_sqrt;
  reg [31:0] GEN_61;
  reg  T_133_round;
  reg [31:0] GEN_62;
  reg  T_133_wflags;
  reg [31:0] GEN_63;
  reg [2:0] T_133_rm;
  reg [31:0] GEN_64;
  reg [1:0] T_133_typ;
  reg [31:0] GEN_65;
  reg [64:0] T_133_in1;
  reg [95:0] GEN_66;
  reg [64:0] T_133_in2;
  reg [95:0] GEN_67;
  reg [64:0] T_133_in3;
  reg [95:0] GEN_68;
  wire [4:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire [64:0] GEN_19;
  wire [64:0] GEN_20;
  wire [64:0] GEN_21;
  wire  in_valid;
  wire [4:0] in_bits_cmd;
  wire  in_bits_ldst;
  wire  in_bits_wen;
  wire  in_bits_ren1;
  wire  in_bits_ren2;
  wire  in_bits_ren3;
  wire  in_bits_swap12;
  wire  in_bits_swap23;
  wire  in_bits_single;
  wire  in_bits_fromint;
  wire  in_bits_toint;
  wire  in_bits_fastpipe;
  wire  in_bits_fma;
  wire  in_bits_div;
  wire  in_bits_sqrt;
  wire  in_bits_round;
  wire  in_bits_wflags;
  wire [2:0] in_bits_rm;
  wire [1:0] in_bits_typ;
  wire [64:0] in_bits_in1;
  wire [64:0] in_bits_in2;
  wire [64:0] in_bits_in3;
  wire [64:0] mux_data;
  wire [4:0] mux_exc;
  wire  T_257;
  wire [7:0] T_258;
  wire [22:0] T_259;
  wire  T_261;
  wire  T_263;
  wire  T_264;
  wire [31:0] GEN_40;
  wire [31:0] T_265;
  wire [15:0] T_266;
  wire [15:0] T_267;
  wire  T_269;
  wire [7:0] T_270;
  wire [7:0] T_271;
  wire  T_273;
  wire [3:0] T_274;
  wire [3:0] T_275;
  wire  T_277;
  wire  T_278;
  wire  T_280;
  wire  T_282;
  wire [1:0] T_284;
  wire [1:0] T_285;
  wire  T_286;
  wire  T_288;
  wire  T_290;
  wire [1:0] T_292;
  wire [1:0] T_293;
  wire [1:0] T_294;
  wire [2:0] T_295;
  wire [3:0] T_296;
  wire [3:0] T_297;
  wire  T_299;
  wire  T_300;
  wire  T_302;
  wire  T_304;
  wire [1:0] T_306;
  wire [1:0] T_307;
  wire  T_308;
  wire  T_310;
  wire  T_312;
  wire [1:0] T_314;
  wire [1:0] T_315;
  wire [1:0] T_316;
  wire [2:0] T_317;
  wire [2:0] T_318;
  wire [3:0] T_319;
  wire [7:0] T_320;
  wire [7:0] T_321;
  wire  T_323;
  wire [3:0] T_324;
  wire [3:0] T_325;
  wire  T_327;
  wire  T_328;
  wire  T_330;
  wire  T_332;
  wire [1:0] T_334;
  wire [1:0] T_335;
  wire  T_336;
  wire  T_338;
  wire  T_340;
  wire [1:0] T_342;
  wire [1:0] T_343;
  wire [1:0] T_344;
  wire [2:0] T_345;
  wire [3:0] T_346;
  wire [3:0] T_347;
  wire  T_349;
  wire  T_350;
  wire  T_352;
  wire  T_354;
  wire [1:0] T_356;
  wire [1:0] T_357;
  wire  T_358;
  wire  T_360;
  wire  T_362;
  wire [1:0] T_364;
  wire [1:0] T_365;
  wire [1:0] T_366;
  wire [2:0] T_367;
  wire [2:0] T_368;
  wire [3:0] T_369;
  wire [3:0] T_370;
  wire [4:0] T_371;
  wire [4:0] T_372;
  wire [53:0] GEN_41;
  wire [53:0] T_373;
  wire [21:0] T_374;
  wire [22:0] T_376;
  wire [8:0] GEN_42;
  wire [8:0] T_382;
  wire [8:0] T_383;
  wire [1:0] T_387;
  wire [7:0] GEN_43;
  wire [7:0] T_388;
  wire [8:0] GEN_44;
  wire [9:0] T_389;
  wire [8:0] T_390;
  wire [1:0] T_391;
  wire  T_393;
  wire  T_395;
  wire  T_396;
  wire [2:0] T_400;
  wire [8:0] GEN_45;
  wire [8:0] T_401;
  wire [8:0] T_402;
  wire [8:0] T_403;
  wire [6:0] GEN_46;
  wire [6:0] T_404;
  wire [8:0] GEN_47;
  wire [8:0] T_405;
  wire [22:0] T_406;
  wire [9:0] T_407;
  wire [32:0] T_408;
  wire  T_410;
  wire  T_411;
  wire [10:0] T_412;
  wire [51:0] T_413;
  wire  T_415;
  wire  T_417;
  wire  T_418;
  wire [63:0] GEN_48;
  wire [63:0] T_419;
  wire [31:0] T_420;
  wire [31:0] T_421;
  wire  T_423;
  wire [15:0] T_424;
  wire [15:0] T_425;
  wire  T_427;
  wire [7:0] T_428;
  wire [7:0] T_429;
  wire  T_431;
  wire [3:0] T_432;
  wire [3:0] T_433;
  wire  T_435;
  wire  T_436;
  wire  T_438;
  wire  T_440;
  wire [1:0] T_442;
  wire [1:0] T_443;
  wire  T_444;
  wire  T_446;
  wire  T_448;
  wire [1:0] T_450;
  wire [1:0] T_451;
  wire [1:0] T_452;
  wire [2:0] T_453;
  wire [3:0] T_454;
  wire [3:0] T_455;
  wire  T_457;
  wire  T_458;
  wire  T_460;
  wire  T_462;
  wire [1:0] T_464;
  wire [1:0] T_465;
  wire  T_466;
  wire  T_468;
  wire  T_470;
  wire [1:0] T_472;
  wire [1:0] T_473;
  wire [1:0] T_474;
  wire [2:0] T_475;
  wire [2:0] T_476;
  wire [3:0] T_477;
  wire [7:0] T_478;
  wire [7:0] T_479;
  wire  T_481;
  wire [3:0] T_482;
  wire [3:0] T_483;
  wire  T_485;
  wire  T_486;
  wire  T_488;
  wire  T_490;
  wire [1:0] T_492;
  wire [1:0] T_493;
  wire  T_494;
  wire  T_496;
  wire  T_498;
  wire [1:0] T_500;
  wire [1:0] T_501;
  wire [1:0] T_502;
  wire [2:0] T_503;
  wire [3:0] T_504;
  wire [3:0] T_505;
  wire  T_507;
  wire  T_508;
  wire  T_510;
  wire  T_512;
  wire [1:0] T_514;
  wire [1:0] T_515;
  wire  T_516;
  wire  T_518;
  wire  T_520;
  wire [1:0] T_522;
  wire [1:0] T_523;
  wire [1:0] T_524;
  wire [2:0] T_525;
  wire [2:0] T_526;
  wire [3:0] T_527;
  wire [3:0] T_528;
  wire [4:0] T_529;
  wire [15:0] T_530;
  wire [15:0] T_531;
  wire  T_533;
  wire [7:0] T_534;
  wire [7:0] T_535;
  wire  T_537;
  wire [3:0] T_538;
  wire [3:0] T_539;
  wire  T_541;
  wire  T_542;
  wire  T_544;
  wire  T_546;
  wire [1:0] T_548;
  wire [1:0] T_549;
  wire  T_550;
  wire  T_552;
  wire  T_554;
  wire [1:0] T_556;
  wire [1:0] T_557;
  wire [1:0] T_558;
  wire [2:0] T_559;
  wire [3:0] T_560;
  wire [3:0] T_561;
  wire  T_563;
  wire  T_564;
  wire  T_566;
  wire  T_568;
  wire [1:0] T_570;
  wire [1:0] T_571;
  wire  T_572;
  wire  T_574;
  wire  T_576;
  wire [1:0] T_578;
  wire [1:0] T_579;
  wire [1:0] T_580;
  wire [2:0] T_581;
  wire [2:0] T_582;
  wire [3:0] T_583;
  wire [7:0] T_584;
  wire [7:0] T_585;
  wire  T_587;
  wire [3:0] T_588;
  wire [3:0] T_589;
  wire  T_591;
  wire  T_592;
  wire  T_594;
  wire  T_596;
  wire [1:0] T_598;
  wire [1:0] T_599;
  wire  T_600;
  wire  T_602;
  wire  T_604;
  wire [1:0] T_606;
  wire [1:0] T_607;
  wire [1:0] T_608;
  wire [2:0] T_609;
  wire [3:0] T_610;
  wire [3:0] T_611;
  wire  T_613;
  wire  T_614;
  wire  T_616;
  wire  T_618;
  wire [1:0] T_620;
  wire [1:0] T_621;
  wire  T_622;
  wire  T_624;
  wire  T_626;
  wire [1:0] T_628;
  wire [1:0] T_629;
  wire [1:0] T_630;
  wire [2:0] T_631;
  wire [2:0] T_632;
  wire [3:0] T_633;
  wire [3:0] T_634;
  wire [4:0] T_635;
  wire [4:0] T_636;
  wire [5:0] T_637;
  wire [5:0] T_638;
  wire [114:0] GEN_49;
  wire [114:0] T_639;
  wire [50:0] T_640;
  wire [51:0] T_642;
  wire [11:0] GEN_50;
  wire [11:0] T_648;
  wire [11:0] T_649;
  wire [1:0] T_653;
  wire [10:0] GEN_51;
  wire [10:0] T_654;
  wire [11:0] GEN_52;
  wire [12:0] T_655;
  wire [11:0] T_656;
  wire [1:0] T_657;
  wire  T_659;
  wire  T_661;
  wire  T_662;
  wire [2:0] T_666;
  wire [11:0] GEN_53;
  wire [11:0] T_667;
  wire [11:0] T_668;
  wire [11:0] T_669;
  wire [9:0] GEN_54;
  wire [9:0] T_670;
  wire [11:0] GEN_55;
  wire [11:0] T_671;
  wire [51:0] T_672;
  wire [12:0] T_673;
  wire [64:0] T_674;
  wire [64:0] GEN_22;
  wire [64:0] T_675;
  wire [64:0] T_676;
  wire [31:0] T_677;
  wire  T_678;
  wire  T_680;
  wire  T_681;
  wire [32:0] T_682;
  wire [31:0] T_683;
  wire [32:0] T_684;
  wire [64:0] GEN_23;
  wire [64:0] intValue;
  wire [4:0] T_687;
  wire  T_688;
  wire  INToRecFN_2_clk;
  wire  INToRecFN_2_reset;
  wire  INToRecFN_2_io_signedIn;
  wire [63:0] INToRecFN_2_io_in;
  wire [1:0] INToRecFN_2_io_roundingMode;
  wire [32:0] INToRecFN_2_io_out;
  wire [4:0] INToRecFN_2_io_exceptionFlags;
  wire  T_690;
  wire [64:0] T_692;
  wire  INToRecFN_1_1_clk;
  wire  INToRecFN_1_1_reset;
  wire  INToRecFN_1_1_io_signedIn;
  wire [63:0] INToRecFN_1_1_io_in;
  wire [1:0] INToRecFN_1_1_io_roundingMode;
  wire [64:0] INToRecFN_1_1_io_out;
  wire [4:0] INToRecFN_1_1_io_exceptionFlags;
  wire [65:0] T_698;
  wire [65:0] GEN_24;
  wire [4:0] GEN_25;
  wire [65:0] GEN_31;
  wire [4:0] GEN_32;
  reg  T_701;
  reg [31:0] GEN_69;
  reg [64:0] T_702_data;
  reg [95:0] GEN_70;
  reg [4:0] T_702_exc;
  reg [31:0] GEN_71;
  wire [64:0] GEN_38;
  wire [4:0] GEN_39;
  wire  T_713_valid;
  wire [64:0] T_713_bits_data;
  wire [4:0] T_713_bits_exc;
  INToRecFN INToRecFN_2 (
    .clk(INToRecFN_2_clk),
    .reset(INToRecFN_2_reset),
    .io_signedIn(INToRecFN_2_io_signedIn),
    .io_in(INToRecFN_2_io_in),
    .io_roundingMode(INToRecFN_2_io_roundingMode),
    .io_out(INToRecFN_2_io_out),
    .io_exceptionFlags(INToRecFN_2_io_exceptionFlags)
  );
  INToRecFN_1 INToRecFN_1_1 (
    .clk(INToRecFN_1_1_clk),
    .reset(INToRecFN_1_1_reset),
    .io_signedIn(INToRecFN_1_1_io_signedIn),
    .io_in(INToRecFN_1_1_io_in),
    .io_roundingMode(INToRecFN_1_1_io_roundingMode),
    .io_out(INToRecFN_1_1_io_out),
    .io_exceptionFlags(INToRecFN_1_1_io_exceptionFlags)
  );
  assign io_out_valid = T_713_valid;
  assign io_out_bits_data = T_713_bits_data;
  assign io_out_bits_exc = T_713_bits_exc;
  assign GEN_0 = io_in_valid ? io_in_bits_cmd : T_133_cmd;
  assign GEN_1 = io_in_valid ? io_in_bits_ldst : T_133_ldst;
  assign GEN_2 = io_in_valid ? io_in_bits_wen : T_133_wen;
  assign GEN_3 = io_in_valid ? io_in_bits_ren1 : T_133_ren1;
  assign GEN_4 = io_in_valid ? io_in_bits_ren2 : T_133_ren2;
  assign GEN_5 = io_in_valid ? io_in_bits_ren3 : T_133_ren3;
  assign GEN_6 = io_in_valid ? io_in_bits_swap12 : T_133_swap12;
  assign GEN_7 = io_in_valid ? io_in_bits_swap23 : T_133_swap23;
  assign GEN_8 = io_in_valid ? io_in_bits_single : T_133_single;
  assign GEN_9 = io_in_valid ? io_in_bits_fromint : T_133_fromint;
  assign GEN_10 = io_in_valid ? io_in_bits_toint : T_133_toint;
  assign GEN_11 = io_in_valid ? io_in_bits_fastpipe : T_133_fastpipe;
  assign GEN_12 = io_in_valid ? io_in_bits_fma : T_133_fma;
  assign GEN_13 = io_in_valid ? io_in_bits_div : T_133_div;
  assign GEN_14 = io_in_valid ? io_in_bits_sqrt : T_133_sqrt;
  assign GEN_15 = io_in_valid ? io_in_bits_round : T_133_round;
  assign GEN_16 = io_in_valid ? io_in_bits_wflags : T_133_wflags;
  assign GEN_17 = io_in_valid ? io_in_bits_rm : T_133_rm;
  assign GEN_18 = io_in_valid ? io_in_bits_typ : T_133_typ;
  assign GEN_19 = io_in_valid ? io_in_bits_in1 : T_133_in1;
  assign GEN_20 = io_in_valid ? io_in_bits_in2 : T_133_in2;
  assign GEN_21 = io_in_valid ? io_in_bits_in3 : T_133_in3;
  assign in_valid = T_132;
  assign in_bits_cmd = T_133_cmd;
  assign in_bits_ldst = T_133_ldst;
  assign in_bits_wen = T_133_wen;
  assign in_bits_ren1 = T_133_ren1;
  assign in_bits_ren2 = T_133_ren2;
  assign in_bits_ren3 = T_133_ren3;
  assign in_bits_swap12 = T_133_swap12;
  assign in_bits_swap23 = T_133_swap23;
  assign in_bits_single = T_133_single;
  assign in_bits_fromint = T_133_fromint;
  assign in_bits_toint = T_133_toint;
  assign in_bits_fastpipe = T_133_fastpipe;
  assign in_bits_fma = T_133_fma;
  assign in_bits_div = T_133_div;
  assign in_bits_sqrt = T_133_sqrt;
  assign in_bits_round = T_133_round;
  assign in_bits_wflags = T_133_wflags;
  assign in_bits_rm = T_133_rm;
  assign in_bits_typ = T_133_typ;
  assign in_bits_in1 = T_133_in1;
  assign in_bits_in2 = T_133_in2;
  assign in_bits_in3 = T_133_in3;
  assign mux_data = GEN_31[64:0];
  assign mux_exc = GEN_32;
  assign T_257 = in_bits_in1[31];
  assign T_258 = in_bits_in1[30:23];
  assign T_259 = in_bits_in1[22:0];
  assign T_261 = T_258 == 8'h0;
  assign T_263 = T_259 == 23'h0;
  assign T_264 = T_261 & T_263;
  assign GEN_40 = {{9'd0}, T_259};
  assign T_265 = GEN_40 << 9;
  assign T_266 = T_265[31:16];
  assign T_267 = T_265[15:0];
  assign T_269 = T_266 != 16'h0;
  assign T_270 = T_266[15:8];
  assign T_271 = T_266[7:0];
  assign T_273 = T_270 != 8'h0;
  assign T_274 = T_270[7:4];
  assign T_275 = T_270[3:0];
  assign T_277 = T_274 != 4'h0;
  assign T_278 = T_274[3];
  assign T_280 = T_274[2];
  assign T_282 = T_274[1];
  assign T_284 = T_280 ? 2'h2 : {{1'd0}, T_282};
  assign T_285 = T_278 ? 2'h3 : T_284;
  assign T_286 = T_275[3];
  assign T_288 = T_275[2];
  assign T_290 = T_275[1];
  assign T_292 = T_288 ? 2'h2 : {{1'd0}, T_290};
  assign T_293 = T_286 ? 2'h3 : T_292;
  assign T_294 = T_277 ? T_285 : T_293;
  assign T_295 = {T_277,T_294};
  assign T_296 = T_271[7:4];
  assign T_297 = T_271[3:0];
  assign T_299 = T_296 != 4'h0;
  assign T_300 = T_296[3];
  assign T_302 = T_296[2];
  assign T_304 = T_296[1];
  assign T_306 = T_302 ? 2'h2 : {{1'd0}, T_304};
  assign T_307 = T_300 ? 2'h3 : T_306;
  assign T_308 = T_297[3];
  assign T_310 = T_297[2];
  assign T_312 = T_297[1];
  assign T_314 = T_310 ? 2'h2 : {{1'd0}, T_312};
  assign T_315 = T_308 ? 2'h3 : T_314;
  assign T_316 = T_299 ? T_307 : T_315;
  assign T_317 = {T_299,T_316};
  assign T_318 = T_273 ? T_295 : T_317;
  assign T_319 = {T_273,T_318};
  assign T_320 = T_267[15:8];
  assign T_321 = T_267[7:0];
  assign T_323 = T_320 != 8'h0;
  assign T_324 = T_320[7:4];
  assign T_325 = T_320[3:0];
  assign T_327 = T_324 != 4'h0;
  assign T_328 = T_324[3];
  assign T_330 = T_324[2];
  assign T_332 = T_324[1];
  assign T_334 = T_330 ? 2'h2 : {{1'd0}, T_332};
  assign T_335 = T_328 ? 2'h3 : T_334;
  assign T_336 = T_325[3];
  assign T_338 = T_325[2];
  assign T_340 = T_325[1];
  assign T_342 = T_338 ? 2'h2 : {{1'd0}, T_340};
  assign T_343 = T_336 ? 2'h3 : T_342;
  assign T_344 = T_327 ? T_335 : T_343;
  assign T_345 = {T_327,T_344};
  assign T_346 = T_321[7:4];
  assign T_347 = T_321[3:0];
  assign T_349 = T_346 != 4'h0;
  assign T_350 = T_346[3];
  assign T_352 = T_346[2];
  assign T_354 = T_346[1];
  assign T_356 = T_352 ? 2'h2 : {{1'd0}, T_354};
  assign T_357 = T_350 ? 2'h3 : T_356;
  assign T_358 = T_347[3];
  assign T_360 = T_347[2];
  assign T_362 = T_347[1];
  assign T_364 = T_360 ? 2'h2 : {{1'd0}, T_362};
  assign T_365 = T_358 ? 2'h3 : T_364;
  assign T_366 = T_349 ? T_357 : T_365;
  assign T_367 = {T_349,T_366};
  assign T_368 = T_323 ? T_345 : T_367;
  assign T_369 = {T_323,T_368};
  assign T_370 = T_269 ? T_319 : T_369;
  assign T_371 = {T_269,T_370};
  assign T_372 = ~ T_371;
  assign GEN_41 = {{31'd0}, T_259};
  assign T_373 = GEN_41 << T_372;
  assign T_374 = T_373[21:0];
  assign T_376 = {T_374,1'h0};
  assign GEN_42 = {{4'd0}, T_372};
  assign T_382 = GEN_42 ^ 9'h1ff;
  assign T_383 = T_261 ? T_382 : {{1'd0}, T_258};
  assign T_387 = T_261 ? 2'h2 : 2'h1;
  assign GEN_43 = {{6'd0}, T_387};
  assign T_388 = 8'h80 | GEN_43;
  assign GEN_44 = {{1'd0}, T_388};
  assign T_389 = T_383 + GEN_44;
  assign T_390 = T_389[8:0];
  assign T_391 = T_390[8:7];
  assign T_393 = T_391 == 2'h3;
  assign T_395 = T_263 == 1'h0;
  assign T_396 = T_393 & T_395;
  assign T_400 = T_264 ? 3'h7 : 3'h0;
  assign GEN_45 = {{6'd0}, T_400};
  assign T_401 = GEN_45 << 6;
  assign T_402 = ~ T_401;
  assign T_403 = T_390 & T_402;
  assign GEN_46 = {{6'd0}, T_396};
  assign T_404 = GEN_46 << 6;
  assign GEN_47 = {{2'd0}, T_404};
  assign T_405 = T_403 | GEN_47;
  assign T_406 = T_261 ? T_376 : T_259;
  assign T_407 = {T_257,T_405};
  assign T_408 = {T_407,T_406};
  assign T_410 = in_bits_single == 1'h0;
  assign T_411 = in_bits_in1[63];
  assign T_412 = in_bits_in1[62:52];
  assign T_413 = in_bits_in1[51:0];
  assign T_415 = T_412 == 11'h0;
  assign T_417 = T_413 == 52'h0;
  assign T_418 = T_415 & T_417;
  assign GEN_48 = {{12'd0}, T_413};
  assign T_419 = GEN_48 << 12;
  assign T_420 = T_419[63:32];
  assign T_421 = T_419[31:0];
  assign T_423 = T_420 != 32'h0;
  assign T_424 = T_420[31:16];
  assign T_425 = T_420[15:0];
  assign T_427 = T_424 != 16'h0;
  assign T_428 = T_424[15:8];
  assign T_429 = T_424[7:0];
  assign T_431 = T_428 != 8'h0;
  assign T_432 = T_428[7:4];
  assign T_433 = T_428[3:0];
  assign T_435 = T_432 != 4'h0;
  assign T_436 = T_432[3];
  assign T_438 = T_432[2];
  assign T_440 = T_432[1];
  assign T_442 = T_438 ? 2'h2 : {{1'd0}, T_440};
  assign T_443 = T_436 ? 2'h3 : T_442;
  assign T_444 = T_433[3];
  assign T_446 = T_433[2];
  assign T_448 = T_433[1];
  assign T_450 = T_446 ? 2'h2 : {{1'd0}, T_448};
  assign T_451 = T_444 ? 2'h3 : T_450;
  assign T_452 = T_435 ? T_443 : T_451;
  assign T_453 = {T_435,T_452};
  assign T_454 = T_429[7:4];
  assign T_455 = T_429[3:0];
  assign T_457 = T_454 != 4'h0;
  assign T_458 = T_454[3];
  assign T_460 = T_454[2];
  assign T_462 = T_454[1];
  assign T_464 = T_460 ? 2'h2 : {{1'd0}, T_462};
  assign T_465 = T_458 ? 2'h3 : T_464;
  assign T_466 = T_455[3];
  assign T_468 = T_455[2];
  assign T_470 = T_455[1];
  assign T_472 = T_468 ? 2'h2 : {{1'd0}, T_470};
  assign T_473 = T_466 ? 2'h3 : T_472;
  assign T_474 = T_457 ? T_465 : T_473;
  assign T_475 = {T_457,T_474};
  assign T_476 = T_431 ? T_453 : T_475;
  assign T_477 = {T_431,T_476};
  assign T_478 = T_425[15:8];
  assign T_479 = T_425[7:0];
  assign T_481 = T_478 != 8'h0;
  assign T_482 = T_478[7:4];
  assign T_483 = T_478[3:0];
  assign T_485 = T_482 != 4'h0;
  assign T_486 = T_482[3];
  assign T_488 = T_482[2];
  assign T_490 = T_482[1];
  assign T_492 = T_488 ? 2'h2 : {{1'd0}, T_490};
  assign T_493 = T_486 ? 2'h3 : T_492;
  assign T_494 = T_483[3];
  assign T_496 = T_483[2];
  assign T_498 = T_483[1];
  assign T_500 = T_496 ? 2'h2 : {{1'd0}, T_498};
  assign T_501 = T_494 ? 2'h3 : T_500;
  assign T_502 = T_485 ? T_493 : T_501;
  assign T_503 = {T_485,T_502};
  assign T_504 = T_479[7:4];
  assign T_505 = T_479[3:0];
  assign T_507 = T_504 != 4'h0;
  assign T_508 = T_504[3];
  assign T_510 = T_504[2];
  assign T_512 = T_504[1];
  assign T_514 = T_510 ? 2'h2 : {{1'd0}, T_512};
  assign T_515 = T_508 ? 2'h3 : T_514;
  assign T_516 = T_505[3];
  assign T_518 = T_505[2];
  assign T_520 = T_505[1];
  assign T_522 = T_518 ? 2'h2 : {{1'd0}, T_520};
  assign T_523 = T_516 ? 2'h3 : T_522;
  assign T_524 = T_507 ? T_515 : T_523;
  assign T_525 = {T_507,T_524};
  assign T_526 = T_481 ? T_503 : T_525;
  assign T_527 = {T_481,T_526};
  assign T_528 = T_427 ? T_477 : T_527;
  assign T_529 = {T_427,T_528};
  assign T_530 = T_421[31:16];
  assign T_531 = T_421[15:0];
  assign T_533 = T_530 != 16'h0;
  assign T_534 = T_530[15:8];
  assign T_535 = T_530[7:0];
  assign T_537 = T_534 != 8'h0;
  assign T_538 = T_534[7:4];
  assign T_539 = T_534[3:0];
  assign T_541 = T_538 != 4'h0;
  assign T_542 = T_538[3];
  assign T_544 = T_538[2];
  assign T_546 = T_538[1];
  assign T_548 = T_544 ? 2'h2 : {{1'd0}, T_546};
  assign T_549 = T_542 ? 2'h3 : T_548;
  assign T_550 = T_539[3];
  assign T_552 = T_539[2];
  assign T_554 = T_539[1];
  assign T_556 = T_552 ? 2'h2 : {{1'd0}, T_554};
  assign T_557 = T_550 ? 2'h3 : T_556;
  assign T_558 = T_541 ? T_549 : T_557;
  assign T_559 = {T_541,T_558};
  assign T_560 = T_535[7:4];
  assign T_561 = T_535[3:0];
  assign T_563 = T_560 != 4'h0;
  assign T_564 = T_560[3];
  assign T_566 = T_560[2];
  assign T_568 = T_560[1];
  assign T_570 = T_566 ? 2'h2 : {{1'd0}, T_568};
  assign T_571 = T_564 ? 2'h3 : T_570;
  assign T_572 = T_561[3];
  assign T_574 = T_561[2];
  assign T_576 = T_561[1];
  assign T_578 = T_574 ? 2'h2 : {{1'd0}, T_576};
  assign T_579 = T_572 ? 2'h3 : T_578;
  assign T_580 = T_563 ? T_571 : T_579;
  assign T_581 = {T_563,T_580};
  assign T_582 = T_537 ? T_559 : T_581;
  assign T_583 = {T_537,T_582};
  assign T_584 = T_531[15:8];
  assign T_585 = T_531[7:0];
  assign T_587 = T_584 != 8'h0;
  assign T_588 = T_584[7:4];
  assign T_589 = T_584[3:0];
  assign T_591 = T_588 != 4'h0;
  assign T_592 = T_588[3];
  assign T_594 = T_588[2];
  assign T_596 = T_588[1];
  assign T_598 = T_594 ? 2'h2 : {{1'd0}, T_596};
  assign T_599 = T_592 ? 2'h3 : T_598;
  assign T_600 = T_589[3];
  assign T_602 = T_589[2];
  assign T_604 = T_589[1];
  assign T_606 = T_602 ? 2'h2 : {{1'd0}, T_604};
  assign T_607 = T_600 ? 2'h3 : T_606;
  assign T_608 = T_591 ? T_599 : T_607;
  assign T_609 = {T_591,T_608};
  assign T_610 = T_585[7:4];
  assign T_611 = T_585[3:0];
  assign T_613 = T_610 != 4'h0;
  assign T_614 = T_610[3];
  assign T_616 = T_610[2];
  assign T_618 = T_610[1];
  assign T_620 = T_616 ? 2'h2 : {{1'd0}, T_618};
  assign T_621 = T_614 ? 2'h3 : T_620;
  assign T_622 = T_611[3];
  assign T_624 = T_611[2];
  assign T_626 = T_611[1];
  assign T_628 = T_624 ? 2'h2 : {{1'd0}, T_626};
  assign T_629 = T_622 ? 2'h3 : T_628;
  assign T_630 = T_613 ? T_621 : T_629;
  assign T_631 = {T_613,T_630};
  assign T_632 = T_587 ? T_609 : T_631;
  assign T_633 = {T_587,T_632};
  assign T_634 = T_533 ? T_583 : T_633;
  assign T_635 = {T_533,T_634};
  assign T_636 = T_423 ? T_529 : T_635;
  assign T_637 = {T_423,T_636};
  assign T_638 = ~ T_637;
  assign GEN_49 = {{63'd0}, T_413};
  assign T_639 = GEN_49 << T_638;
  assign T_640 = T_639[50:0];
  assign T_642 = {T_640,1'h0};
  assign GEN_50 = {{6'd0}, T_638};
  assign T_648 = GEN_50 ^ 12'hfff;
  assign T_649 = T_415 ? T_648 : {{1'd0}, T_412};
  assign T_653 = T_415 ? 2'h2 : 2'h1;
  assign GEN_51 = {{9'd0}, T_653};
  assign T_654 = 11'h400 | GEN_51;
  assign GEN_52 = {{1'd0}, T_654};
  assign T_655 = T_649 + GEN_52;
  assign T_656 = T_655[11:0];
  assign T_657 = T_656[11:10];
  assign T_659 = T_657 == 2'h3;
  assign T_661 = T_417 == 1'h0;
  assign T_662 = T_659 & T_661;
  assign T_666 = T_418 ? 3'h7 : 3'h0;
  assign GEN_53 = {{9'd0}, T_666};
  assign T_667 = GEN_53 << 9;
  assign T_668 = ~ T_667;
  assign T_669 = T_656 & T_668;
  assign GEN_54 = {{9'd0}, T_662};
  assign T_670 = GEN_54 << 9;
  assign GEN_55 = {{2'd0}, T_670};
  assign T_671 = T_669 | GEN_55;
  assign T_672 = T_415 ? T_642 : T_413;
  assign T_673 = {T_411,T_671};
  assign T_674 = {T_673,T_672};
  assign GEN_22 = T_410 ? T_674 : {{32'd0}, T_408};
  assign T_675 = $signed(in_bits_in1);
  assign T_676 = GEN_23;
  assign T_677 = in_bits_in1[31:0];
  assign T_678 = in_bits_typ[1];
  assign T_680 = T_678 == 1'h0;
  assign T_681 = in_bits_typ[0];
  assign T_682 = {1'b0,$signed(T_677)};
  assign T_683 = $signed(T_677);
  assign T_684 = T_681 ? $signed(T_682) : $signed({{1{T_683[31]}},T_683});
  assign GEN_23 = T_680 ? $signed({{32{T_684[32]}},T_684}) : $signed(T_675);
  assign intValue = $unsigned(T_676);
  assign T_687 = in_bits_cmd & 5'h4;
  assign T_688 = 5'h0 == T_687;
  assign INToRecFN_2_clk = clk;
  assign INToRecFN_2_reset = reset;
  assign INToRecFN_2_io_signedIn = T_690;
  assign INToRecFN_2_io_in = intValue[63:0];
  assign INToRecFN_2_io_roundingMode = in_bits_rm[1:0];
  assign T_690 = ~ T_681;
  assign T_692 = {32'hffffffff,INToRecFN_2_io_out};
  assign INToRecFN_1_1_clk = clk;
  assign INToRecFN_1_1_reset = reset;
  assign INToRecFN_1_1_io_signedIn = T_690;
  assign INToRecFN_1_1_io_in = intValue[63:0];
  assign INToRecFN_1_1_io_roundingMode = in_bits_rm[1:0];
  assign T_698 = {1'h0,INToRecFN_1_1_io_out};
  assign GEN_24 = T_410 ? T_698 : {{1'd0}, T_692};
  assign GEN_25 = T_410 ? INToRecFN_1_1_io_exceptionFlags : INToRecFN_2_io_exceptionFlags;
  assign GEN_31 = T_688 ? GEN_24 : {{1'd0}, GEN_22};
  assign GEN_32 = T_688 ? GEN_25 : 5'h0;
  assign GEN_38 = in_valid ? mux_data : T_702_data;
  assign GEN_39 = in_valid ? mux_exc : T_702_exc;
  assign T_713_valid = T_701;
  assign T_713_bits_data = T_702_data;
  assign T_713_bits_exc = T_702_exc;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  T_132 = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  T_133_cmd = GEN_27[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  T_133_ldst = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  T_133_wen = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  T_133_ren1 = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  T_133_ren2 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  T_133_ren3 = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  T_133_swap12 = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  T_133_swap23 = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  T_133_single = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  T_133_fromint = GEN_56[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  T_133_toint = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  T_133_fastpipe = GEN_58[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  T_133_fma = GEN_59[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {1{$random}};
  T_133_div = GEN_60[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_61 = {1{$random}};
  T_133_sqrt = GEN_61[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_62 = {1{$random}};
  T_133_round = GEN_62[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_63 = {1{$random}};
  T_133_wflags = GEN_63[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_64 = {1{$random}};
  T_133_rm = GEN_64[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_65 = {1{$random}};
  T_133_typ = GEN_65[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_66 = {3{$random}};
  T_133_in1 = GEN_66[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_67 = {3{$random}};
  T_133_in2 = GEN_67[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_68 = {3{$random}};
  T_133_in3 = GEN_68[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_69 = {1{$random}};
  T_701 = GEN_69[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_70 = {3{$random}};
  T_702_data = GEN_70[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_71 = {1{$random}};
  T_702_exc = GEN_71[4:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_132 <= 1'h0;
    end else begin
      T_132 <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_cmd <= io_in_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_ldst <= io_in_bits_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_wen <= io_in_bits_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_ren1 <= io_in_bits_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_ren2 <= io_in_bits_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_ren3 <= io_in_bits_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_swap12 <= io_in_bits_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_swap23 <= io_in_bits_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_single <= io_in_bits_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_fromint <= io_in_bits_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_toint <= io_in_bits_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_fastpipe <= io_in_bits_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_fma <= io_in_bits_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_div <= io_in_bits_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_sqrt <= io_in_bits_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_round <= io_in_bits_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_wflags <= io_in_bits_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_rm <= io_in_bits_rm;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_typ <= io_in_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_in1 <= io_in_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_in2 <= io_in_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_133_in3 <= io_in_bits_in3;
      end
    end
    if(reset) begin
      T_701 <= 1'h0;
    end else begin
      T_701 <= in_valid;
    end
    if(1'h0) begin
    end else begin
      if(in_valid) begin
        T_702_data <= mux_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(in_valid) begin
        T_702_exc <= mux_exc;
      end
    end
  end
endmodule
module RoundRawFNToRecFN(
  input   clk,
  input   reset,
  input   io_invalidExc,
  input   io_infiniteExc,
  input   io_in_sign,
  input   io_in_isNaN,
  input   io_in_isInf,
  input   io_in_isZero,
  input  [9:0] io_in_sExp,
  input  [26:0] io_in_sig,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  T_19;
  wire  T_21;
  wire  T_22;
  wire  roundMagUp;
  wire  doShiftSigDown1;
  wire  isNegExp;
  wire [24:0] T_27;
  wire [8:0] T_28;
  wire [8:0] T_29;
  wire  T_30;
  wire [7:0] T_31;
  wire  T_32;
  wire [6:0] T_33;
  wire  T_34;
  wire [5:0] T_35;
  wire [64:0] T_38;
  wire [21:0] T_39;
  wire [15:0] T_40;
  wire [7:0] T_45;
  wire [15:0] T_46;
  wire [7:0] T_47;
  wire [15:0] GEN_0;
  wire [15:0] T_48;
  wire [15:0] T_50;
  wire [15:0] T_51;
  wire [11:0] T_55;
  wire [15:0] GEN_1;
  wire [15:0] T_56;
  wire [11:0] T_57;
  wire [15:0] GEN_2;
  wire [15:0] T_58;
  wire [15:0] T_60;
  wire [15:0] T_61;
  wire [13:0] T_65;
  wire [15:0] GEN_3;
  wire [15:0] T_66;
  wire [13:0] T_67;
  wire [15:0] GEN_4;
  wire [15:0] T_68;
  wire [15:0] T_70;
  wire [15:0] T_71;
  wire [14:0] T_75;
  wire [15:0] GEN_5;
  wire [15:0] T_76;
  wire [14:0] T_77;
  wire [15:0] GEN_6;
  wire [15:0] T_78;
  wire [15:0] T_80;
  wire [15:0] T_81;
  wire [5:0] T_82;
  wire [3:0] T_83;
  wire [1:0] T_84;
  wire  T_85;
  wire  T_86;
  wire [1:0] T_87;
  wire [1:0] T_88;
  wire  T_89;
  wire  T_90;
  wire [1:0] T_91;
  wire [3:0] T_92;
  wire [1:0] T_93;
  wire  T_94;
  wire  T_95;
  wire [1:0] T_96;
  wire [5:0] T_97;
  wire [21:0] T_98;
  wire [21:0] T_99;
  wire [21:0] T_100;
  wire [21:0] T_101;
  wire [24:0] T_103;
  wire [2:0] T_108;
  wire [1:0] T_109;
  wire  T_110;
  wire  T_111;
  wire [1:0] T_112;
  wire  T_113;
  wire [2:0] T_114;
  wire [2:0] T_116;
  wire [24:0] T_117;
  wire [24:0] T_119;
  wire [24:0] T_120;
  wire [24:0] GEN_7;
  wire [24:0] T_121;
  wire [26:0] roundMask;
  wire [27:0] T_123;
  wire [26:0] shiftedRoundMask;
  wire [26:0] T_124;
  wire [26:0] roundPosMask;
  wire [26:0] T_125;
  wire  roundPosBit;
  wire [26:0] T_127;
  wire  anyRoundExtra;
  wire  common_inexact;
  wire  T_129;
  wire  T_130;
  wire  T_131;
  wire [26:0] T_132;
  wire [24:0] T_133;
  wire [25:0] T_135;
  wire  T_138;
  wire  T_139;
  wire [25:0] T_140;
  wire [25:0] T_142;
  wire [25:0] T_143;
  wire [25:0] T_144;
  wire [26:0] T_145;
  wire [26:0] T_146;
  wire [24:0] T_147;
  wire [25:0] roundedSig;
  wire [1:0] T_148;
  wire [2:0] T_149;
  wire [9:0] GEN_8;
  wire [10:0] sRoundedExp;
  wire [8:0] common_expOut;
  wire [22:0] T_150;
  wire [22:0] T_151;
  wire [22:0] common_fractOut;
  wire [3:0] T_152;
  wire  common_overflow;
  wire  common_totalUnderflow;
  wire [8:0] T_157;
  wire [9:0] GEN_9;
  wire  T_158;
  wire  common_underflow;
  wire  isNaNOut;
  wire  notNaN_isSpecialInfOut;
  wire  T_160;
  wire  T_162;
  wire  T_163;
  wire  T_165;
  wire  commonCase;
  wire  overflow;
  wire  underflow;
  wire  T_166;
  wire  inexact;
  wire  overflow_roundMagUp;
  wire  T_167;
  wire  pegMinNonzeroMagOut;
  wire  T_168;
  wire  T_170;
  wire  pegMaxFiniteMagOut;
  wire  T_171;
  wire  notNaN_isInfOut;
  wire  signOut;
  wire  T_173;
  wire [8:0] T_176;
  wire [8:0] T_177;
  wire [8:0] T_178;
  wire [8:0] T_182;
  wire [8:0] T_183;
  wire [8:0] T_184;
  wire [8:0] T_187;
  wire [8:0] T_188;
  wire [8:0] T_189;
  wire [8:0] T_192;
  wire [8:0] T_193;
  wire [8:0] T_194;
  wire [8:0] T_197;
  wire [8:0] T_198;
  wire [8:0] T_201;
  wire [8:0] T_202;
  wire [8:0] T_205;
  wire [8:0] T_206;
  wire [8:0] T_209;
  wire [8:0] expOut;
  wire  T_210;
  wire [22:0] T_214;
  wire [22:0] T_215;
  wire [22:0] T_219;
  wire [22:0] fractOut;
  wire [9:0] T_220;
  wire [32:0] T_221;
  wire [1:0] T_222;
  wire [1:0] T_223;
  wire [2:0] T_224;
  wire [4:0] T_225;
  assign io_out = T_221;
  assign io_exceptionFlags = T_225;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign T_19 = roundingMode_min & io_in_sign;
  assign T_21 = io_in_sign == 1'h0;
  assign T_22 = roundingMode_max & T_21;
  assign roundMagUp = T_19 | T_22;
  assign doShiftSigDown1 = io_in_sig[26];
  assign isNegExp = $signed(io_in_sExp) < $signed(10'sh0);
  assign T_27 = isNegExp ? 25'h1ffffff : 25'h0;
  assign T_28 = io_in_sExp[8:0];
  assign T_29 = ~ T_28;
  assign T_30 = T_29[8];
  assign T_31 = T_29[7:0];
  assign T_32 = T_31[7];
  assign T_33 = T_31[6:0];
  assign T_34 = T_33[6];
  assign T_35 = T_33[5:0];
  assign T_38 = $signed(65'sh10000000000000000) >>> T_35;
  assign T_39 = T_38[63:42];
  assign T_40 = T_39[15:0];
  assign T_45 = T_40[15:8];
  assign T_46 = {{8'd0}, T_45};
  assign T_47 = T_40[7:0];
  assign GEN_0 = {{8'd0}, T_47};
  assign T_48 = GEN_0 << 8;
  assign T_50 = T_48 & 16'hff00;
  assign T_51 = T_46 | T_50;
  assign T_55 = T_51[15:4];
  assign GEN_1 = {{4'd0}, T_55};
  assign T_56 = GEN_1 & 16'hf0f;
  assign T_57 = T_51[11:0];
  assign GEN_2 = {{4'd0}, T_57};
  assign T_58 = GEN_2 << 4;
  assign T_60 = T_58 & 16'hf0f0;
  assign T_61 = T_56 | T_60;
  assign T_65 = T_61[15:2];
  assign GEN_3 = {{2'd0}, T_65};
  assign T_66 = GEN_3 & 16'h3333;
  assign T_67 = T_61[13:0];
  assign GEN_4 = {{2'd0}, T_67};
  assign T_68 = GEN_4 << 2;
  assign T_70 = T_68 & 16'hcccc;
  assign T_71 = T_66 | T_70;
  assign T_75 = T_71[15:1];
  assign GEN_5 = {{1'd0}, T_75};
  assign T_76 = GEN_5 & 16'h5555;
  assign T_77 = T_71[14:0];
  assign GEN_6 = {{1'd0}, T_77};
  assign T_78 = GEN_6 << 1;
  assign T_80 = T_78 & 16'haaaa;
  assign T_81 = T_76 | T_80;
  assign T_82 = T_39[21:16];
  assign T_83 = T_82[3:0];
  assign T_84 = T_83[1:0];
  assign T_85 = T_84[0];
  assign T_86 = T_84[1];
  assign T_87 = {T_85,T_86};
  assign T_88 = T_83[3:2];
  assign T_89 = T_88[0];
  assign T_90 = T_88[1];
  assign T_91 = {T_89,T_90};
  assign T_92 = {T_87,T_91};
  assign T_93 = T_82[5:4];
  assign T_94 = T_93[0];
  assign T_95 = T_93[1];
  assign T_96 = {T_94,T_95};
  assign T_97 = {T_92,T_96};
  assign T_98 = {T_81,T_97};
  assign T_99 = ~ T_98;
  assign T_100 = T_34 ? 22'h0 : T_99;
  assign T_101 = ~ T_100;
  assign T_103 = {T_101,3'h7};
  assign T_108 = T_38[2:0];
  assign T_109 = T_108[1:0];
  assign T_110 = T_109[0];
  assign T_111 = T_109[1];
  assign T_112 = {T_110,T_111};
  assign T_113 = T_108[2];
  assign T_114 = {T_112,T_113};
  assign T_116 = T_34 ? T_114 : 3'h0;
  assign T_117 = T_32 ? T_103 : {{22'd0}, T_116};
  assign T_119 = T_30 ? T_117 : 25'h0;
  assign T_120 = T_27 | T_119;
  assign GEN_7 = {{24'd0}, doShiftSigDown1};
  assign T_121 = T_120 | GEN_7;
  assign roundMask = {T_121,2'h3};
  assign T_123 = {isNegExp,roundMask};
  assign shiftedRoundMask = T_123[27:1];
  assign T_124 = ~ shiftedRoundMask;
  assign roundPosMask = T_124 & roundMask;
  assign T_125 = io_in_sig & roundPosMask;
  assign roundPosBit = T_125 != 27'h0;
  assign T_127 = io_in_sig & shiftedRoundMask;
  assign anyRoundExtra = T_127 != 27'h0;
  assign common_inexact = roundPosBit | anyRoundExtra;
  assign T_129 = roundingMode_nearest_even & roundPosBit;
  assign T_130 = roundMagUp & common_inexact;
  assign T_131 = T_129 | T_130;
  assign T_132 = io_in_sig | roundMask;
  assign T_133 = T_132[26:2];
  assign T_135 = T_133 + 25'h1;
  assign T_138 = anyRoundExtra == 1'h0;
  assign T_139 = T_129 & T_138;
  assign T_140 = roundMask[26:1];
  assign T_142 = T_139 ? T_140 : 26'h0;
  assign T_143 = ~ T_142;
  assign T_144 = T_135 & T_143;
  assign T_145 = ~ roundMask;
  assign T_146 = io_in_sig & T_145;
  assign T_147 = T_146[26:2];
  assign roundedSig = T_131 ? T_144 : {{1'd0}, T_147};
  assign T_148 = roundedSig[25:24];
  assign T_149 = {1'b0,$signed(T_148)};
  assign GEN_8 = {{7{T_149[2]}},T_149};
  assign sRoundedExp = $signed(io_in_sExp) + $signed(GEN_8);
  assign common_expOut = sRoundedExp[8:0];
  assign T_150 = roundedSig[23:1];
  assign T_151 = roundedSig[22:0];
  assign common_fractOut = doShiftSigDown1 ? T_150 : T_151;
  assign T_152 = sRoundedExp[10:7];
  assign common_overflow = $signed(T_152) >= $signed(4'sh3);
  assign common_totalUnderflow = $signed(sRoundedExp) < $signed(11'sh6b);
  assign T_157 = doShiftSigDown1 ? $signed(9'sh81) : $signed(9'sh82);
  assign GEN_9 = {{1{T_157[8]}},T_157};
  assign T_158 = $signed(io_in_sExp) < $signed(GEN_9);
  assign common_underflow = common_inexact & T_158;
  assign isNaNOut = io_invalidExc | io_in_isNaN;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T_160 = isNaNOut == 1'h0;
  assign T_162 = notNaN_isSpecialInfOut == 1'h0;
  assign T_163 = T_160 & T_162;
  assign T_165 = io_in_isZero == 1'h0;
  assign commonCase = T_163 & T_165;
  assign overflow = commonCase & common_overflow;
  assign underflow = commonCase & common_underflow;
  assign T_166 = commonCase & common_inexact;
  assign inexact = overflow | T_166;
  assign overflow_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign T_167 = commonCase & common_totalUnderflow;
  assign pegMinNonzeroMagOut = T_167 & roundMagUp;
  assign T_168 = commonCase & overflow;
  assign T_170 = overflow_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = T_168 & T_170;
  assign T_171 = overflow & overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T_171;
  assign signOut = isNaNOut ? 1'h0 : io_in_sign;
  assign T_173 = io_in_isZero | common_totalUnderflow;
  assign T_176 = T_173 ? 9'h1c0 : 9'h0;
  assign T_177 = ~ T_176;
  assign T_178 = common_expOut & T_177;
  assign T_182 = pegMinNonzeroMagOut ? 9'h194 : 9'h0;
  assign T_183 = ~ T_182;
  assign T_184 = T_178 & T_183;
  assign T_187 = pegMaxFiniteMagOut ? 9'h80 : 9'h0;
  assign T_188 = ~ T_187;
  assign T_189 = T_184 & T_188;
  assign T_192 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T_193 = ~ T_192;
  assign T_194 = T_189 & T_193;
  assign T_197 = pegMinNonzeroMagOut ? 9'h6b : 9'h0;
  assign T_198 = T_194 | T_197;
  assign T_201 = pegMaxFiniteMagOut ? 9'h17f : 9'h0;
  assign T_202 = T_198 | T_201;
  assign T_205 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign T_206 = T_202 | T_205;
  assign T_209 = isNaNOut ? 9'h1c0 : 9'h0;
  assign expOut = T_206 | T_209;
  assign T_210 = common_totalUnderflow | isNaNOut;
  assign T_214 = isNaNOut ? 23'h400000 : 23'h0;
  assign T_215 = T_210 ? T_214 : common_fractOut;
  assign T_219 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0;
  assign fractOut = T_215 | T_219;
  assign T_220 = {signOut,expOut};
  assign T_221 = {T_220,fractOut};
  assign T_222 = {underflow,inexact};
  assign T_223 = {io_invalidExc,io_infiniteExc};
  assign T_224 = {T_223,overflow};
  assign T_225 = {T_224,T_222};
endmodule
module RecFNToRecFN(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_4;
  wire [2:0] T_5;
  wire  T_7;
  wire [1:0] T_8;
  wire  T_10;
  wire  T_18_sign;
  wire  T_18_isNaN;
  wire  T_18_isInf;
  wire  T_18_isZero;
  wire [12:0] T_18_sExp;
  wire [55:0] T_18_sig;
  wire  T_25;
  wire  T_26;
  wire  T_27;
  wire  T_30;
  wire  T_31;
  wire [12:0] T_32;
  wire  T_35;
  wire [51:0] T_36;
  wire [53:0] T_38;
  wire [1:0] T_39;
  wire [55:0] T_40;
  wire [13:0] T_42;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [9:0] outRawFloat_sExp;
  wire [26:0] outRawFloat_sig;
  wire  T_57;
  wire [3:0] T_58;
  wire  T_60;
  wire [8:0] T_68;
  wire [8:0] T_69;
  wire [9:0] T_70;
  wire [9:0] T_71;
  wire [25:0] T_72;
  wire [29:0] T_73;
  wire  T_75;
  wire [26:0] T_76;
  wire  T_77;
  wire  T_79;
  wire  invalidExc;
  wire  RoundRawFNToRecFN_1_clk;
  wire  RoundRawFNToRecFN_1_reset;
  wire  RoundRawFNToRecFN_1_io_invalidExc;
  wire  RoundRawFNToRecFN_1_io_infiniteExc;
  wire  RoundRawFNToRecFN_1_io_in_sign;
  wire  RoundRawFNToRecFN_1_io_in_isNaN;
  wire  RoundRawFNToRecFN_1_io_in_isInf;
  wire  RoundRawFNToRecFN_1_io_in_isZero;
  wire [9:0] RoundRawFNToRecFN_1_io_in_sExp;
  wire [26:0] RoundRawFNToRecFN_1_io_in_sig;
  wire [1:0] RoundRawFNToRecFN_1_io_roundingMode;
  wire [32:0] RoundRawFNToRecFN_1_io_out;
  wire [4:0] RoundRawFNToRecFN_1_io_exceptionFlags;
  RoundRawFNToRecFN RoundRawFNToRecFN_1 (
    .clk(RoundRawFNToRecFN_1_clk),
    .reset(RoundRawFNToRecFN_1_reset),
    .io_invalidExc(RoundRawFNToRecFN_1_io_invalidExc),
    .io_infiniteExc(RoundRawFNToRecFN_1_io_infiniteExc),
    .io_in_sign(RoundRawFNToRecFN_1_io_in_sign),
    .io_in_isNaN(RoundRawFNToRecFN_1_io_in_isNaN),
    .io_in_isInf(RoundRawFNToRecFN_1_io_in_isInf),
    .io_in_isZero(RoundRawFNToRecFN_1_io_in_isZero),
    .io_in_sExp(RoundRawFNToRecFN_1_io_in_sExp),
    .io_in_sig(RoundRawFNToRecFN_1_io_in_sig),
    .io_roundingMode(RoundRawFNToRecFN_1_io_roundingMode),
    .io_out(RoundRawFNToRecFN_1_io_out),
    .io_exceptionFlags(RoundRawFNToRecFN_1_io_exceptionFlags)
  );
  assign io_out = RoundRawFNToRecFN_1_io_out;
  assign io_exceptionFlags = RoundRawFNToRecFN_1_io_exceptionFlags;
  assign T_4 = io_in[63:52];
  assign T_5 = T_4[11:9];
  assign T_7 = T_5 == 3'h0;
  assign T_8 = T_4[11:10];
  assign T_10 = T_8 == 2'h3;
  assign T_18_sign = T_25;
  assign T_18_isNaN = T_27;
  assign T_18_isInf = T_31;
  assign T_18_isZero = T_7;
  assign T_18_sExp = T_32;
  assign T_18_sig = T_40;
  assign T_25 = io_in[64];
  assign T_26 = T_4[9];
  assign T_27 = T_10 & T_26;
  assign T_30 = T_26 == 1'h0;
  assign T_31 = T_10 & T_30;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_35 = T_7 == 1'h0;
  assign T_36 = io_in[51:0];
  assign T_38 = {T_36,2'h0};
  assign T_39 = {1'h0,T_35};
  assign T_40 = {T_39,T_38};
  assign T_42 = $signed(T_18_sExp) + $signed(13'sh1900);
  assign outRawFloat_sign = T_18_sign;
  assign outRawFloat_isNaN = T_18_isNaN;
  assign outRawFloat_isInf = T_18_isInf;
  assign outRawFloat_isZero = T_18_isZero;
  assign outRawFloat_sExp = T_71;
  assign outRawFloat_sig = T_76;
  assign T_57 = $signed(T_42) < $signed(14'sh0);
  assign T_58 = T_42[12:9];
  assign T_60 = T_58 != 4'h0;
  assign T_68 = T_42[8:0];
  assign T_69 = T_60 ? 9'h1fc : T_68;
  assign T_70 = {T_57,T_69};
  assign T_71 = $signed(T_70);
  assign T_72 = T_18_sig[55:30];
  assign T_73 = T_18_sig[29:0];
  assign T_75 = T_73 != 30'h0;
  assign T_76 = {T_72,T_75};
  assign T_77 = outRawFloat_sig[24];
  assign T_79 = T_77 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_79;
  assign RoundRawFNToRecFN_1_clk = clk;
  assign RoundRawFNToRecFN_1_reset = reset;
  assign RoundRawFNToRecFN_1_io_invalidExc = invalidExc;
  assign RoundRawFNToRecFN_1_io_infiniteExc = 1'h0;
  assign RoundRawFNToRecFN_1_io_in_sign = outRawFloat_sign;
  assign RoundRawFNToRecFN_1_io_in_isNaN = outRawFloat_isNaN;
  assign RoundRawFNToRecFN_1_io_in_isInf = outRawFloat_isInf;
  assign RoundRawFNToRecFN_1_io_in_isZero = outRawFloat_isZero;
  assign RoundRawFNToRecFN_1_io_in_sExp = outRawFloat_sExp;
  assign RoundRawFNToRecFN_1_io_in_sig = outRawFloat_sig;
  assign RoundRawFNToRecFN_1_io_roundingMode = io_roundingMode;
endmodule
module RecFNToRecFN_1(
  input   clk,
  input   reset,
  input  [32:0] io_in,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [8:0] T_4;
  wire [2:0] T_5;
  wire  T_7;
  wire [1:0] T_8;
  wire  T_10;
  wire  T_18_sign;
  wire  T_18_isNaN;
  wire  T_18_isInf;
  wire  T_18_isZero;
  wire [9:0] T_18_sExp;
  wire [26:0] T_18_sig;
  wire  T_25;
  wire  T_26;
  wire  T_27;
  wire  T_30;
  wire  T_31;
  wire [9:0] T_32;
  wire  T_35;
  wire [22:0] T_36;
  wire [24:0] T_38;
  wire [1:0] T_39;
  wire [26:0] T_40;
  wire [11:0] GEN_0;
  wire [12:0] T_42;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [12:0] outRawFloat_sExp;
  wire [55:0] outRawFloat_sig;
  wire [55:0] GEN_1;
  wire [55:0] T_56;
  wire  T_57;
  wire  T_59;
  wire  invalidExc;
  wire  T_61;
  wire  T_62;
  wire [11:0] T_63;
  wire [11:0] T_66;
  wire [11:0] T_67;
  wire [11:0] T_68;
  wire  T_69;
  wire [11:0] T_72;
  wire [11:0] T_73;
  wire [11:0] T_74;
  wire [11:0] T_77;
  wire [11:0] T_78;
  wire [11:0] T_81;
  wire [11:0] T_82;
  wire [51:0] T_85;
  wire [51:0] T_86;
  wire [12:0] T_87;
  wire [64:0] T_88;
  wire [4:0] T_90;
  assign io_out = T_88;
  assign io_exceptionFlags = T_90;
  assign T_4 = io_in[31:23];
  assign T_5 = T_4[8:6];
  assign T_7 = T_5 == 3'h0;
  assign T_8 = T_4[8:7];
  assign T_10 = T_8 == 2'h3;
  assign T_18_sign = T_25;
  assign T_18_isNaN = T_27;
  assign T_18_isInf = T_31;
  assign T_18_isZero = T_7;
  assign T_18_sExp = T_32;
  assign T_18_sig = T_40;
  assign T_25 = io_in[32];
  assign T_26 = T_4[6];
  assign T_27 = T_10 & T_26;
  assign T_30 = T_26 == 1'h0;
  assign T_31 = T_10 & T_30;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_35 = T_7 == 1'h0;
  assign T_36 = io_in[22:0];
  assign T_38 = {T_36,2'h0};
  assign T_39 = {1'h0,T_35};
  assign T_40 = {T_39,T_38};
  assign GEN_0 = {{2{T_18_sExp[9]}},T_18_sExp};
  assign T_42 = $signed(GEN_0) + $signed(12'sh700);
  assign outRawFloat_sign = T_18_sign;
  assign outRawFloat_isNaN = T_18_isNaN;
  assign outRawFloat_isInf = T_18_isInf;
  assign outRawFloat_isZero = T_18_isZero;
  assign outRawFloat_sExp = T_42;
  assign outRawFloat_sig = T_56;
  assign GEN_1 = {{29'd0}, T_18_sig};
  assign T_56 = GEN_1 << 29;
  assign T_57 = outRawFloat_sig[53];
  assign T_59 = T_57 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_59;
  assign T_61 = outRawFloat_isNaN == 1'h0;
  assign T_62 = outRawFloat_sign & T_61;
  assign T_63 = outRawFloat_sExp[11:0];
  assign T_66 = outRawFloat_isZero ? 12'hc00 : 12'h0;
  assign T_67 = ~ T_66;
  assign T_68 = T_63 & T_67;
  assign T_69 = outRawFloat_isZero | outRawFloat_isInf;
  assign T_72 = T_69 ? 12'h200 : 12'h0;
  assign T_73 = ~ T_72;
  assign T_74 = T_68 & T_73;
  assign T_77 = outRawFloat_isInf ? 12'hc00 : 12'h0;
  assign T_78 = T_74 | T_77;
  assign T_81 = outRawFloat_isNaN ? 12'he00 : 12'h0;
  assign T_82 = T_78 | T_81;
  assign T_85 = outRawFloat_sig[53:2];
  assign T_86 = outRawFloat_isNaN ? 52'h8000000000000 : T_85;
  assign T_87 = {T_62,T_82};
  assign T_88 = {T_87,T_86};
  assign T_90 = {invalidExc,4'h0};
endmodule
module FPToFP(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  input   io_lt
);
  reg  T_133;
  reg [31:0] GEN_25;
  reg [4:0] T_134_cmd;
  reg [31:0] GEN_26;
  reg  T_134_ldst;
  reg [31:0] GEN_27;
  reg  T_134_wen;
  reg [31:0] GEN_28;
  reg  T_134_ren1;
  reg [31:0] GEN_31;
  reg  T_134_ren2;
  reg [31:0] GEN_32;
  reg  T_134_ren3;
  reg [31:0] GEN_33;
  reg  T_134_swap12;
  reg [31:0] GEN_34;
  reg  T_134_swap23;
  reg [31:0] GEN_37;
  reg  T_134_single;
  reg [31:0] GEN_38;
  reg  T_134_fromint;
  reg [31:0] GEN_39;
  reg  T_134_toint;
  reg [31:0] GEN_40;
  reg  T_134_fastpipe;
  reg [31:0] GEN_43;
  reg  T_134_fma;
  reg [31:0] GEN_44;
  reg  T_134_div;
  reg [31:0] GEN_45;
  reg  T_134_sqrt;
  reg [31:0] GEN_46;
  reg  T_134_round;
  reg [31:0] GEN_50;
  reg  T_134_wflags;
  reg [31:0] GEN_51;
  reg [2:0] T_134_rm;
  reg [31:0] GEN_52;
  reg [1:0] T_134_typ;
  reg [31:0] GEN_53;
  reg [64:0] T_134_in1;
  reg [95:0] GEN_54;
  reg [64:0] T_134_in2;
  reg [95:0] GEN_55;
  reg [64:0] T_134_in3;
  reg [95:0] GEN_56;
  wire [4:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire [64:0] GEN_19;
  wire [64:0] GEN_20;
  wire [64:0] GEN_21;
  wire  in_valid;
  wire [4:0] in_bits_cmd;
  wire  in_bits_ldst;
  wire  in_bits_wen;
  wire  in_bits_ren1;
  wire  in_bits_ren2;
  wire  in_bits_ren3;
  wire  in_bits_swap12;
  wire  in_bits_swap23;
  wire  in_bits_single;
  wire  in_bits_fromint;
  wire  in_bits_toint;
  wire  in_bits_fastpipe;
  wire  in_bits_fma;
  wire  in_bits_div;
  wire  in_bits_sqrt;
  wire  in_bits_round;
  wire  in_bits_wflags;
  wire [2:0] in_bits_rm;
  wire [1:0] in_bits_typ;
  wire [64:0] in_bits_in1;
  wire [64:0] in_bits_in2;
  wire [64:0] in_bits_in3;
  wire  T_252;
  wire [64:0] T_253;
  wire  T_254;
  wire [64:0] T_255;
  wire [64:0] T_256;
  wire [64:0] signNum;
  wire  T_257;
  wire [31:0] T_258;
  wire [32:0] fsgnj_s;
  wire [31:0] T_259;
  wire [64:0] T_260;
  wire  T_261;
  wire [63:0] T_262;
  wire [64:0] T_263;
  wire [64:0] fsgnj;
  wire [64:0] mux_data;
  wire [4:0] mux_exc;
  wire [4:0] T_272;
  wire  T_273;
  wire [2:0] T_274;
  wire [2:0] T_275;
  wire  T_277;
  wire [2:0] T_278;
  wire [2:0] T_279;
  wire  T_281;
  wire  T_286;
  wire  T_288;
  wire  T_289;
  wire  T_294;
  wire  T_296;
  wire  T_297;
  wire  T_299;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_304;
  wire [2:0] T_305;
  wire [2:0] T_306;
  wire  T_308;
  wire [2:0] T_309;
  wire [2:0] T_310;
  wire  T_312;
  wire  T_317;
  wire  T_319;
  wire  T_320;
  wire  T_325;
  wire  T_327;
  wire  T_328;
  wire  T_332;
  wire  T_333;
  wire  T_334;
  wire  T_335;
  wire  T_336;
  wire  T_337;
  wire [4:0] GEN_49;
  wire [4:0] T_338;
  wire  T_340;
  wire [64:0] GEN_22;
  wire [4:0] GEN_23;
  wire [64:0] GEN_24;
  wire [4:0] T_343;
  wire  T_344;
  wire  RecFNToRecFN_2_clk;
  wire  RecFNToRecFN_2_reset;
  wire [64:0] RecFNToRecFN_2_io_in;
  wire [1:0] RecFNToRecFN_2_io_roundingMode;
  wire [32:0] RecFNToRecFN_2_io_out;
  wire [4:0] RecFNToRecFN_2_io_exceptionFlags;
  wire [64:0] T_346;
  wire [64:0] GEN_29;
  wire [4:0] GEN_30;
  wire  T_348;
  wire  RecFNToRecFN_1_1_clk;
  wire  RecFNToRecFN_1_1_reset;
  wire [32:0] RecFNToRecFN_1_1_io_in;
  wire [1:0] RecFNToRecFN_1_1_io_roundingMode;
  wire [64:0] RecFNToRecFN_1_1_io_out;
  wire [4:0] RecFNToRecFN_1_1_io_exceptionFlags;
  wire [64:0] GEN_35;
  wire [4:0] GEN_36;
  wire [64:0] GEN_41;
  wire [4:0] GEN_42;
  reg  T_351;
  reg [31:0] GEN_57;
  reg [64:0] T_352_data;
  reg [95:0] GEN_58;
  reg [4:0] T_352_exc;
  reg [31:0] GEN_59;
  wire [64:0] GEN_47;
  wire [4:0] GEN_48;
  wire  T_363_valid;
  wire [64:0] T_363_bits_data;
  wire [4:0] T_363_bits_exc;
  RecFNToRecFN RecFNToRecFN_2 (
    .clk(RecFNToRecFN_2_clk),
    .reset(RecFNToRecFN_2_reset),
    .io_in(RecFNToRecFN_2_io_in),
    .io_roundingMode(RecFNToRecFN_2_io_roundingMode),
    .io_out(RecFNToRecFN_2_io_out),
    .io_exceptionFlags(RecFNToRecFN_2_io_exceptionFlags)
  );
  RecFNToRecFN_1 RecFNToRecFN_1_1 (
    .clk(RecFNToRecFN_1_1_clk),
    .reset(RecFNToRecFN_1_1_reset),
    .io_in(RecFNToRecFN_1_1_io_in),
    .io_roundingMode(RecFNToRecFN_1_1_io_roundingMode),
    .io_out(RecFNToRecFN_1_1_io_out),
    .io_exceptionFlags(RecFNToRecFN_1_1_io_exceptionFlags)
  );
  assign io_out_valid = T_363_valid;
  assign io_out_bits_data = T_363_bits_data;
  assign io_out_bits_exc = T_363_bits_exc;
  assign GEN_0 = io_in_valid ? io_in_bits_cmd : T_134_cmd;
  assign GEN_1 = io_in_valid ? io_in_bits_ldst : T_134_ldst;
  assign GEN_2 = io_in_valid ? io_in_bits_wen : T_134_wen;
  assign GEN_3 = io_in_valid ? io_in_bits_ren1 : T_134_ren1;
  assign GEN_4 = io_in_valid ? io_in_bits_ren2 : T_134_ren2;
  assign GEN_5 = io_in_valid ? io_in_bits_ren3 : T_134_ren3;
  assign GEN_6 = io_in_valid ? io_in_bits_swap12 : T_134_swap12;
  assign GEN_7 = io_in_valid ? io_in_bits_swap23 : T_134_swap23;
  assign GEN_8 = io_in_valid ? io_in_bits_single : T_134_single;
  assign GEN_9 = io_in_valid ? io_in_bits_fromint : T_134_fromint;
  assign GEN_10 = io_in_valid ? io_in_bits_toint : T_134_toint;
  assign GEN_11 = io_in_valid ? io_in_bits_fastpipe : T_134_fastpipe;
  assign GEN_12 = io_in_valid ? io_in_bits_fma : T_134_fma;
  assign GEN_13 = io_in_valid ? io_in_bits_div : T_134_div;
  assign GEN_14 = io_in_valid ? io_in_bits_sqrt : T_134_sqrt;
  assign GEN_15 = io_in_valid ? io_in_bits_round : T_134_round;
  assign GEN_16 = io_in_valid ? io_in_bits_wflags : T_134_wflags;
  assign GEN_17 = io_in_valid ? io_in_bits_rm : T_134_rm;
  assign GEN_18 = io_in_valid ? io_in_bits_typ : T_134_typ;
  assign GEN_19 = io_in_valid ? io_in_bits_in1 : T_134_in1;
  assign GEN_20 = io_in_valid ? io_in_bits_in2 : T_134_in2;
  assign GEN_21 = io_in_valid ? io_in_bits_in3 : T_134_in3;
  assign in_valid = T_133;
  assign in_bits_cmd = T_134_cmd;
  assign in_bits_ldst = T_134_ldst;
  assign in_bits_wen = T_134_wen;
  assign in_bits_ren1 = T_134_ren1;
  assign in_bits_ren2 = T_134_ren2;
  assign in_bits_ren3 = T_134_ren3;
  assign in_bits_swap12 = T_134_swap12;
  assign in_bits_swap23 = T_134_swap23;
  assign in_bits_single = T_134_single;
  assign in_bits_fromint = T_134_fromint;
  assign in_bits_toint = T_134_toint;
  assign in_bits_fastpipe = T_134_fastpipe;
  assign in_bits_fma = T_134_fma;
  assign in_bits_div = T_134_div;
  assign in_bits_sqrt = T_134_sqrt;
  assign in_bits_round = T_134_round;
  assign in_bits_wflags = T_134_wflags;
  assign in_bits_rm = T_134_rm;
  assign in_bits_typ = T_134_typ;
  assign in_bits_in1 = T_134_in1;
  assign in_bits_in2 = T_134_in2;
  assign in_bits_in3 = T_134_in3;
  assign T_252 = in_bits_rm[1];
  assign T_253 = in_bits_in1 ^ in_bits_in2;
  assign T_254 = in_bits_rm[0];
  assign T_255 = ~ in_bits_in2;
  assign T_256 = T_254 ? T_255 : in_bits_in2;
  assign signNum = T_252 ? T_253 : T_256;
  assign T_257 = signNum[32];
  assign T_258 = in_bits_in1[31:0];
  assign fsgnj_s = {T_257,T_258};
  assign T_259 = in_bits_in1[64:33];
  assign T_260 = {T_259,fsgnj_s};
  assign T_261 = signNum[64];
  assign T_262 = in_bits_in1[63:0];
  assign T_263 = {T_261,T_262};
  assign fsgnj = in_bits_single ? T_260 : T_263;
  assign mux_data = GEN_41;
  assign mux_exc = GEN_42;
  assign T_272 = in_bits_cmd & 5'hd;
  assign T_273 = 5'h5 == T_272;
  assign T_274 = in_bits_in1[31:29];
  assign T_275 = ~ T_274;
  assign T_277 = T_275 == 3'h0;
  assign T_278 = in_bits_in2[31:29];
  assign T_279 = ~ T_278;
  assign T_281 = T_279 == 3'h0;
  assign T_286 = in_bits_in1[22];
  assign T_288 = T_286 == 1'h0;
  assign T_289 = T_277 & T_288;
  assign T_294 = in_bits_in2[22];
  assign T_296 = T_294 == 1'h0;
  assign T_297 = T_281 & T_296;
  assign T_299 = T_254 != io_lt;
  assign T_301 = T_277 == 1'h0;
  assign T_302 = T_299 & T_301;
  assign T_303 = T_281 | T_302;
  assign T_304 = T_289 | T_297;
  assign T_305 = in_bits_in1[63:61];
  assign T_306 = ~ T_305;
  assign T_308 = T_306 == 3'h0;
  assign T_309 = in_bits_in2[63:61];
  assign T_310 = ~ T_309;
  assign T_312 = T_310 == 3'h0;
  assign T_317 = in_bits_in1[51];
  assign T_319 = T_317 == 1'h0;
  assign T_320 = T_308 & T_319;
  assign T_325 = in_bits_in2[51];
  assign T_327 = T_325 == 1'h0;
  assign T_328 = T_312 & T_327;
  assign T_332 = T_308 == 1'h0;
  assign T_333 = T_299 & T_332;
  assign T_334 = T_312 | T_333;
  assign T_335 = T_320 | T_328;
  assign T_336 = in_bits_single ? T_303 : T_334;
  assign T_337 = in_bits_single ? T_304 : T_335;
  assign GEN_49 = {{4'd0}, T_337};
  assign T_338 = GEN_49 << 4;
  assign T_340 = T_336 == 1'h0;
  assign GEN_22 = T_340 ? in_bits_in2 : in_bits_in1;
  assign GEN_23 = T_273 ? T_338 : 5'h0;
  assign GEN_24 = T_273 ? GEN_22 : fsgnj;
  assign T_343 = in_bits_cmd & 5'h4;
  assign T_344 = 5'h0 == T_343;
  assign RecFNToRecFN_2_clk = clk;
  assign RecFNToRecFN_2_reset = reset;
  assign RecFNToRecFN_2_io_in = in_bits_in1;
  assign RecFNToRecFN_2_io_roundingMode = in_bits_rm[1:0];
  assign T_346 = {32'hffffffff,RecFNToRecFN_2_io_out};
  assign GEN_29 = in_bits_single ? T_346 : GEN_24;
  assign GEN_30 = in_bits_single ? RecFNToRecFN_2_io_exceptionFlags : GEN_23;
  assign T_348 = in_bits_single == 1'h0;
  assign RecFNToRecFN_1_1_clk = clk;
  assign RecFNToRecFN_1_1_reset = reset;
  assign RecFNToRecFN_1_1_io_in = in_bits_in1[32:0];
  assign RecFNToRecFN_1_1_io_roundingMode = in_bits_rm[1:0];
  assign GEN_35 = T_348 ? RecFNToRecFN_1_1_io_out : GEN_29;
  assign GEN_36 = T_348 ? RecFNToRecFN_1_1_io_exceptionFlags : GEN_30;
  assign GEN_41 = T_344 ? GEN_35 : GEN_24;
  assign GEN_42 = T_344 ? GEN_36 : GEN_23;
  assign GEN_47 = in_valid ? mux_data : T_352_data;
  assign GEN_48 = in_valid ? mux_exc : T_352_exc;
  assign T_363_valid = T_351;
  assign T_363_bits_data = T_352_data;
  assign T_363_bits_exc = T_352_exc;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_25 = {1{$random}};
  T_133 = GEN_25[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  T_134_cmd = GEN_26[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  T_134_ldst = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  T_134_wen = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  T_134_ren1 = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  T_134_ren2 = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  T_134_ren3 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  T_134_swap12 = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  T_134_swap23 = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  T_134_single = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  T_134_fromint = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  T_134_toint = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  T_134_fastpipe = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  T_134_fma = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  T_134_div = GEN_45[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  T_134_sqrt = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  T_134_round = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  T_134_wflags = GEN_51[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  T_134_rm = GEN_52[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {1{$random}};
  T_134_typ = GEN_53[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {3{$random}};
  T_134_in1 = GEN_54[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {3{$random}};
  T_134_in2 = GEN_55[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {3{$random}};
  T_134_in3 = GEN_56[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  T_351 = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {3{$random}};
  T_352_data = GEN_58[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  T_352_exc = GEN_59[4:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_133 <= 1'h0;
    end else begin
      T_133 <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_cmd <= io_in_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_ldst <= io_in_bits_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_wen <= io_in_bits_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_ren1 <= io_in_bits_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_ren2 <= io_in_bits_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_ren3 <= io_in_bits_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_swap12 <= io_in_bits_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_swap23 <= io_in_bits_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_single <= io_in_bits_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_fromint <= io_in_bits_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_toint <= io_in_bits_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_fastpipe <= io_in_bits_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_fma <= io_in_bits_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_div <= io_in_bits_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_sqrt <= io_in_bits_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_round <= io_in_bits_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_wflags <= io_in_bits_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_rm <= io_in_bits_rm;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_typ <= io_in_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_in1 <= io_in_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_in2 <= io_in_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        T_134_in3 <= io_in_bits_in3;
      end
    end
    if(reset) begin
      T_351 <= 1'h0;
    end else begin
      T_351 <= in_valid;
    end
    if(1'h0) begin
    end else begin
      if(in_valid) begin
        T_352_data <= mux_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(in_valid) begin
        T_352_exc <= mux_exc;
      end
    end
  end
endmodule
module MulAddRecFN_preMul_1(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [1:0] io_roundingMode,
  output [52:0] io_mulAddA,
  output [52:0] io_mulAddB,
  output [105:0] io_mulAddC,
  output [2:0] io_toPostMul_highExpA,
  output  io_toPostMul_isNaN_isQuietNaNA,
  output [2:0] io_toPostMul_highExpB,
  output  io_toPostMul_isNaN_isQuietNaNB,
  output  io_toPostMul_signProd,
  output  io_toPostMul_isZeroProd,
  output  io_toPostMul_opSignC,
  output [2:0] io_toPostMul_highExpC,
  output  io_toPostMul_isNaN_isQuietNaNC,
  output  io_toPostMul_isCDominant,
  output  io_toPostMul_CAlignDist_0,
  output [7:0] io_toPostMul_CAlignDist,
  output  io_toPostMul_bit0AlignedNegSigC,
  output [54:0] io_toPostMul_highAlignedNegSigC,
  output [13:0] io_toPostMul_sExpSum,
  output [1:0] io_toPostMul_roundingMode
);
  wire  signA;
  wire [11:0] expA;
  wire [51:0] fractA;
  wire [2:0] T_42;
  wire  isZeroA;
  wire  T_45;
  wire [52:0] sigA;
  wire  signB;
  wire [11:0] expB;
  wire [51:0] fractB;
  wire [2:0] T_46;
  wire  isZeroB;
  wire  T_49;
  wire [52:0] sigB;
  wire  T_50;
  wire  T_51;
  wire  opSignC;
  wire [11:0] expC;
  wire [51:0] fractC;
  wire [2:0] T_52;
  wire  isZeroC;
  wire  T_55;
  wire [52:0] sigC;
  wire  T_56;
  wire  T_57;
  wire  signProd;
  wire  isZeroProd;
  wire  T_58;
  wire  T_60;
  wire [2:0] T_64;
  wire [10:0] T_65;
  wire [13:0] T_66;
  wire [13:0] GEN_0;
  wire [14:0] T_67;
  wire [13:0] T_68;
  wire [14:0] T_70;
  wire [13:0] sExpAlignedProd;
  wire  doSubMags;
  wire [13:0] GEN_1;
  wire [14:0] T_71;
  wire [13:0] sNatCAlignDist;
  wire  T_72;
  wire  CAlignDist_floor;
  wire [12:0] T_73;
  wire  T_75;
  wire  CAlignDist_0;
  wire  T_80;
  wire  T_81;
  wire  isCDominant;
  wire  T_85;
  wire [7:0] T_86;
  wire [7:0] T_88;
  wire [7:0] CAlignDist;
  wire [13:0] sExpSum;
  wire  T_89;
  wire [6:0] T_90;
  wire  T_91;
  wire [5:0] T_92;
  wire [64:0] T_95;
  wire [32:0] T_96;
  wire [31:0] T_97;
  wire [15:0] T_102;
  wire [31:0] T_103;
  wire [15:0] T_104;
  wire [31:0] GEN_2;
  wire [31:0] T_105;
  wire [31:0] T_107;
  wire [31:0] T_108;
  wire [23:0] T_112;
  wire [31:0] GEN_3;
  wire [31:0] T_113;
  wire [23:0] T_114;
  wire [31:0] GEN_4;
  wire [31:0] T_115;
  wire [31:0] T_117;
  wire [31:0] T_118;
  wire [27:0] T_122;
  wire [31:0] GEN_5;
  wire [31:0] T_123;
  wire [27:0] T_124;
  wire [31:0] GEN_6;
  wire [31:0] T_125;
  wire [31:0] T_127;
  wire [31:0] T_128;
  wire [29:0] T_132;
  wire [31:0] GEN_7;
  wire [31:0] T_133;
  wire [29:0] T_134;
  wire [31:0] GEN_8;
  wire [31:0] T_135;
  wire [31:0] T_137;
  wire [31:0] T_138;
  wire [30:0] T_142;
  wire [31:0] GEN_9;
  wire [31:0] T_143;
  wire [30:0] T_144;
  wire [31:0] GEN_10;
  wire [31:0] T_145;
  wire [31:0] T_147;
  wire [31:0] T_148;
  wire  T_149;
  wire [32:0] T_150;
  wire [32:0] T_151;
  wire [32:0] T_152;
  wire [32:0] T_153;
  wire [52:0] T_155;
  wire [19:0] T_160;
  wire [15:0] T_161;
  wire [7:0] T_166;
  wire [15:0] T_167;
  wire [7:0] T_168;
  wire [15:0] GEN_11;
  wire [15:0] T_169;
  wire [15:0] T_171;
  wire [15:0] T_172;
  wire [11:0] T_176;
  wire [15:0] GEN_12;
  wire [15:0] T_177;
  wire [11:0] T_178;
  wire [15:0] GEN_13;
  wire [15:0] T_179;
  wire [15:0] T_181;
  wire [15:0] T_182;
  wire [13:0] T_186;
  wire [15:0] GEN_14;
  wire [15:0] T_187;
  wire [13:0] T_188;
  wire [15:0] GEN_15;
  wire [15:0] T_189;
  wire [15:0] T_191;
  wire [15:0] T_192;
  wire [14:0] T_196;
  wire [15:0] GEN_16;
  wire [15:0] T_197;
  wire [14:0] T_198;
  wire [15:0] GEN_17;
  wire [15:0] T_199;
  wire [15:0] T_201;
  wire [15:0] T_202;
  wire [3:0] T_203;
  wire [1:0] T_204;
  wire  T_205;
  wire  T_206;
  wire [1:0] T_207;
  wire [1:0] T_208;
  wire  T_209;
  wire  T_210;
  wire [1:0] T_211;
  wire [3:0] T_212;
  wire [19:0] T_213;
  wire [19:0] T_215;
  wire [52:0] CExtraMask;
  wire [52:0] T_216;
  wire [52:0] negSigC;
  wire [107:0] T_220;
  wire [53:0] T_221;
  wire [161:0] T_222;
  wire [161:0] T_223;
  wire [161:0] T_224;
  wire [52:0] T_225;
  wire  T_227;
  wire  T_228;
  wire [161:0] T_229;
  wire [162:0] T_230;
  wire [161:0] alignedNegSigC;
  wire [105:0] T_231;
  wire  T_233;
  wire  T_235;
  wire  T_237;
  wire  T_238;
  wire [54:0] T_239;
  assign io_mulAddA = sigA;
  assign io_mulAddB = sigB;
  assign io_mulAddC = T_231;
  assign io_toPostMul_highExpA = T_42;
  assign io_toPostMul_isNaN_isQuietNaNA = T_233;
  assign io_toPostMul_highExpB = T_46;
  assign io_toPostMul_isNaN_isQuietNaNB = T_235;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_highExpC = T_52;
  assign io_toPostMul_isNaN_isQuietNaNC = T_237;
  assign io_toPostMul_isCDominant = isCDominant;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_bit0AlignedNegSigC = T_238;
  assign io_toPostMul_highAlignedNegSigC = T_239;
  assign io_toPostMul_sExpSum = sExpSum;
  assign io_toPostMul_roundingMode = io_roundingMode;
  assign signA = io_a[64];
  assign expA = io_a[63:52];
  assign fractA = io_a[51:0];
  assign T_42 = expA[11:9];
  assign isZeroA = T_42 == 3'h0;
  assign T_45 = isZeroA == 1'h0;
  assign sigA = {T_45,fractA};
  assign signB = io_b[64];
  assign expB = io_b[63:52];
  assign fractB = io_b[51:0];
  assign T_46 = expB[11:9];
  assign isZeroB = T_46 == 3'h0;
  assign T_49 = isZeroB == 1'h0;
  assign sigB = {T_49,fractB};
  assign T_50 = io_c[64];
  assign T_51 = io_op[0];
  assign opSignC = T_50 ^ T_51;
  assign expC = io_c[63:52];
  assign fractC = io_c[51:0];
  assign T_52 = expC[11:9];
  assign isZeroC = T_52 == 3'h0;
  assign T_55 = isZeroC == 1'h0;
  assign sigC = {T_55,fractC};
  assign T_56 = signA ^ signB;
  assign T_57 = io_op[1];
  assign signProd = T_56 ^ T_57;
  assign isZeroProd = isZeroA | isZeroB;
  assign T_58 = expB[11];
  assign T_60 = T_58 == 1'h0;
  assign T_64 = T_60 ? 3'h7 : 3'h0;
  assign T_65 = expB[10:0];
  assign T_66 = {T_64,T_65};
  assign GEN_0 = {{2'd0}, expA};
  assign T_67 = GEN_0 + T_66;
  assign T_68 = T_67[13:0];
  assign T_70 = T_68 + 14'h38;
  assign sExpAlignedProd = T_70[13:0];
  assign doSubMags = signProd ^ opSignC;
  assign GEN_1 = {{2'd0}, expC};
  assign T_71 = sExpAlignedProd - GEN_1;
  assign sNatCAlignDist = T_71[13:0];
  assign T_72 = sNatCAlignDist[13];
  assign CAlignDist_floor = isZeroProd | T_72;
  assign T_73 = sNatCAlignDist[12:0];
  assign T_75 = T_73 == 13'h0;
  assign CAlignDist_0 = CAlignDist_floor | T_75;
  assign T_80 = T_73 < 13'h36;
  assign T_81 = CAlignDist_floor | T_80;
  assign isCDominant = T_55 & T_81;
  assign T_85 = T_73 < 13'ha1;
  assign T_86 = sNatCAlignDist[7:0];
  assign T_88 = T_85 ? T_86 : 8'ha1;
  assign CAlignDist = CAlignDist_floor ? 8'h0 : T_88;
  assign sExpSum = CAlignDist_floor ? {{2'd0}, expC} : sExpAlignedProd;
  assign T_89 = CAlignDist[7];
  assign T_90 = CAlignDist[6:0];
  assign T_91 = T_90[6];
  assign T_92 = T_90[5:0];
  assign T_95 = $signed(65'sh10000000000000000) >>> T_92;
  assign T_96 = T_95[63:31];
  assign T_97 = T_96[31:0];
  assign T_102 = T_97[31:16];
  assign T_103 = {{16'd0}, T_102};
  assign T_104 = T_97[15:0];
  assign GEN_2 = {{16'd0}, T_104};
  assign T_105 = GEN_2 << 16;
  assign T_107 = T_105 & 32'hffff0000;
  assign T_108 = T_103 | T_107;
  assign T_112 = T_108[31:8];
  assign GEN_3 = {{8'd0}, T_112};
  assign T_113 = GEN_3 & 32'hff00ff;
  assign T_114 = T_108[23:0];
  assign GEN_4 = {{8'd0}, T_114};
  assign T_115 = GEN_4 << 8;
  assign T_117 = T_115 & 32'hff00ff00;
  assign T_118 = T_113 | T_117;
  assign T_122 = T_118[31:4];
  assign GEN_5 = {{4'd0}, T_122};
  assign T_123 = GEN_5 & 32'hf0f0f0f;
  assign T_124 = T_118[27:0];
  assign GEN_6 = {{4'd0}, T_124};
  assign T_125 = GEN_6 << 4;
  assign T_127 = T_125 & 32'hf0f0f0f0;
  assign T_128 = T_123 | T_127;
  assign T_132 = T_128[31:2];
  assign GEN_7 = {{2'd0}, T_132};
  assign T_133 = GEN_7 & 32'h33333333;
  assign T_134 = T_128[29:0];
  assign GEN_8 = {{2'd0}, T_134};
  assign T_135 = GEN_8 << 2;
  assign T_137 = T_135 & 32'hcccccccc;
  assign T_138 = T_133 | T_137;
  assign T_142 = T_138[31:1];
  assign GEN_9 = {{1'd0}, T_142};
  assign T_143 = GEN_9 & 32'h55555555;
  assign T_144 = T_138[30:0];
  assign GEN_10 = {{1'd0}, T_144};
  assign T_145 = GEN_10 << 1;
  assign T_147 = T_145 & 32'haaaaaaaa;
  assign T_148 = T_143 | T_147;
  assign T_149 = T_96[32];
  assign T_150 = {T_148,T_149};
  assign T_151 = ~ T_150;
  assign T_152 = T_91 ? 33'h0 : T_151;
  assign T_153 = ~ T_152;
  assign T_155 = {T_153,20'hfffff};
  assign T_160 = T_95[19:0];
  assign T_161 = T_160[15:0];
  assign T_166 = T_161[15:8];
  assign T_167 = {{8'd0}, T_166};
  assign T_168 = T_161[7:0];
  assign GEN_11 = {{8'd0}, T_168};
  assign T_169 = GEN_11 << 8;
  assign T_171 = T_169 & 16'hff00;
  assign T_172 = T_167 | T_171;
  assign T_176 = T_172[15:4];
  assign GEN_12 = {{4'd0}, T_176};
  assign T_177 = GEN_12 & 16'hf0f;
  assign T_178 = T_172[11:0];
  assign GEN_13 = {{4'd0}, T_178};
  assign T_179 = GEN_13 << 4;
  assign T_181 = T_179 & 16'hf0f0;
  assign T_182 = T_177 | T_181;
  assign T_186 = T_182[15:2];
  assign GEN_14 = {{2'd0}, T_186};
  assign T_187 = GEN_14 & 16'h3333;
  assign T_188 = T_182[13:0];
  assign GEN_15 = {{2'd0}, T_188};
  assign T_189 = GEN_15 << 2;
  assign T_191 = T_189 & 16'hcccc;
  assign T_192 = T_187 | T_191;
  assign T_196 = T_192[15:1];
  assign GEN_16 = {{1'd0}, T_196};
  assign T_197 = GEN_16 & 16'h5555;
  assign T_198 = T_192[14:0];
  assign GEN_17 = {{1'd0}, T_198};
  assign T_199 = GEN_17 << 1;
  assign T_201 = T_199 & 16'haaaa;
  assign T_202 = T_197 | T_201;
  assign T_203 = T_160[19:16];
  assign T_204 = T_203[1:0];
  assign T_205 = T_204[0];
  assign T_206 = T_204[1];
  assign T_207 = {T_205,T_206};
  assign T_208 = T_203[3:2];
  assign T_209 = T_208[0];
  assign T_210 = T_208[1];
  assign T_211 = {T_209,T_210};
  assign T_212 = {T_207,T_211};
  assign T_213 = {T_202,T_212};
  assign T_215 = T_91 ? T_213 : 20'h0;
  assign CExtraMask = T_89 ? T_155 : {{33'd0}, T_215};
  assign T_216 = ~ sigC;
  assign negSigC = doSubMags ? T_216 : sigC;
  assign T_220 = doSubMags ? 108'hfffffffffffffffffffffffffff : 108'h0;
  assign T_221 = {doSubMags,negSigC};
  assign T_222 = {T_221,T_220};
  assign T_223 = $signed(T_222);
  assign T_224 = $signed(T_223) >>> CAlignDist;
  assign T_225 = sigC & CExtraMask;
  assign T_227 = T_225 != 53'h0;
  assign T_228 = T_227 ^ doSubMags;
  assign T_229 = $unsigned(T_224);
  assign T_230 = {T_229,T_228};
  assign alignedNegSigC = T_230[161:0];
  assign T_231 = alignedNegSigC[106:1];
  assign T_233 = fractA[51];
  assign T_235 = fractB[51];
  assign T_237 = fractC[51];
  assign T_238 = alignedNegSigC[0];
  assign T_239 = alignedNegSigC[161:107];
endmodule
module MulAddRecFN_postMul_1(
  input   clk,
  input   reset,
  input  [2:0] io_fromPreMul_highExpA,
  input   io_fromPreMul_isNaN_isQuietNaNA,
  input  [2:0] io_fromPreMul_highExpB,
  input   io_fromPreMul_isNaN_isQuietNaNB,
  input   io_fromPreMul_signProd,
  input   io_fromPreMul_isZeroProd,
  input   io_fromPreMul_opSignC,
  input  [2:0] io_fromPreMul_highExpC,
  input   io_fromPreMul_isNaN_isQuietNaNC,
  input   io_fromPreMul_isCDominant,
  input   io_fromPreMul_CAlignDist_0,
  input  [7:0] io_fromPreMul_CAlignDist,
  input   io_fromPreMul_bit0AlignedNegSigC,
  input  [54:0] io_fromPreMul_highAlignedNegSigC,
  input  [13:0] io_fromPreMul_sExpSum,
  input  [1:0] io_fromPreMul_roundingMode,
  input  [106:0] io_mulAddResult,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  isZeroA;
  wire [1:0] T_38;
  wire  isSpecialA;
  wire  T_40;
  wire  T_42;
  wire  isInfA;
  wire  isNaNA;
  wire  T_45;
  wire  isSigNaNA;
  wire  isZeroB;
  wire [1:0] T_47;
  wire  isSpecialB;
  wire  T_49;
  wire  T_51;
  wire  isInfB;
  wire  isNaNB;
  wire  T_54;
  wire  isSigNaNB;
  wire  isZeroC;
  wire [1:0] T_56;
  wire  isSpecialC;
  wire  T_58;
  wire  T_60;
  wire  isInfC;
  wire  isNaNC;
  wire  T_63;
  wire  isSigNaNC;
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  doSubMags;
  wire  T_66;
  wire [55:0] T_68;
  wire [54:0] T_69;
  wire [54:0] T_70;
  wire [105:0] T_71;
  wire [160:0] T_72;
  wire [161:0] sigSum;
  wire [107:0] T_74;
  wire [108:0] GEN_0;
  wire [108:0] T_77;
  wire [108:0] T_78;
  wire [107:0] T_80;
  wire [43:0] T_81;
  wire [63:0] T_82;
  wire  T_84;
  wire [11:0] T_85;
  wire [31:0] T_86;
  wire  T_88;
  wire [3:0] T_89;
  wire [7:0] T_90;
  wire  T_92;
  wire  T_93;
  wire  T_95;
  wire  T_97;
  wire [1:0] T_99;
  wire [1:0] T_100;
  wire [3:0] T_101;
  wire [3:0] T_102;
  wire  T_104;
  wire  T_105;
  wire  T_107;
  wire  T_109;
  wire [1:0] T_111;
  wire [1:0] T_112;
  wire  T_113;
  wire  T_115;
  wire  T_117;
  wire [1:0] T_119;
  wire [1:0] T_120;
  wire [1:0] T_121;
  wire [2:0] T_122;
  wire [2:0] T_123;
  wire [3:0] T_124;
  wire [15:0] T_125;
  wire [15:0] T_126;
  wire  T_128;
  wire [7:0] T_129;
  wire [7:0] T_130;
  wire  T_132;
  wire [3:0] T_133;
  wire [3:0] T_134;
  wire  T_136;
  wire  T_137;
  wire  T_139;
  wire  T_141;
  wire [1:0] T_143;
  wire [1:0] T_144;
  wire  T_145;
  wire  T_147;
  wire  T_149;
  wire [1:0] T_151;
  wire [1:0] T_152;
  wire [1:0] T_153;
  wire [2:0] T_154;
  wire [3:0] T_155;
  wire [3:0] T_156;
  wire  T_158;
  wire  T_159;
  wire  T_161;
  wire  T_163;
  wire [1:0] T_165;
  wire [1:0] T_166;
  wire  T_167;
  wire  T_169;
  wire  T_171;
  wire [1:0] T_173;
  wire [1:0] T_174;
  wire [1:0] T_175;
  wire [2:0] T_176;
  wire [2:0] T_177;
  wire [3:0] T_178;
  wire [7:0] T_179;
  wire [7:0] T_180;
  wire  T_182;
  wire [3:0] T_183;
  wire [3:0] T_184;
  wire  T_186;
  wire  T_187;
  wire  T_189;
  wire  T_191;
  wire [1:0] T_193;
  wire [1:0] T_194;
  wire  T_195;
  wire  T_197;
  wire  T_199;
  wire [1:0] T_201;
  wire [1:0] T_202;
  wire [1:0] T_203;
  wire [2:0] T_204;
  wire [3:0] T_205;
  wire [3:0] T_206;
  wire  T_208;
  wire  T_209;
  wire  T_211;
  wire  T_213;
  wire [1:0] T_215;
  wire [1:0] T_216;
  wire  T_217;
  wire  T_219;
  wire  T_221;
  wire [1:0] T_223;
  wire [1:0] T_224;
  wire [1:0] T_225;
  wire [2:0] T_226;
  wire [2:0] T_227;
  wire [3:0] T_228;
  wire [3:0] T_229;
  wire [4:0] T_230;
  wire [4:0] T_231;
  wire [5:0] T_232;
  wire [31:0] T_233;
  wire [31:0] T_234;
  wire  T_236;
  wire [15:0] T_237;
  wire [15:0] T_238;
  wire  T_240;
  wire [7:0] T_241;
  wire [7:0] T_242;
  wire  T_244;
  wire [3:0] T_245;
  wire [3:0] T_246;
  wire  T_248;
  wire  T_249;
  wire  T_251;
  wire  T_253;
  wire [1:0] T_255;
  wire [1:0] T_256;
  wire  T_257;
  wire  T_259;
  wire  T_261;
  wire [1:0] T_263;
  wire [1:0] T_264;
  wire [1:0] T_265;
  wire [2:0] T_266;
  wire [3:0] T_267;
  wire [3:0] T_268;
  wire  T_270;
  wire  T_271;
  wire  T_273;
  wire  T_275;
  wire [1:0] T_277;
  wire [1:0] T_278;
  wire  T_279;
  wire  T_281;
  wire  T_283;
  wire [1:0] T_285;
  wire [1:0] T_286;
  wire [1:0] T_287;
  wire [2:0] T_288;
  wire [2:0] T_289;
  wire [3:0] T_290;
  wire [7:0] T_291;
  wire [7:0] T_292;
  wire  T_294;
  wire [3:0] T_295;
  wire [3:0] T_296;
  wire  T_298;
  wire  T_299;
  wire  T_301;
  wire  T_303;
  wire [1:0] T_305;
  wire [1:0] T_306;
  wire  T_307;
  wire  T_309;
  wire  T_311;
  wire [1:0] T_313;
  wire [1:0] T_314;
  wire [1:0] T_315;
  wire [2:0] T_316;
  wire [3:0] T_317;
  wire [3:0] T_318;
  wire  T_320;
  wire  T_321;
  wire  T_323;
  wire  T_325;
  wire [1:0] T_327;
  wire [1:0] T_328;
  wire  T_329;
  wire  T_331;
  wire  T_333;
  wire [1:0] T_335;
  wire [1:0] T_336;
  wire [1:0] T_337;
  wire [2:0] T_338;
  wire [2:0] T_339;
  wire [3:0] T_340;
  wire [3:0] T_341;
  wire [4:0] T_342;
  wire [15:0] T_343;
  wire [15:0] T_344;
  wire  T_346;
  wire [7:0] T_347;
  wire [7:0] T_348;
  wire  T_350;
  wire [3:0] T_351;
  wire [3:0] T_352;
  wire  T_354;
  wire  T_355;
  wire  T_357;
  wire  T_359;
  wire [1:0] T_361;
  wire [1:0] T_362;
  wire  T_363;
  wire  T_365;
  wire  T_367;
  wire [1:0] T_369;
  wire [1:0] T_370;
  wire [1:0] T_371;
  wire [2:0] T_372;
  wire [3:0] T_373;
  wire [3:0] T_374;
  wire  T_376;
  wire  T_377;
  wire  T_379;
  wire  T_381;
  wire [1:0] T_383;
  wire [1:0] T_384;
  wire  T_385;
  wire  T_387;
  wire  T_389;
  wire [1:0] T_391;
  wire [1:0] T_392;
  wire [1:0] T_393;
  wire [2:0] T_394;
  wire [2:0] T_395;
  wire [3:0] T_396;
  wire [7:0] T_397;
  wire [7:0] T_398;
  wire  T_400;
  wire [3:0] T_401;
  wire [3:0] T_402;
  wire  T_404;
  wire  T_405;
  wire  T_407;
  wire  T_409;
  wire [1:0] T_411;
  wire [1:0] T_412;
  wire  T_413;
  wire  T_415;
  wire  T_417;
  wire [1:0] T_419;
  wire [1:0] T_420;
  wire [1:0] T_421;
  wire [2:0] T_422;
  wire [3:0] T_423;
  wire [3:0] T_424;
  wire  T_426;
  wire  T_427;
  wire  T_429;
  wire  T_431;
  wire [1:0] T_433;
  wire [1:0] T_434;
  wire  T_435;
  wire  T_437;
  wire  T_439;
  wire [1:0] T_441;
  wire [1:0] T_442;
  wire [1:0] T_443;
  wire [2:0] T_444;
  wire [2:0] T_445;
  wire [3:0] T_446;
  wire [3:0] T_447;
  wire [4:0] T_448;
  wire [4:0] T_449;
  wire [5:0] T_450;
  wire [5:0] T_451;
  wire [6:0] T_452;
  wire [7:0] GEN_2;
  wire [8:0] T_453;
  wire [7:0] estNormPos_dist;
  wire [31:0] T_454;
  wire  T_456;
  wire [43:0] T_457;
  wire  T_459;
  wire [1:0] firstReduceSigSum;
  wire [161:0] complSigSum;
  wire [31:0] T_460;
  wire  T_462;
  wire [43:0] T_463;
  wire  T_465;
  wire [1:0] firstReduceComplSigSum;
  wire  T_466;
  wire [8:0] T_468;
  wire [7:0] T_469;
  wire [5:0] T_470;
  wire [7:0] CDom_estNormDist;
  wire  T_472;
  wire  T_473;
  wire  T_475;
  wire  T_476;
  wire [85:0] T_477;
  wire  T_479;
  wire [86:0] T_480;
  wire [86:0] T_482;
  wire  T_486;
  wire [85:0] T_487;
  wire  T_488;
  wire [86:0] T_489;
  wire [86:0] T_491;
  wire [86:0] T_492;
  wire  T_496;
  wire [85:0] T_497;
  wire  T_499;
  wire [86:0] T_500;
  wire [86:0] T_502;
  wire [86:0] T_503;
  wire  T_505;
  wire [85:0] T_506;
  wire  T_507;
  wire [86:0] T_508;
  wire [86:0] T_510;
  wire [86:0] CDom_firstNormAbsSigSum;
  wire [64:0] T_511;
  wire  T_514;
  wire  T_516;
  wire [65:0] T_517;
  wire  T_519;
  wire  T_520;
  wire [85:0] T_524;
  wire [86:0] T_525;
  wire [86:0] T_526;
  wire [85:0] T_527;
  wire [10:0] T_528;
  wire  T_530;
  wire [10:0] T_531;
  wire  T_533;
  wire  T_534;
  wire [86:0] T_535;
  wire  T_536;
  wire  T_537;
  wire [64:0] T_538;
  wire [21:0] T_542;
  wire [86:0] T_543;
  wire [86:0] T_544;
  wire [32:0] T_546;
  wire [53:0] T_550;
  wire [86:0] T_551;
  wire [86:0] T_552;
  wire [86:0] notCDom_pos_firstNormAbsSigSum;
  wire [63:0] T_553;
  wire [64:0] T_555;
  wire [1:0] T_558;
  wire [87:0] GEN_3;
  wire [87:0] T_559;
  wire [87:0] T_560;
  wire [86:0] T_561;
  wire  T_564;
  wire [87:0] T_565;
  wire [65:0] T_568;
  wire [87:0] GEN_4;
  wire [87:0] T_569;
  wire [87:0] T_570;
  wire [33:0] T_572;
  wire [87:0] GEN_5;
  wire [87:0] T_573;
  wire [87:0] T_574;
  wire [87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire  notCDom_signSigSum;
  wire  T_576;
  wire  T_577;
  wire  doNegSignSum;
  wire [7:0] estNormDist;
  wire [87:0] T_579;
  wire [86:0] T_580;
  wire [87:0] cFirstNormAbsSigSum;
  wire  T_582;
  wire  T_584;
  wire  T_585;
  wire  doIncrSig;
  wire [4:0] estNormDist_5;
  wire [4:0] normTo2ShiftDist;
  wire [32:0] T_587;
  wire [30:0] T_588;
  wire [15:0] T_589;
  wire [7:0] T_594;
  wire [15:0] T_595;
  wire [7:0] T_596;
  wire [15:0] GEN_6;
  wire [15:0] T_597;
  wire [15:0] T_599;
  wire [15:0] T_600;
  wire [11:0] T_604;
  wire [15:0] GEN_7;
  wire [15:0] T_605;
  wire [11:0] T_606;
  wire [15:0] GEN_8;
  wire [15:0] T_607;
  wire [15:0] T_609;
  wire [15:0] T_610;
  wire [13:0] T_614;
  wire [15:0] GEN_9;
  wire [15:0] T_615;
  wire [13:0] T_616;
  wire [15:0] GEN_10;
  wire [15:0] T_617;
  wire [15:0] T_619;
  wire [15:0] T_620;
  wire [14:0] T_624;
  wire [15:0] GEN_11;
  wire [15:0] T_625;
  wire [14:0] T_626;
  wire [15:0] GEN_12;
  wire [15:0] T_627;
  wire [15:0] T_629;
  wire [15:0] T_630;
  wire [14:0] T_631;
  wire [7:0] T_632;
  wire [3:0] T_637;
  wire [7:0] T_638;
  wire [3:0] T_639;
  wire [7:0] GEN_13;
  wire [7:0] T_640;
  wire [7:0] T_642;
  wire [7:0] T_643;
  wire [5:0] T_647;
  wire [7:0] GEN_14;
  wire [7:0] T_648;
  wire [5:0] T_649;
  wire [7:0] GEN_15;
  wire [7:0] T_650;
  wire [7:0] T_652;
  wire [7:0] T_653;
  wire [6:0] T_657;
  wire [7:0] GEN_16;
  wire [7:0] T_658;
  wire [6:0] T_659;
  wire [7:0] GEN_17;
  wire [7:0] T_660;
  wire [7:0] T_662;
  wire [7:0] T_663;
  wire [6:0] T_664;
  wire [3:0] T_665;
  wire [1:0] T_666;
  wire  T_667;
  wire  T_668;
  wire [1:0] T_669;
  wire [1:0] T_670;
  wire  T_671;
  wire  T_672;
  wire [1:0] T_673;
  wire [3:0] T_674;
  wire [2:0] T_675;
  wire [1:0] T_676;
  wire  T_677;
  wire  T_678;
  wire [1:0] T_679;
  wire  T_680;
  wire [2:0] T_681;
  wire [6:0] T_682;
  wire [14:0] T_683;
  wire [30:0] T_684;
  wire [31:0] absSigSumExtraMask;
  wire [86:0] T_686;
  wire [86:0] T_687;
  wire [31:0] T_688;
  wire [31:0] T_689;
  wire [31:0] T_690;
  wire  T_692;
  wire [31:0] T_694;
  wire  T_696;
  wire  T_697;
  wire [87:0] T_698;
  wire [56:0] sigX3;
  wire [1:0] T_699;
  wire  sigX3Shift1;
  wire [13:0] GEN_18;
  wire [14:0] T_701;
  wire [13:0] sExpX3;
  wire [2:0] T_702;
  wire  isZeroY;
  wire  T_704;
  wire  signY;
  wire [12:0] sExpX3_13;
  wire  T_705;
  wire [55:0] T_709;
  wire [12:0] T_710;
  wire  T_711;
  wire [11:0] T_712;
  wire  T_713;
  wire [10:0] T_714;
  wire  T_715;
  wire [9:0] T_716;
  wire  T_717;
  wire [8:0] T_718;
  wire  T_720;
  wire [7:0] T_721;
  wire  T_723;
  wire [6:0] T_724;
  wire  T_726;
  wire [5:0] T_727;
  wire [64:0] T_730;
  wire [49:0] T_731;
  wire [31:0] T_732;
  wire [15:0] T_737;
  wire [31:0] T_738;
  wire [15:0] T_739;
  wire [31:0] GEN_19;
  wire [31:0] T_740;
  wire [31:0] T_742;
  wire [31:0] T_743;
  wire [23:0] T_747;
  wire [31:0] GEN_20;
  wire [31:0] T_748;
  wire [23:0] T_749;
  wire [31:0] GEN_21;
  wire [31:0] T_750;
  wire [31:0] T_752;
  wire [31:0] T_753;
  wire [27:0] T_757;
  wire [31:0] GEN_22;
  wire [31:0] T_758;
  wire [27:0] T_759;
  wire [31:0] GEN_23;
  wire [31:0] T_760;
  wire [31:0] T_762;
  wire [31:0] T_763;
  wire [29:0] T_767;
  wire [31:0] GEN_24;
  wire [31:0] T_768;
  wire [29:0] T_769;
  wire [31:0] GEN_25;
  wire [31:0] T_770;
  wire [31:0] T_772;
  wire [31:0] T_773;
  wire [30:0] T_777;
  wire [31:0] GEN_26;
  wire [31:0] T_778;
  wire [30:0] T_779;
  wire [31:0] GEN_27;
  wire [31:0] T_780;
  wire [31:0] T_782;
  wire [31:0] T_783;
  wire [17:0] T_784;
  wire [15:0] T_785;
  wire [7:0] T_790;
  wire [15:0] T_791;
  wire [7:0] T_792;
  wire [15:0] GEN_28;
  wire [15:0] T_793;
  wire [15:0] T_795;
  wire [15:0] T_796;
  wire [11:0] T_800;
  wire [15:0] GEN_29;
  wire [15:0] T_801;
  wire [11:0] T_802;
  wire [15:0] GEN_30;
  wire [15:0] T_803;
  wire [15:0] T_805;
  wire [15:0] T_806;
  wire [13:0] T_810;
  wire [15:0] GEN_31;
  wire [15:0] T_811;
  wire [13:0] T_812;
  wire [15:0] GEN_32;
  wire [15:0] T_813;
  wire [15:0] T_815;
  wire [15:0] T_816;
  wire [14:0] T_820;
  wire [15:0] GEN_33;
  wire [15:0] T_821;
  wire [14:0] T_822;
  wire [15:0] GEN_34;
  wire [15:0] T_823;
  wire [15:0] T_825;
  wire [15:0] T_826;
  wire [1:0] T_827;
  wire  T_828;
  wire  T_829;
  wire [1:0] T_830;
  wire [17:0] T_831;
  wire [49:0] T_832;
  wire [49:0] T_833;
  wire [49:0] T_834;
  wire [49:0] T_835;
  wire [49:0] T_836;
  wire [49:0] T_837;
  wire [49:0] T_838;
  wire [49:0] T_839;
  wire [49:0] T_840;
  wire [49:0] T_841;
  wire [49:0] T_842;
  wire [49:0] T_843;
  wire [49:0] T_844;
  wire [53:0] T_846;
  wire [3:0] T_857;
  wire [1:0] T_858;
  wire  T_859;
  wire  T_860;
  wire [1:0] T_861;
  wire [1:0] T_862;
  wire  T_863;
  wire  T_864;
  wire [1:0] T_865;
  wire [3:0] T_866;
  wire [3:0] T_868;
  wire [3:0] T_870;
  wire [3:0] T_872;
  wire [3:0] T_874;
  wire [53:0] T_875;
  wire [53:0] T_877;
  wire [53:0] T_879;
  wire  T_880;
  wire [53:0] GEN_35;
  wire [53:0] T_881;
  wire [55:0] T_883;
  wire [55:0] roundMask;
  wire [54:0] T_884;
  wire [54:0] T_885;
  wire [55:0] GEN_36;
  wire [55:0] roundPosMask;
  wire [56:0] GEN_37;
  wire [56:0] T_886;
  wire  roundPosBit;
  wire [56:0] GEN_38;
  wire [56:0] T_889;
  wire  anyRoundExtra;
  wire [56:0] T_891;
  wire [56:0] T_893;
  wire  allRoundExtra;
  wire  anyRound;
  wire  allRound;
  wire  roundDirectUp;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire  T_902;
  wire  T_903;
  wire  T_904;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_908;
  wire  T_909;
  wire  T_910;
  wire  roundUp;
  wire  T_914;
  wire  T_915;
  wire  T_916;
  wire  T_917;
  wire  T_919;
  wire  T_920;
  wire  roundEven;
  wire  T_922;
  wire  roundInexact;
  wire [56:0] GEN_40;
  wire [56:0] T_923;
  wire [54:0] T_924;
  wire [55:0] T_926;
  wire [54:0] T_927;
  wire  T_929;
  wire  T_931;
  wire  T_932;
  wire [55:0] T_933;
  wire [56:0] GEN_41;
  wire [56:0] T_934;
  wire [54:0] T_935;
  wire [54:0] T_937;
  wire [54:0] T_939;
  wire [54:0] T_940;
  wire [54:0] T_943;
  wire [54:0] T_945;
  wire [54:0] sigY3;
  wire  T_946;
  wire [14:0] T_948;
  wire [13:0] T_949;
  wire [13:0] T_951;
  wire  T_952;
  wire [13:0] T_954;
  wire [13:0] T_955;
  wire [1:0] T_956;
  wire  T_958;
  wire [14:0] T_960;
  wire [13:0] T_961;
  wire [13:0] T_963;
  wire [13:0] sExpY;
  wire [11:0] expY;
  wire [51:0] T_964;
  wire [51:0] T_965;
  wire [51:0] fractY;
  wire [2:0] T_966;
  wire  overflowY;
  wire  T_969;
  wire  T_970;
  wire  T_973;
  wire  T_974;
  wire  totalUnderflowY;
  wire [10:0] T_978;
  wire [12:0] GEN_42;
  wire  T_979;
  wire  T_980;
  wire  underflowY;
  wire  T_981;
  wire  T_983;
  wire  T_984;
  wire  roundMagUp;
  wire  overflowY_roundMagUp;
  wire  mulSpecial;
  wire  addSpecial;
  wire  notSpecial_addZeros;
  wire  T_986;
  wire  T_988;
  wire  commonCase;
  wire  T_989;
  wire  T_990;
  wire  T_991;
  wire  T_993;
  wire  T_995;
  wire  T_996;
  wire  T_997;
  wire  T_998;
  wire  T_999;
  wire  T_1000;
  wire  notSigNaN_invalid;
  wire  T_1001;
  wire  T_1002;
  wire  invalid;
  wire  overflow;
  wire  underflow;
  wire  T_1003;
  wire  inexact;
  wire  T_1004;
  wire  notSpecial_isZeroOut;
  wire  T_1005;
  wire  pegMinFiniteMagOut;
  wire  T_1007;
  wire  pegMaxFiniteMagOut;
  wire  T_1009;
  wire  T_1010;
  wire  notNaN_isInfOut;
  wire  T_1011;
  wire  T_1012;
  wire  isNaNOut;
  wire  T_1015;
  wire  T_1017;
  wire  T_1018;
  wire  T_1019;
  wire  T_1020;
  wire  T_1022;
  wire  T_1023;
  wire  T_1024;
  wire  T_1025;
  wire  T_1028;
  wire  T_1029;
  wire  T_1030;
  wire  uncommonCaseSignOut;
  wire  T_1032;
  wire  T_1033;
  wire  T_1034;
  wire  signOut;
  wire [11:0] T_1037;
  wire [11:0] T_1038;
  wire [11:0] T_1039;
  wire [11:0] T_1043;
  wire [11:0] T_1044;
  wire [11:0] T_1045;
  wire [11:0] T_1048;
  wire [11:0] T_1049;
  wire [11:0] T_1050;
  wire [11:0] T_1053;
  wire [11:0] T_1054;
  wire [11:0] T_1055;
  wire [11:0] T_1058;
  wire [11:0] T_1059;
  wire [11:0] T_1062;
  wire [11:0] T_1063;
  wire [11:0] T_1066;
  wire [11:0] T_1067;
  wire [11:0] T_1070;
  wire [11:0] expOut;
  wire  T_1071;
  wire  T_1072;
  wire [51:0] T_1076;
  wire [51:0] T_1077;
  wire [51:0] T_1081;
  wire [51:0] fractOut;
  wire [12:0] T_1082;
  wire [64:0] T_1083;
  wire [1:0] T_1085;
  wire [1:0] T_1086;
  wire [2:0] T_1087;
  wire [4:0] T_1088;
  assign io_out = T_1083;
  assign io_exceptionFlags = T_1088;
  assign isZeroA = io_fromPreMul_highExpA == 3'h0;
  assign T_38 = io_fromPreMul_highExpA[2:1];
  assign isSpecialA = T_38 == 2'h3;
  assign T_40 = io_fromPreMul_highExpA[0];
  assign T_42 = T_40 == 1'h0;
  assign isInfA = isSpecialA & T_42;
  assign isNaNA = isSpecialA & T_40;
  assign T_45 = io_fromPreMul_isNaN_isQuietNaNA == 1'h0;
  assign isSigNaNA = isNaNA & T_45;
  assign isZeroB = io_fromPreMul_highExpB == 3'h0;
  assign T_47 = io_fromPreMul_highExpB[2:1];
  assign isSpecialB = T_47 == 2'h3;
  assign T_49 = io_fromPreMul_highExpB[0];
  assign T_51 = T_49 == 1'h0;
  assign isInfB = isSpecialB & T_51;
  assign isNaNB = isSpecialB & T_49;
  assign T_54 = io_fromPreMul_isNaN_isQuietNaNB == 1'h0;
  assign isSigNaNB = isNaNB & T_54;
  assign isZeroC = io_fromPreMul_highExpC == 3'h0;
  assign T_56 = io_fromPreMul_highExpC[2:1];
  assign isSpecialC = T_56 == 2'h3;
  assign T_58 = io_fromPreMul_highExpC[0];
  assign T_60 = T_58 == 1'h0;
  assign isInfC = isSpecialC & T_60;
  assign isNaNC = isSpecialC & T_58;
  assign T_63 = io_fromPreMul_isNaN_isQuietNaNC == 1'h0;
  assign isSigNaNC = isNaNC & T_63;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T_66 = io_mulAddResult[106];
  assign T_68 = io_fromPreMul_highAlignedNegSigC + 55'h1;
  assign T_69 = T_68[54:0];
  assign T_70 = T_66 ? T_69 : io_fromPreMul_highAlignedNegSigC;
  assign T_71 = io_mulAddResult[105:0];
  assign T_72 = {T_70,T_71};
  assign sigSum = {T_72,io_fromPreMul_bit0AlignedNegSigC};
  assign T_74 = sigSum[108:1];
  assign GEN_0 = {{1'd0}, T_74};
  assign T_77 = GEN_0 << 1;
  assign T_78 = GEN_0 ^ T_77;
  assign T_80 = T_78[107:0];
  assign T_81 = T_80[107:64];
  assign T_82 = T_80[63:0];
  assign T_84 = T_81 != 44'h0;
  assign T_85 = T_81[43:32];
  assign T_86 = T_81[31:0];
  assign T_88 = T_85 != 12'h0;
  assign T_89 = T_85[11:8];
  assign T_90 = T_85[7:0];
  assign T_92 = T_89 != 4'h0;
  assign T_93 = T_89[3];
  assign T_95 = T_89[2];
  assign T_97 = T_89[1];
  assign T_99 = T_95 ? 2'h2 : {{1'd0}, T_97};
  assign T_100 = T_93 ? 2'h3 : T_99;
  assign T_101 = T_90[7:4];
  assign T_102 = T_90[3:0];
  assign T_104 = T_101 != 4'h0;
  assign T_105 = T_101[3];
  assign T_107 = T_101[2];
  assign T_109 = T_101[1];
  assign T_111 = T_107 ? 2'h2 : {{1'd0}, T_109};
  assign T_112 = T_105 ? 2'h3 : T_111;
  assign T_113 = T_102[3];
  assign T_115 = T_102[2];
  assign T_117 = T_102[1];
  assign T_119 = T_115 ? 2'h2 : {{1'd0}, T_117};
  assign T_120 = T_113 ? 2'h3 : T_119;
  assign T_121 = T_104 ? T_112 : T_120;
  assign T_122 = {T_104,T_121};
  assign T_123 = T_92 ? {{1'd0}, T_100} : T_122;
  assign T_124 = {T_92,T_123};
  assign T_125 = T_86[31:16];
  assign T_126 = T_86[15:0];
  assign T_128 = T_125 != 16'h0;
  assign T_129 = T_125[15:8];
  assign T_130 = T_125[7:0];
  assign T_132 = T_129 != 8'h0;
  assign T_133 = T_129[7:4];
  assign T_134 = T_129[3:0];
  assign T_136 = T_133 != 4'h0;
  assign T_137 = T_133[3];
  assign T_139 = T_133[2];
  assign T_141 = T_133[1];
  assign T_143 = T_139 ? 2'h2 : {{1'd0}, T_141};
  assign T_144 = T_137 ? 2'h3 : T_143;
  assign T_145 = T_134[3];
  assign T_147 = T_134[2];
  assign T_149 = T_134[1];
  assign T_151 = T_147 ? 2'h2 : {{1'd0}, T_149};
  assign T_152 = T_145 ? 2'h3 : T_151;
  assign T_153 = T_136 ? T_144 : T_152;
  assign T_154 = {T_136,T_153};
  assign T_155 = T_130[7:4];
  assign T_156 = T_130[3:0];
  assign T_158 = T_155 != 4'h0;
  assign T_159 = T_155[3];
  assign T_161 = T_155[2];
  assign T_163 = T_155[1];
  assign T_165 = T_161 ? 2'h2 : {{1'd0}, T_163};
  assign T_166 = T_159 ? 2'h3 : T_165;
  assign T_167 = T_156[3];
  assign T_169 = T_156[2];
  assign T_171 = T_156[1];
  assign T_173 = T_169 ? 2'h2 : {{1'd0}, T_171};
  assign T_174 = T_167 ? 2'h3 : T_173;
  assign T_175 = T_158 ? T_166 : T_174;
  assign T_176 = {T_158,T_175};
  assign T_177 = T_132 ? T_154 : T_176;
  assign T_178 = {T_132,T_177};
  assign T_179 = T_126[15:8];
  assign T_180 = T_126[7:0];
  assign T_182 = T_179 != 8'h0;
  assign T_183 = T_179[7:4];
  assign T_184 = T_179[3:0];
  assign T_186 = T_183 != 4'h0;
  assign T_187 = T_183[3];
  assign T_189 = T_183[2];
  assign T_191 = T_183[1];
  assign T_193 = T_189 ? 2'h2 : {{1'd0}, T_191};
  assign T_194 = T_187 ? 2'h3 : T_193;
  assign T_195 = T_184[3];
  assign T_197 = T_184[2];
  assign T_199 = T_184[1];
  assign T_201 = T_197 ? 2'h2 : {{1'd0}, T_199};
  assign T_202 = T_195 ? 2'h3 : T_201;
  assign T_203 = T_186 ? T_194 : T_202;
  assign T_204 = {T_186,T_203};
  assign T_205 = T_180[7:4];
  assign T_206 = T_180[3:0];
  assign T_208 = T_205 != 4'h0;
  assign T_209 = T_205[3];
  assign T_211 = T_205[2];
  assign T_213 = T_205[1];
  assign T_215 = T_211 ? 2'h2 : {{1'd0}, T_213};
  assign T_216 = T_209 ? 2'h3 : T_215;
  assign T_217 = T_206[3];
  assign T_219 = T_206[2];
  assign T_221 = T_206[1];
  assign T_223 = T_219 ? 2'h2 : {{1'd0}, T_221};
  assign T_224 = T_217 ? 2'h3 : T_223;
  assign T_225 = T_208 ? T_216 : T_224;
  assign T_226 = {T_208,T_225};
  assign T_227 = T_182 ? T_204 : T_226;
  assign T_228 = {T_182,T_227};
  assign T_229 = T_128 ? T_178 : T_228;
  assign T_230 = {T_128,T_229};
  assign T_231 = T_88 ? {{1'd0}, T_124} : T_230;
  assign T_232 = {T_88,T_231};
  assign T_233 = T_82[63:32];
  assign T_234 = T_82[31:0];
  assign T_236 = T_233 != 32'h0;
  assign T_237 = T_233[31:16];
  assign T_238 = T_233[15:0];
  assign T_240 = T_237 != 16'h0;
  assign T_241 = T_237[15:8];
  assign T_242 = T_237[7:0];
  assign T_244 = T_241 != 8'h0;
  assign T_245 = T_241[7:4];
  assign T_246 = T_241[3:0];
  assign T_248 = T_245 != 4'h0;
  assign T_249 = T_245[3];
  assign T_251 = T_245[2];
  assign T_253 = T_245[1];
  assign T_255 = T_251 ? 2'h2 : {{1'd0}, T_253};
  assign T_256 = T_249 ? 2'h3 : T_255;
  assign T_257 = T_246[3];
  assign T_259 = T_246[2];
  assign T_261 = T_246[1];
  assign T_263 = T_259 ? 2'h2 : {{1'd0}, T_261};
  assign T_264 = T_257 ? 2'h3 : T_263;
  assign T_265 = T_248 ? T_256 : T_264;
  assign T_266 = {T_248,T_265};
  assign T_267 = T_242[7:4];
  assign T_268 = T_242[3:0];
  assign T_270 = T_267 != 4'h0;
  assign T_271 = T_267[3];
  assign T_273 = T_267[2];
  assign T_275 = T_267[1];
  assign T_277 = T_273 ? 2'h2 : {{1'd0}, T_275};
  assign T_278 = T_271 ? 2'h3 : T_277;
  assign T_279 = T_268[3];
  assign T_281 = T_268[2];
  assign T_283 = T_268[1];
  assign T_285 = T_281 ? 2'h2 : {{1'd0}, T_283};
  assign T_286 = T_279 ? 2'h3 : T_285;
  assign T_287 = T_270 ? T_278 : T_286;
  assign T_288 = {T_270,T_287};
  assign T_289 = T_244 ? T_266 : T_288;
  assign T_290 = {T_244,T_289};
  assign T_291 = T_238[15:8];
  assign T_292 = T_238[7:0];
  assign T_294 = T_291 != 8'h0;
  assign T_295 = T_291[7:4];
  assign T_296 = T_291[3:0];
  assign T_298 = T_295 != 4'h0;
  assign T_299 = T_295[3];
  assign T_301 = T_295[2];
  assign T_303 = T_295[1];
  assign T_305 = T_301 ? 2'h2 : {{1'd0}, T_303};
  assign T_306 = T_299 ? 2'h3 : T_305;
  assign T_307 = T_296[3];
  assign T_309 = T_296[2];
  assign T_311 = T_296[1];
  assign T_313 = T_309 ? 2'h2 : {{1'd0}, T_311};
  assign T_314 = T_307 ? 2'h3 : T_313;
  assign T_315 = T_298 ? T_306 : T_314;
  assign T_316 = {T_298,T_315};
  assign T_317 = T_292[7:4];
  assign T_318 = T_292[3:0];
  assign T_320 = T_317 != 4'h0;
  assign T_321 = T_317[3];
  assign T_323 = T_317[2];
  assign T_325 = T_317[1];
  assign T_327 = T_323 ? 2'h2 : {{1'd0}, T_325};
  assign T_328 = T_321 ? 2'h3 : T_327;
  assign T_329 = T_318[3];
  assign T_331 = T_318[2];
  assign T_333 = T_318[1];
  assign T_335 = T_331 ? 2'h2 : {{1'd0}, T_333};
  assign T_336 = T_329 ? 2'h3 : T_335;
  assign T_337 = T_320 ? T_328 : T_336;
  assign T_338 = {T_320,T_337};
  assign T_339 = T_294 ? T_316 : T_338;
  assign T_340 = {T_294,T_339};
  assign T_341 = T_240 ? T_290 : T_340;
  assign T_342 = {T_240,T_341};
  assign T_343 = T_234[31:16];
  assign T_344 = T_234[15:0];
  assign T_346 = T_343 != 16'h0;
  assign T_347 = T_343[15:8];
  assign T_348 = T_343[7:0];
  assign T_350 = T_347 != 8'h0;
  assign T_351 = T_347[7:4];
  assign T_352 = T_347[3:0];
  assign T_354 = T_351 != 4'h0;
  assign T_355 = T_351[3];
  assign T_357 = T_351[2];
  assign T_359 = T_351[1];
  assign T_361 = T_357 ? 2'h2 : {{1'd0}, T_359};
  assign T_362 = T_355 ? 2'h3 : T_361;
  assign T_363 = T_352[3];
  assign T_365 = T_352[2];
  assign T_367 = T_352[1];
  assign T_369 = T_365 ? 2'h2 : {{1'd0}, T_367};
  assign T_370 = T_363 ? 2'h3 : T_369;
  assign T_371 = T_354 ? T_362 : T_370;
  assign T_372 = {T_354,T_371};
  assign T_373 = T_348[7:4];
  assign T_374 = T_348[3:0];
  assign T_376 = T_373 != 4'h0;
  assign T_377 = T_373[3];
  assign T_379 = T_373[2];
  assign T_381 = T_373[1];
  assign T_383 = T_379 ? 2'h2 : {{1'd0}, T_381};
  assign T_384 = T_377 ? 2'h3 : T_383;
  assign T_385 = T_374[3];
  assign T_387 = T_374[2];
  assign T_389 = T_374[1];
  assign T_391 = T_387 ? 2'h2 : {{1'd0}, T_389};
  assign T_392 = T_385 ? 2'h3 : T_391;
  assign T_393 = T_376 ? T_384 : T_392;
  assign T_394 = {T_376,T_393};
  assign T_395 = T_350 ? T_372 : T_394;
  assign T_396 = {T_350,T_395};
  assign T_397 = T_344[15:8];
  assign T_398 = T_344[7:0];
  assign T_400 = T_397 != 8'h0;
  assign T_401 = T_397[7:4];
  assign T_402 = T_397[3:0];
  assign T_404 = T_401 != 4'h0;
  assign T_405 = T_401[3];
  assign T_407 = T_401[2];
  assign T_409 = T_401[1];
  assign T_411 = T_407 ? 2'h2 : {{1'd0}, T_409};
  assign T_412 = T_405 ? 2'h3 : T_411;
  assign T_413 = T_402[3];
  assign T_415 = T_402[2];
  assign T_417 = T_402[1];
  assign T_419 = T_415 ? 2'h2 : {{1'd0}, T_417};
  assign T_420 = T_413 ? 2'h3 : T_419;
  assign T_421 = T_404 ? T_412 : T_420;
  assign T_422 = {T_404,T_421};
  assign T_423 = T_398[7:4];
  assign T_424 = T_398[3:0];
  assign T_426 = T_423 != 4'h0;
  assign T_427 = T_423[3];
  assign T_429 = T_423[2];
  assign T_431 = T_423[1];
  assign T_433 = T_429 ? 2'h2 : {{1'd0}, T_431};
  assign T_434 = T_427 ? 2'h3 : T_433;
  assign T_435 = T_424[3];
  assign T_437 = T_424[2];
  assign T_439 = T_424[1];
  assign T_441 = T_437 ? 2'h2 : {{1'd0}, T_439};
  assign T_442 = T_435 ? 2'h3 : T_441;
  assign T_443 = T_426 ? T_434 : T_442;
  assign T_444 = {T_426,T_443};
  assign T_445 = T_400 ? T_422 : T_444;
  assign T_446 = {T_400,T_445};
  assign T_447 = T_346 ? T_396 : T_446;
  assign T_448 = {T_346,T_447};
  assign T_449 = T_236 ? T_342 : T_448;
  assign T_450 = {T_236,T_449};
  assign T_451 = T_84 ? T_232 : T_450;
  assign T_452 = {T_84,T_451};
  assign GEN_2 = {{1'd0}, T_452};
  assign T_453 = 8'ha0 - GEN_2;
  assign estNormPos_dist = T_453[7:0];
  assign T_454 = sigSum[75:44];
  assign T_456 = T_454 != 32'h0;
  assign T_457 = sigSum[43:0];
  assign T_459 = T_457 != 44'h0;
  assign firstReduceSigSum = {T_456,T_459};
  assign complSigSum = ~ sigSum;
  assign T_460 = complSigSum[75:44];
  assign T_462 = T_460 != 32'h0;
  assign T_463 = complSigSum[43:0];
  assign T_465 = T_463 != 44'h0;
  assign firstReduceComplSigSum = {T_462,T_465};
  assign T_466 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign T_468 = io_fromPreMul_CAlignDist - 8'h1;
  assign T_469 = T_468[7:0];
  assign T_470 = T_469[5:0];
  assign CDom_estNormDist = T_466 ? io_fromPreMul_CAlignDist : {{2'd0}, T_470};
  assign T_472 = doSubMags == 1'h0;
  assign T_473 = CDom_estNormDist[5];
  assign T_475 = T_473 == 1'h0;
  assign T_476 = T_472 & T_475;
  assign T_477 = sigSum[161:76];
  assign T_479 = firstReduceSigSum != 2'h0;
  assign T_480 = {T_477,T_479};
  assign T_482 = T_476 ? T_480 : 87'h0;
  assign T_486 = T_472 & T_473;
  assign T_487 = sigSum[129:44];
  assign T_488 = firstReduceSigSum[0];
  assign T_489 = {T_487,T_488};
  assign T_491 = T_486 ? T_489 : 87'h0;
  assign T_492 = T_482 | T_491;
  assign T_496 = doSubMags & T_475;
  assign T_497 = complSigSum[161:76];
  assign T_499 = firstReduceComplSigSum != 2'h0;
  assign T_500 = {T_497,T_499};
  assign T_502 = T_496 ? T_500 : 87'h0;
  assign T_503 = T_492 | T_502;
  assign T_505 = doSubMags & T_473;
  assign T_506 = complSigSum[129:44];
  assign T_507 = firstReduceComplSigSum[0];
  assign T_508 = {T_506,T_507};
  assign T_510 = T_505 ? T_508 : 87'h0;
  assign CDom_firstNormAbsSigSum = T_503 | T_510;
  assign T_511 = sigSum[108:44];
  assign T_514 = T_507 == 1'h0;
  assign T_516 = doSubMags ? T_514 : T_488;
  assign T_517 = {T_511,T_516};
  assign T_519 = estNormPos_dist[4];
  assign T_520 = sigSum[1];
  assign T_524 = doSubMags ? 86'h3fffffffffffffffffffff : 86'h0;
  assign T_525 = {T_520,T_524};
  assign T_526 = T_519 ? {{21'd0}, T_517} : T_525;
  assign T_527 = sigSum[97:12];
  assign T_528 = complSigSum[11:1];
  assign T_530 = T_528 == 11'h0;
  assign T_531 = sigSum[11:1];
  assign T_533 = T_531 != 11'h0;
  assign T_534 = doSubMags ? T_530 : T_533;
  assign T_535 = {T_527,T_534};
  assign T_536 = estNormPos_dist[6];
  assign T_537 = estNormPos_dist[5];
  assign T_538 = sigSum[65:1];
  assign T_542 = doSubMags ? 22'h3fffff : 22'h0;
  assign T_543 = {T_538,T_542};
  assign T_544 = T_537 ? T_543 : T_535;
  assign T_546 = sigSum[33:1];
  assign T_550 = doSubMags ? 54'h3fffffffffffff : 54'h0;
  assign T_551 = {T_546,T_550};
  assign T_552 = T_537 ? T_526 : T_551;
  assign notCDom_pos_firstNormAbsSigSum = T_536 ? T_544 : T_552;
  assign T_553 = complSigSum[107:44];
  assign T_555 = {T_553,T_507};
  assign T_558 = complSigSum[2:1];
  assign GEN_3 = {{86'd0}, T_558};
  assign T_559 = GEN_3 << 86;
  assign T_560 = T_519 ? {{23'd0}, T_555} : T_559;
  assign T_561 = complSigSum[98:12];
  assign T_564 = T_528 != 11'h0;
  assign T_565 = {T_561,T_564};
  assign T_568 = complSigSum[66:1];
  assign GEN_4 = {{22'd0}, T_568};
  assign T_569 = GEN_4 << 22;
  assign T_570 = T_537 ? T_569 : T_565;
  assign T_572 = complSigSum[34:1];
  assign GEN_5 = {{54'd0}, T_572};
  assign T_573 = GEN_5 << 54;
  assign T_574 = T_537 ? T_560 : T_573;
  assign notCDom_neg_cFirstNormAbsSigSum = T_536 ? T_570 : T_574;
  assign notCDom_signSigSum = sigSum[109];
  assign T_576 = isZeroC == 1'h0;
  assign T_577 = doSubMags & T_576;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T_577 : notCDom_signSigSum;
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : estNormPos_dist;
  assign T_579 = io_fromPreMul_isCDominant ? {{1'd0}, CDom_firstNormAbsSigSum} : notCDom_neg_cFirstNormAbsSigSum;
  assign T_580 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T_579 : {{1'd0}, T_580};
  assign T_582 = io_fromPreMul_isCDominant == 1'h0;
  assign T_584 = notCDom_signSigSum == 1'h0;
  assign T_585 = T_582 & T_584;
  assign doIncrSig = T_585 & doSubMags;
  assign estNormDist_5 = estNormDist[4:0];
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign T_587 = $signed(33'sh100000000) >>> normTo2ShiftDist;
  assign T_588 = T_587[31:1];
  assign T_589 = T_588[15:0];
  assign T_594 = T_589[15:8];
  assign T_595 = {{8'd0}, T_594};
  assign T_596 = T_589[7:0];
  assign GEN_6 = {{8'd0}, T_596};
  assign T_597 = GEN_6 << 8;
  assign T_599 = T_597 & 16'hff00;
  assign T_600 = T_595 | T_599;
  assign T_604 = T_600[15:4];
  assign GEN_7 = {{4'd0}, T_604};
  assign T_605 = GEN_7 & 16'hf0f;
  assign T_606 = T_600[11:0];
  assign GEN_8 = {{4'd0}, T_606};
  assign T_607 = GEN_8 << 4;
  assign T_609 = T_607 & 16'hf0f0;
  assign T_610 = T_605 | T_609;
  assign T_614 = T_610[15:2];
  assign GEN_9 = {{2'd0}, T_614};
  assign T_615 = GEN_9 & 16'h3333;
  assign T_616 = T_610[13:0];
  assign GEN_10 = {{2'd0}, T_616};
  assign T_617 = GEN_10 << 2;
  assign T_619 = T_617 & 16'hcccc;
  assign T_620 = T_615 | T_619;
  assign T_624 = T_620[15:1];
  assign GEN_11 = {{1'd0}, T_624};
  assign T_625 = GEN_11 & 16'h5555;
  assign T_626 = T_620[14:0];
  assign GEN_12 = {{1'd0}, T_626};
  assign T_627 = GEN_12 << 1;
  assign T_629 = T_627 & 16'haaaa;
  assign T_630 = T_625 | T_629;
  assign T_631 = T_588[30:16];
  assign T_632 = T_631[7:0];
  assign T_637 = T_632[7:4];
  assign T_638 = {{4'd0}, T_637};
  assign T_639 = T_632[3:0];
  assign GEN_13 = {{4'd0}, T_639};
  assign T_640 = GEN_13 << 4;
  assign T_642 = T_640 & 8'hf0;
  assign T_643 = T_638 | T_642;
  assign T_647 = T_643[7:2];
  assign GEN_14 = {{2'd0}, T_647};
  assign T_648 = GEN_14 & 8'h33;
  assign T_649 = T_643[5:0];
  assign GEN_15 = {{2'd0}, T_649};
  assign T_650 = GEN_15 << 2;
  assign T_652 = T_650 & 8'hcc;
  assign T_653 = T_648 | T_652;
  assign T_657 = T_653[7:1];
  assign GEN_16 = {{1'd0}, T_657};
  assign T_658 = GEN_16 & 8'h55;
  assign T_659 = T_653[6:0];
  assign GEN_17 = {{1'd0}, T_659};
  assign T_660 = GEN_17 << 1;
  assign T_662 = T_660 & 8'haa;
  assign T_663 = T_658 | T_662;
  assign T_664 = T_631[14:8];
  assign T_665 = T_664[3:0];
  assign T_666 = T_665[1:0];
  assign T_667 = T_666[0];
  assign T_668 = T_666[1];
  assign T_669 = {T_667,T_668};
  assign T_670 = T_665[3:2];
  assign T_671 = T_670[0];
  assign T_672 = T_670[1];
  assign T_673 = {T_671,T_672};
  assign T_674 = {T_669,T_673};
  assign T_675 = T_664[6:4];
  assign T_676 = T_675[1:0];
  assign T_677 = T_676[0];
  assign T_678 = T_676[1];
  assign T_679 = {T_677,T_678};
  assign T_680 = T_675[2];
  assign T_681 = {T_679,T_680};
  assign T_682 = {T_674,T_681};
  assign T_683 = {T_663,T_682};
  assign T_684 = {T_630,T_683};
  assign absSigSumExtraMask = {T_684,1'h1};
  assign T_686 = cFirstNormAbsSigSum[87:1];
  assign T_687 = T_686 >> normTo2ShiftDist;
  assign T_688 = cFirstNormAbsSigSum[31:0];
  assign T_689 = ~ T_688;
  assign T_690 = T_689 & absSigSumExtraMask;
  assign T_692 = T_690 == 32'h0;
  assign T_694 = T_688 & absSigSumExtraMask;
  assign T_696 = T_694 != 32'h0;
  assign T_697 = doIncrSig ? T_692 : T_696;
  assign T_698 = {T_687,T_697};
  assign sigX3 = T_698[56:0];
  assign T_699 = sigX3[56:55];
  assign sigX3Shift1 = T_699 == 2'h0;
  assign GEN_18 = {{6'd0}, estNormDist};
  assign T_701 = io_fromPreMul_sExpSum - GEN_18;
  assign sExpX3 = T_701[13:0];
  assign T_702 = sigX3[56:54];
  assign isZeroY = T_702 == 3'h0;
  assign T_704 = io_fromPreMul_signProd ^ doNegSignSum;
  assign signY = isZeroY ? roundingMode_min : T_704;
  assign sExpX3_13 = sExpX3[12:0];
  assign T_705 = sExpX3[13];
  assign T_709 = T_705 ? 56'hffffffffffffff : 56'h0;
  assign T_710 = ~ sExpX3_13;
  assign T_711 = T_710[12];
  assign T_712 = T_710[11:0];
  assign T_713 = T_712[11];
  assign T_714 = T_712[10:0];
  assign T_715 = T_714[10];
  assign T_716 = T_714[9:0];
  assign T_717 = T_716[9];
  assign T_718 = T_716[8:0];
  assign T_720 = T_718[8];
  assign T_721 = T_718[7:0];
  assign T_723 = T_721[7];
  assign T_724 = T_721[6:0];
  assign T_726 = T_724[6];
  assign T_727 = T_724[5:0];
  assign T_730 = $signed(65'sh10000000000000000) >>> T_727;
  assign T_731 = T_730[63:14];
  assign T_732 = T_731[31:0];
  assign T_737 = T_732[31:16];
  assign T_738 = {{16'd0}, T_737};
  assign T_739 = T_732[15:0];
  assign GEN_19 = {{16'd0}, T_739};
  assign T_740 = GEN_19 << 16;
  assign T_742 = T_740 & 32'hffff0000;
  assign T_743 = T_738 | T_742;
  assign T_747 = T_743[31:8];
  assign GEN_20 = {{8'd0}, T_747};
  assign T_748 = GEN_20 & 32'hff00ff;
  assign T_749 = T_743[23:0];
  assign GEN_21 = {{8'd0}, T_749};
  assign T_750 = GEN_21 << 8;
  assign T_752 = T_750 & 32'hff00ff00;
  assign T_753 = T_748 | T_752;
  assign T_757 = T_753[31:4];
  assign GEN_22 = {{4'd0}, T_757};
  assign T_758 = GEN_22 & 32'hf0f0f0f;
  assign T_759 = T_753[27:0];
  assign GEN_23 = {{4'd0}, T_759};
  assign T_760 = GEN_23 << 4;
  assign T_762 = T_760 & 32'hf0f0f0f0;
  assign T_763 = T_758 | T_762;
  assign T_767 = T_763[31:2];
  assign GEN_24 = {{2'd0}, T_767};
  assign T_768 = GEN_24 & 32'h33333333;
  assign T_769 = T_763[29:0];
  assign GEN_25 = {{2'd0}, T_769};
  assign T_770 = GEN_25 << 2;
  assign T_772 = T_770 & 32'hcccccccc;
  assign T_773 = T_768 | T_772;
  assign T_777 = T_773[31:1];
  assign GEN_26 = {{1'd0}, T_777};
  assign T_778 = GEN_26 & 32'h55555555;
  assign T_779 = T_773[30:0];
  assign GEN_27 = {{1'd0}, T_779};
  assign T_780 = GEN_27 << 1;
  assign T_782 = T_780 & 32'haaaaaaaa;
  assign T_783 = T_778 | T_782;
  assign T_784 = T_731[49:32];
  assign T_785 = T_784[15:0];
  assign T_790 = T_785[15:8];
  assign T_791 = {{8'd0}, T_790};
  assign T_792 = T_785[7:0];
  assign GEN_28 = {{8'd0}, T_792};
  assign T_793 = GEN_28 << 8;
  assign T_795 = T_793 & 16'hff00;
  assign T_796 = T_791 | T_795;
  assign T_800 = T_796[15:4];
  assign GEN_29 = {{4'd0}, T_800};
  assign T_801 = GEN_29 & 16'hf0f;
  assign T_802 = T_796[11:0];
  assign GEN_30 = {{4'd0}, T_802};
  assign T_803 = GEN_30 << 4;
  assign T_805 = T_803 & 16'hf0f0;
  assign T_806 = T_801 | T_805;
  assign T_810 = T_806[15:2];
  assign GEN_31 = {{2'd0}, T_810};
  assign T_811 = GEN_31 & 16'h3333;
  assign T_812 = T_806[13:0];
  assign GEN_32 = {{2'd0}, T_812};
  assign T_813 = GEN_32 << 2;
  assign T_815 = T_813 & 16'hcccc;
  assign T_816 = T_811 | T_815;
  assign T_820 = T_816[15:1];
  assign GEN_33 = {{1'd0}, T_820};
  assign T_821 = GEN_33 & 16'h5555;
  assign T_822 = T_816[14:0];
  assign GEN_34 = {{1'd0}, T_822};
  assign T_823 = GEN_34 << 1;
  assign T_825 = T_823 & 16'haaaa;
  assign T_826 = T_821 | T_825;
  assign T_827 = T_784[17:16];
  assign T_828 = T_827[0];
  assign T_829 = T_827[1];
  assign T_830 = {T_828,T_829};
  assign T_831 = {T_826,T_830};
  assign T_832 = {T_783,T_831};
  assign T_833 = ~ T_832;
  assign T_834 = T_726 ? 50'h0 : T_833;
  assign T_835 = ~ T_834;
  assign T_836 = ~ T_835;
  assign T_837 = T_723 ? 50'h0 : T_836;
  assign T_838 = ~ T_837;
  assign T_839 = ~ T_838;
  assign T_840 = T_720 ? 50'h0 : T_839;
  assign T_841 = ~ T_840;
  assign T_842 = ~ T_841;
  assign T_843 = T_717 ? 50'h0 : T_842;
  assign T_844 = ~ T_843;
  assign T_846 = {T_844,4'hf};
  assign T_857 = T_730[3:0];
  assign T_858 = T_857[1:0];
  assign T_859 = T_858[0];
  assign T_860 = T_858[1];
  assign T_861 = {T_859,T_860};
  assign T_862 = T_857[3:2];
  assign T_863 = T_862[0];
  assign T_864 = T_862[1];
  assign T_865 = {T_863,T_864};
  assign T_866 = {T_861,T_865};
  assign T_868 = T_726 ? T_866 : 4'h0;
  assign T_870 = T_723 ? T_868 : 4'h0;
  assign T_872 = T_720 ? T_870 : 4'h0;
  assign T_874 = T_717 ? T_872 : 4'h0;
  assign T_875 = T_715 ? T_846 : {{50'd0}, T_874};
  assign T_877 = T_713 ? T_875 : 54'h0;
  assign T_879 = T_711 ? T_877 : 54'h0;
  assign T_880 = sigX3[55];
  assign GEN_35 = {{53'd0}, T_880};
  assign T_881 = T_879 | GEN_35;
  assign T_883 = {T_881,2'h3};
  assign roundMask = T_709 | T_883;
  assign T_884 = roundMask[55:1];
  assign T_885 = ~ T_884;
  assign GEN_36 = {{1'd0}, T_885};
  assign roundPosMask = GEN_36 & roundMask;
  assign GEN_37 = {{1'd0}, roundPosMask};
  assign T_886 = sigX3 & GEN_37;
  assign roundPosBit = T_886 != 57'h0;
  assign GEN_38 = {{2'd0}, T_884};
  assign T_889 = sigX3 & GEN_38;
  assign anyRoundExtra = T_889 != 57'h0;
  assign T_891 = ~ sigX3;
  assign T_893 = T_891 & GEN_38;
  assign allRoundExtra = T_893 == 57'h0;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign allRound = roundPosBit & allRoundExtra;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign T_896 = doIncrSig == 1'h0;
  assign T_897 = T_896 & roundingMode_nearest_even;
  assign T_898 = T_897 & roundPosBit;
  assign T_899 = T_898 & anyRoundExtra;
  assign T_902 = T_896 & roundDirectUp;
  assign T_903 = T_902 & anyRound;
  assign T_904 = T_899 | T_903;
  assign T_905 = doIncrSig & allRound;
  assign T_906 = T_904 | T_905;
  assign T_907 = doIncrSig & roundingMode_nearest_even;
  assign T_908 = T_907 & roundPosBit;
  assign T_909 = T_906 | T_908;
  assign T_910 = doIncrSig & roundDirectUp;
  assign roundUp = T_909 | T_910;
  assign T_914 = roundPosBit == 1'h0;
  assign T_915 = roundingMode_nearest_even & T_914;
  assign T_916 = T_915 & allRoundExtra;
  assign T_917 = roundingMode_nearest_even & roundPosBit;
  assign T_919 = anyRoundExtra == 1'h0;
  assign T_920 = T_917 & T_919;
  assign roundEven = doIncrSig ? T_916 : T_920;
  assign T_922 = allRound == 1'h0;
  assign roundInexact = doIncrSig ? T_922 : anyRound;
  assign GEN_40 = {{1'd0}, roundMask};
  assign T_923 = sigX3 | GEN_40;
  assign T_924 = T_923[56:2];
  assign T_926 = T_924 + 55'h1;
  assign T_927 = T_926[54:0];
  assign T_929 = roundUp == 1'h0;
  assign T_931 = roundEven == 1'h0;
  assign T_932 = T_929 & T_931;
  assign T_933 = ~ roundMask;
  assign GEN_41 = {{1'd0}, T_933};
  assign T_934 = sigX3 & GEN_41;
  assign T_935 = T_934[56:2];
  assign T_937 = T_932 ? T_935 : 55'h0;
  assign T_939 = roundUp ? T_927 : 55'h0;
  assign T_940 = T_937 | T_939;
  assign T_943 = T_927 & T_885;
  assign T_945 = roundEven ? T_943 : 55'h0;
  assign sigY3 = T_940 | T_945;
  assign T_946 = sigY3[54];
  assign T_948 = sExpX3 + 14'h1;
  assign T_949 = T_948[13:0];
  assign T_951 = T_946 ? T_949 : 14'h0;
  assign T_952 = sigY3[53];
  assign T_954 = T_952 ? sExpX3 : 14'h0;
  assign T_955 = T_951 | T_954;
  assign T_956 = sigY3[54:53];
  assign T_958 = T_956 == 2'h0;
  assign T_960 = sExpX3 - 14'h1;
  assign T_961 = T_960[13:0];
  assign T_963 = T_958 ? T_961 : 14'h0;
  assign sExpY = T_955 | T_963;
  assign expY = sExpY[11:0];
  assign T_964 = sigY3[51:0];
  assign T_965 = sigY3[52:1];
  assign fractY = sigX3Shift1 ? T_964 : T_965;
  assign T_966 = sExpY[12:10];
  assign overflowY = T_966 == 3'h3;
  assign T_969 = isZeroY == 1'h0;
  assign T_970 = sExpY[12];
  assign T_973 = expY < 12'h3ce;
  assign T_974 = T_970 | T_973;
  assign totalUnderflowY = T_969 & T_974;
  assign T_978 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign GEN_42 = {{2'd0}, T_978};
  assign T_979 = sExpX3_13 <= GEN_42;
  assign T_980 = T_705 | T_979;
  assign underflowY = roundInexact & T_980;
  assign T_981 = roundingMode_min & signY;
  assign T_983 = signY == 1'h0;
  assign T_984 = roundingMode_max & T_983;
  assign roundMagUp = T_981 | T_984;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign mulSpecial = isSpecialA | isSpecialB;
  assign addSpecial = mulSpecial | isSpecialC;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign T_986 = addSpecial == 1'h0;
  assign T_988 = notSpecial_addZeros == 1'h0;
  assign commonCase = T_986 & T_988;
  assign T_989 = isInfA & isZeroB;
  assign T_990 = isZeroA & isInfB;
  assign T_991 = T_989 | T_990;
  assign T_993 = isNaNA == 1'h0;
  assign T_995 = isNaNB == 1'h0;
  assign T_996 = T_993 & T_995;
  assign T_997 = isInfA | isInfB;
  assign T_998 = T_996 & T_997;
  assign T_999 = T_998 & isInfC;
  assign T_1000 = T_999 & doSubMags;
  assign notSigNaN_invalid = T_991 | T_1000;
  assign T_1001 = isSigNaNA | isSigNaNB;
  assign T_1002 = T_1001 | isSigNaNC;
  assign invalid = T_1002 | notSigNaN_invalid;
  assign overflow = commonCase & overflowY;
  assign underflow = commonCase & underflowY;
  assign T_1003 = commonCase & roundInexact;
  assign inexact = overflow | T_1003;
  assign T_1004 = notSpecial_addZeros | isZeroY;
  assign notSpecial_isZeroOut = T_1004 | totalUnderflowY;
  assign T_1005 = commonCase & totalUnderflowY;
  assign pegMinFiniteMagOut = T_1005 & roundMagUp;
  assign T_1007 = overflowY_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = overflow & T_1007;
  assign T_1009 = T_997 | isInfC;
  assign T_1010 = overflow & overflowY_roundMagUp;
  assign notNaN_isInfOut = T_1009 | T_1010;
  assign T_1011 = isNaNA | isNaNB;
  assign T_1012 = T_1011 | isNaNC;
  assign isNaNOut = T_1012 | notSigNaN_invalid;
  assign T_1015 = T_472 & io_fromPreMul_opSignC;
  assign T_1017 = isSpecialC == 1'h0;
  assign T_1018 = mulSpecial & T_1017;
  assign T_1019 = T_1018 & io_fromPreMul_signProd;
  assign T_1020 = T_1015 | T_1019;
  assign T_1022 = mulSpecial == 1'h0;
  assign T_1023 = T_1022 & isSpecialC;
  assign T_1024 = T_1023 & io_fromPreMul_opSignC;
  assign T_1025 = T_1020 | T_1024;
  assign T_1028 = T_1022 & notSpecial_addZeros;
  assign T_1029 = T_1028 & doSubMags;
  assign T_1030 = T_1029 & roundingMode_min;
  assign uncommonCaseSignOut = T_1025 | T_1030;
  assign T_1032 = isNaNOut == 1'h0;
  assign T_1033 = T_1032 & uncommonCaseSignOut;
  assign T_1034 = commonCase & signY;
  assign signOut = T_1033 | T_1034;
  assign T_1037 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign T_1038 = ~ T_1037;
  assign T_1039 = expY & T_1038;
  assign T_1043 = pegMinFiniteMagOut ? 12'hc31 : 12'h0;
  assign T_1044 = ~ T_1043;
  assign T_1045 = T_1039 & T_1044;
  assign T_1048 = pegMaxFiniteMagOut ? 12'h400 : 12'h0;
  assign T_1049 = ~ T_1048;
  assign T_1050 = T_1045 & T_1049;
  assign T_1053 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T_1054 = ~ T_1053;
  assign T_1055 = T_1050 & T_1054;
  assign T_1058 = pegMinFiniteMagOut ? 12'h3ce : 12'h0;
  assign T_1059 = T_1055 | T_1058;
  assign T_1062 = pegMaxFiniteMagOut ? 12'hbff : 12'h0;
  assign T_1063 = T_1059 | T_1062;
  assign T_1066 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign T_1067 = T_1063 | T_1066;
  assign T_1070 = isNaNOut ? 12'he00 : 12'h0;
  assign expOut = T_1067 | T_1070;
  assign T_1071 = totalUnderflowY & roundMagUp;
  assign T_1072 = T_1071 | isNaNOut;
  assign T_1076 = isNaNOut ? 52'h8000000000000 : 52'h0;
  assign T_1077 = T_1072 ? T_1076 : fractY;
  assign T_1081 = pegMaxFiniteMagOut ? 52'hfffffffffffff : 52'h0;
  assign fractOut = T_1077 | T_1081;
  assign T_1082 = {signOut,expOut};
  assign T_1083 = {T_1082,fractOut};
  assign T_1085 = {underflow,inexact};
  assign T_1086 = {invalid,1'h0};
  assign T_1087 = {T_1086,overflow};
  assign T_1088 = {T_1087,T_1085};
endmodule
module MulAddRecFN_1(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  mulAddRecFN_preMul_clk;
  wire  mulAddRecFN_preMul_reset;
  wire [1:0] mulAddRecFN_preMul_io_op;
  wire [64:0] mulAddRecFN_preMul_io_a;
  wire [64:0] mulAddRecFN_preMul_io_b;
  wire [64:0] mulAddRecFN_preMul_io_c;
  wire [1:0] mulAddRecFN_preMul_io_roundingMode;
  wire [52:0] mulAddRecFN_preMul_io_mulAddA;
  wire [52:0] mulAddRecFN_preMul_io_mulAddB;
  wire [105:0] mulAddRecFN_preMul_io_mulAddC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_preMul_io_toPostMul_signProd;
  wire  mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire  mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire  mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire [7:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire  mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire [54:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire [13:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire [1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire  mulAddRecFN_postMul_clk;
  wire  mulAddRecFN_postMul_reset;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpA;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpB;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_postMul_io_fromPreMul_signProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_isZeroProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_opSignC;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isCDominant;
  wire  mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0;
  wire [7:0] mulAddRecFN_postMul_io_fromPreMul_CAlignDist;
  wire  mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC;
  wire [54:0] mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC;
  wire [13:0] mulAddRecFN_postMul_io_fromPreMul_sExpSum;
  wire [1:0] mulAddRecFN_postMul_io_fromPreMul_roundingMode;
  wire [106:0] mulAddRecFN_postMul_io_mulAddResult;
  wire [64:0] mulAddRecFN_postMul_io_out;
  wire [4:0] mulAddRecFN_postMul_io_exceptionFlags;
  wire [105:0] T_7;
  wire [106:0] T_9;
  wire [106:0] GEN_0;
  wire [107:0] T_10;
  wire [106:0] T_11;
  MulAddRecFN_preMul_1 mulAddRecFN_preMul (
    .clk(mulAddRecFN_preMul_clk),
    .reset(mulAddRecFN_preMul_reset),
    .io_op(mulAddRecFN_preMul_io_op),
    .io_a(mulAddRecFN_preMul_io_a),
    .io_b(mulAddRecFN_preMul_io_b),
    .io_c(mulAddRecFN_preMul_io_c),
    .io_roundingMode(mulAddRecFN_preMul_io_roundingMode),
    .io_mulAddA(mulAddRecFN_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFN_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFN_preMul_io_mulAddC),
    .io_toPostMul_highExpA(mulAddRecFN_preMul_io_toPostMul_highExpA),
    .io_toPostMul_isNaN_isQuietNaNA(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA),
    .io_toPostMul_highExpB(mulAddRecFN_preMul_io_toPostMul_highExpB),
    .io_toPostMul_isNaN_isQuietNaNB(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB),
    .io_toPostMul_signProd(mulAddRecFN_preMul_io_toPostMul_signProd),
    .io_toPostMul_isZeroProd(mulAddRecFN_preMul_io_toPostMul_isZeroProd),
    .io_toPostMul_opSignC(mulAddRecFN_preMul_io_toPostMul_opSignC),
    .io_toPostMul_highExpC(mulAddRecFN_preMul_io_toPostMul_highExpC),
    .io_toPostMul_isNaN_isQuietNaNC(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC),
    .io_toPostMul_isCDominant(mulAddRecFN_preMul_io_toPostMul_isCDominant),
    .io_toPostMul_CAlignDist_0(mulAddRecFN_preMul_io_toPostMul_CAlignDist_0),
    .io_toPostMul_CAlignDist(mulAddRecFN_preMul_io_toPostMul_CAlignDist),
    .io_toPostMul_bit0AlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC),
    .io_toPostMul_highAlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC),
    .io_toPostMul_sExpSum(mulAddRecFN_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_roundingMode(mulAddRecFN_preMul_io_toPostMul_roundingMode)
  );
  MulAddRecFN_postMul_1 mulAddRecFN_postMul (
    .clk(mulAddRecFN_postMul_clk),
    .reset(mulAddRecFN_postMul_reset),
    .io_fromPreMul_highExpA(mulAddRecFN_postMul_io_fromPreMul_highExpA),
    .io_fromPreMul_isNaN_isQuietNaNA(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA),
    .io_fromPreMul_highExpB(mulAddRecFN_postMul_io_fromPreMul_highExpB),
    .io_fromPreMul_isNaN_isQuietNaNB(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB),
    .io_fromPreMul_signProd(mulAddRecFN_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isZeroProd(mulAddRecFN_postMul_io_fromPreMul_isZeroProd),
    .io_fromPreMul_opSignC(mulAddRecFN_postMul_io_fromPreMul_opSignC),
    .io_fromPreMul_highExpC(mulAddRecFN_postMul_io_fromPreMul_highExpC),
    .io_fromPreMul_isNaN_isQuietNaNC(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC),
    .io_fromPreMul_isCDominant(mulAddRecFN_postMul_io_fromPreMul_isCDominant),
    .io_fromPreMul_CAlignDist_0(mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0),
    .io_fromPreMul_CAlignDist(mulAddRecFN_postMul_io_fromPreMul_CAlignDist),
    .io_fromPreMul_bit0AlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC),
    .io_fromPreMul_highAlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC),
    .io_fromPreMul_sExpSum(mulAddRecFN_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_roundingMode(mulAddRecFN_postMul_io_fromPreMul_roundingMode),
    .io_mulAddResult(mulAddRecFN_postMul_io_mulAddResult),
    .io_out(mulAddRecFN_postMul_io_out),
    .io_exceptionFlags(mulAddRecFN_postMul_io_exceptionFlags)
  );
  assign io_out = mulAddRecFN_postMul_io_out;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign mulAddRecFN_preMul_clk = clk;
  assign mulAddRecFN_preMul_reset = reset;
  assign mulAddRecFN_preMul_io_op = io_op;
  assign mulAddRecFN_preMul_io_a = io_a;
  assign mulAddRecFN_preMul_io_b = io_b;
  assign mulAddRecFN_preMul_io_c = io_c;
  assign mulAddRecFN_preMul_io_roundingMode = io_roundingMode;
  assign mulAddRecFN_postMul_clk = clk;
  assign mulAddRecFN_postMul_reset = reset;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpA = mulAddRecFN_preMul_io_toPostMul_highExpA;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpB = mulAddRecFN_preMul_io_toPostMul_highExpB;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  assign mulAddRecFN_postMul_io_fromPreMul_signProd = mulAddRecFN_preMul_io_toPostMul_signProd;
  assign mulAddRecFN_postMul_io_fromPreMul_isZeroProd = mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  assign mulAddRecFN_postMul_io_fromPreMul_opSignC = mulAddRecFN_preMul_io_toPostMul_opSignC;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpC = mulAddRecFN_preMul_io_toPostMul_highExpC;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  assign mulAddRecFN_postMul_io_fromPreMul_isCDominant = mulAddRecFN_preMul_io_toPostMul_isCDominant;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0 = mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist = mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  assign mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_sExpSum = mulAddRecFN_preMul_io_toPostMul_sExpSum;
  assign mulAddRecFN_postMul_io_fromPreMul_roundingMode = mulAddRecFN_preMul_io_toPostMul_roundingMode;
  assign mulAddRecFN_postMul_io_mulAddResult = T_11;
  assign T_7 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign T_9 = {1'h0,mulAddRecFN_preMul_io_mulAddC};
  assign GEN_0 = {{1'd0}, T_7};
  assign T_10 = GEN_0 + T_9;
  assign T_11 = T_10[106:0];
endmodule
module FPUFMAPipe_1(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [64:0] GEN_28;
  wire [64:0] zero;
  reg  valid;
  reg [31:0] GEN_29;
  reg [4:0] in_cmd;
  reg [31:0] GEN_30;
  reg  in_ldst;
  reg [31:0] GEN_31;
  reg  in_wen;
  reg [31:0] GEN_32;
  reg  in_ren1;
  reg [31:0] GEN_33;
  reg  in_ren2;
  reg [31:0] GEN_34;
  reg  in_ren3;
  reg [31:0] GEN_35;
  reg  in_swap12;
  reg [31:0] GEN_36;
  reg  in_swap23;
  reg [31:0] GEN_37;
  reg  in_single;
  reg [31:0] GEN_38;
  reg  in_fromint;
  reg [31:0] GEN_39;
  reg  in_toint;
  reg [31:0] GEN_40;
  reg  in_fastpipe;
  reg [31:0] GEN_41;
  reg  in_fma;
  reg [31:0] GEN_42;
  reg  in_div;
  reg [31:0] GEN_43;
  reg  in_sqrt;
  reg [31:0] GEN_44;
  reg  in_round;
  reg [31:0] GEN_45;
  reg  in_wflags;
  reg [31:0] GEN_46;
  reg [2:0] in_rm;
  reg [31:0] GEN_47;
  reg [1:0] in_typ;
  reg [31:0] GEN_48;
  reg [64:0] in_in1;
  reg [95:0] GEN_49;
  reg [64:0] in_in2;
  reg [95:0] GEN_50;
  reg [64:0] in_in3;
  reg [95:0] GEN_51;
  wire  T_179;
  wire  T_180;
  wire  T_181;
  wire  T_182;
  wire [1:0] T_183;
  wire [64:0] GEN_0;
  wire  T_186;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  fma_clk;
  wire  fma_reset;
  wire [1:0] fma_io_op;
  wire [64:0] fma_io_a;
  wire [64:0] fma_io_b;
  wire [64:0] fma_io_c;
  wire [1:0] fma_io_roundingMode;
  wire [64:0] fma_io_out;
  wire [4:0] fma_io_exceptionFlags;
  wire [64:0] res_data;
  wire [4:0] res_exc;
  wire [65:0] T_193;
  reg  T_196;
  reg [31:0] GEN_52;
  reg [64:0] T_197_data;
  reg [95:0] GEN_53;
  reg [4:0] T_197_exc;
  reg [31:0] GEN_54;
  wire [64:0] GEN_24;
  wire [4:0] GEN_25;
  reg  T_202;
  reg [31:0] GEN_55;
  reg [64:0] T_203_data;
  reg [95:0] GEN_56;
  reg [4:0] T_203_exc;
  reg [31:0] GEN_57;
  wire [64:0] GEN_26;
  wire [4:0] GEN_27;
  wire  T_214_valid;
  wire [64:0] T_214_bits_data;
  wire [4:0] T_214_bits_exc;
  MulAddRecFN_1 fma (
    .clk(fma_clk),
    .reset(fma_reset),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags)
  );
  assign io_out_valid = T_214_valid;
  assign io_out_bits_data = T_214_bits_data;
  assign io_out_bits_exc = T_214_bits_exc;
  assign T_131 = io_in_bits_in1[64];
  assign T_132 = io_in_bits_in2[64];
  assign T_133 = T_131 ^ T_132;
  assign GEN_28 = {{64'd0}, T_133};
  assign zero = GEN_28 << 64;
  assign T_179 = io_in_bits_cmd[1];
  assign T_180 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T_181 = T_179 & T_180;
  assign T_182 = io_in_bits_cmd[0];
  assign T_183 = {T_181,T_182};
  assign GEN_0 = io_in_bits_swap23 ? 65'h8000000000000000 : io_in_bits_in2;
  assign T_186 = T_180 == 1'h0;
  assign GEN_1 = T_186 ? zero : io_in_bits_in3;
  assign GEN_2 = io_in_valid ? {{3'd0}, T_183} : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_0 : in_in2;
  assign GEN_23 = io_in_valid ? GEN_1 : in_in3;
  assign fma_clk = clk;
  assign fma_reset = reset;
  assign fma_io_op = in_cmd[1:0];
  assign fma_io_a = in_in1;
  assign fma_io_b = in_in2;
  assign fma_io_c = in_in3;
  assign fma_io_roundingMode = in_rm[1:0];
  assign res_data = T_193[64:0];
  assign res_exc = fma_io_exceptionFlags;
  assign T_193 = {1'h0,fma_io_out};
  assign GEN_24 = valid ? res_data : T_197_data;
  assign GEN_25 = valid ? res_exc : T_197_exc;
  assign GEN_26 = T_196 ? T_197_data : T_203_data;
  assign GEN_27 = T_196 ? T_197_exc : T_203_exc;
  assign T_214_valid = T_202;
  assign T_214_bits_data = T_203_data;
  assign T_214_bits_exc = T_203_exc;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  valid = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  in_cmd = GEN_30[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  in_ldst = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  in_wen = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  in_ren1 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_34 = {1{$random}};
  in_ren2 = GEN_34[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  in_ren3 = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  in_swap12 = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_37 = {1{$random}};
  in_swap23 = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_38 = {1{$random}};
  in_single = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  in_fromint = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  in_toint = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  in_fastpipe = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  in_fma = GEN_42[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  in_div = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  in_sqrt = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  in_round = GEN_45[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  in_wflags = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  in_rm = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  in_typ = GEN_48[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {3{$random}};
  in_in1 = GEN_49[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {3{$random}};
  in_in2 = GEN_50[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {3{$random}};
  in_in3 = GEN_51[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  T_196 = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_53 = {3{$random}};
  T_197_data = GEN_53[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_54 = {1{$random}};
  T_197_exc = GEN_54[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  T_202 = GEN_55[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {3{$random}};
  T_203_data = GEN_56[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  T_203_exc = GEN_57[4:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_cmd <= {{3'd0}, T_183};
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ldst <= io_in_bits_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wen <= io_in_bits_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren1 <= io_in_bits_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren2 <= io_in_bits_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_ren3 <= io_in_bits_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap12 <= io_in_bits_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_swap23 <= io_in_bits_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_single <= io_in_bits_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fromint <= io_in_bits_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_toint <= io_in_bits_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fastpipe <= io_in_bits_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_fma <= io_in_bits_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_div <= io_in_bits_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_sqrt <= io_in_bits_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_round <= io_in_bits_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_wflags <= io_in_bits_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_rm <= io_in_bits_rm;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_typ <= io_in_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        in_in1 <= io_in_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(io_in_bits_swap23) begin
          in_in2 <= 65'h8000000000000000;
        end else begin
          in_in2 <= io_in_bits_in2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_in_valid) begin
        if(T_186) begin
          in_in3 <= zero;
        end else begin
          in_in3 <= io_in_bits_in3;
        end
      end
    end
    if(reset) begin
      T_196 <= 1'h0;
    end else begin
      T_196 <= valid;
    end
    if(1'h0) begin
    end else begin
      if(valid) begin
        T_197_data <= res_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(valid) begin
        T_197_exc <= res_exc;
      end
    end
    if(reset) begin
      T_202 <= 1'h0;
    end else begin
      T_202 <= T_196;
    end
    if(1'h0) begin
    end else begin
      if(T_196) begin
        T_203_data <= T_197_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_196) begin
        T_203_exc <= T_197_exc;
      end
    end
  end
endmodule
module DivSqrtRecF64_mulAddZ31(
  input   clk,
  input   reset,
  output  io_inReady_div,
  output  io_inReady_sqrt,
  input   io_inValid,
  input   io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [1:0] io_roundingMode,
  output  io_outValid_div,
  output  io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [3:0] io_usingMulAdd,
  output  io_latchMulAddA_0,
  output [53:0] io_mulAddA_0,
  output  io_latchMulAddB_0,
  output [53:0] io_mulAddB_0,
  output [104:0] io_mulAddC_2,
  input  [104:0] io_mulAddResult_3
);
  reg  valid_PA;
  reg [31:0] GEN_115;
  reg  sqrtOp_PA;
  reg [31:0] GEN_119;
  reg  sign_PA;
  reg [31:0] GEN_120;
  reg [2:0] specialCodeB_PA;
  reg [31:0] GEN_121;
  reg  fractB_51_PA;
  reg [31:0] GEN_122;
  reg [1:0] roundingMode_PA;
  reg [31:0] GEN_123;
  reg [2:0] specialCodeA_PA;
  reg [31:0] GEN_124;
  reg  fractA_51_PA;
  reg [31:0] GEN_125;
  reg [13:0] exp_PA;
  reg [31:0] GEN_126;
  reg [50:0] fractB_other_PA;
  reg [63:0] GEN_127;
  reg [50:0] fractA_other_PA;
  reg [63:0] GEN_128;
  reg  valid_PB;
  reg [31:0] GEN_129;
  reg  sqrtOp_PB;
  reg [31:0] GEN_130;
  reg  sign_PB;
  reg [31:0] GEN_131;
  reg [2:0] specialCodeA_PB;
  reg [31:0] GEN_132;
  reg  fractA_51_PB;
  reg [31:0] GEN_133;
  reg [2:0] specialCodeB_PB;
  reg [31:0] GEN_134;
  reg  fractB_51_PB;
  reg [31:0] GEN_135;
  reg [1:0] roundingMode_PB;
  reg [31:0] GEN_136;
  reg [13:0] exp_PB;
  reg [31:0] GEN_137;
  reg  fractA_0_PB;
  reg [31:0] GEN_138;
  reg [50:0] fractB_other_PB;
  reg [63:0] GEN_139;
  reg  valid_PC;
  reg [31:0] GEN_140;
  reg  sqrtOp_PC;
  reg [31:0] GEN_141;
  reg  sign_PC;
  reg [31:0] GEN_142;
  reg [2:0] specialCodeA_PC;
  reg [31:0] GEN_143;
  reg  fractA_51_PC;
  reg [31:0] GEN_144;
  reg [2:0] specialCodeB_PC;
  reg [31:0] GEN_145;
  reg  fractB_51_PC;
  reg [31:0] GEN_146;
  reg [1:0] roundingMode_PC;
  reg [31:0] GEN_147;
  reg [13:0] exp_PC;
  reg [31:0] GEN_148;
  reg  fractA_0_PC;
  reg [31:0] GEN_149;
  reg [50:0] fractB_other_PC;
  reg [63:0] GEN_150;
  reg [2:0] cycleNum_A;
  reg [31:0] GEN_151;
  reg [3:0] cycleNum_B;
  reg [31:0] GEN_152;
  reg [2:0] cycleNum_C;
  reg [31:0] GEN_153;
  reg [2:0] cycleNum_E;
  reg [31:0] GEN_154;
  reg [8:0] fractR0_A;
  reg [31:0] GEN_155;
  reg [9:0] hiSqrR0_A_sqrt;
  reg [31:0] GEN_156;
  reg [20:0] partNegSigma0_A;
  reg [31:0] GEN_157;
  reg [8:0] nextMulAdd9A_A;
  reg [31:0] GEN_158;
  reg [8:0] nextMulAdd9B_A;
  reg [31:0] GEN_159;
  reg [16:0] ER1_B_sqrt;
  reg [31:0] GEN_160;
  reg [31:0] ESqrR1_B_sqrt;
  reg [31:0] GEN_161;
  reg [57:0] sigX1_B;
  reg [63:0] GEN_162;
  reg [32:0] sqrSigma1_C;
  reg [63:0] GEN_163;
  reg [57:0] sigXN_C;
  reg [63:0] GEN_164;
  reg [30:0] u_C_sqrt;
  reg [31:0] GEN_165;
  reg  E_E_div;
  reg [31:0] GEN_166;
  reg [52:0] sigT_E;
  reg [63:0] GEN_167;
  reg  extraT_E;
  reg [31:0] GEN_168;
  reg  isNegRemT_E;
  reg [31:0] GEN_169;
  reg  trueEqX_E1;
  reg [31:0] GEN_170;
  wire  ready_PA;
  wire  ready_PB;
  wire  ready_PC;
  wire  leaving_PA;
  wire  leaving_PB;
  wire  leaving_PC;
  wire  cyc_B10_sqrt;
  wire  cyc_B9_sqrt;
  wire  cyc_B8_sqrt;
  wire  cyc_B7_sqrt;
  wire  cyc_B6;
  wire  cyc_B5;
  wire  cyc_B4;
  wire  cyc_B3;
  wire  cyc_B2;
  wire  cyc_B1;
  wire  cyc_B6_div;
  wire  cyc_B5_div;
  wire  cyc_B4_div;
  wire  cyc_B3_div;
  wire  cyc_B2_div;
  wire  cyc_B1_div;
  wire  cyc_B6_sqrt;
  wire  cyc_B5_sqrt;
  wire  cyc_B4_sqrt;
  wire  cyc_B3_sqrt;
  wire  cyc_B2_sqrt;
  wire  cyc_B1_sqrt;
  wire  cyc_C5;
  wire  cyc_C4;
  wire  valid_normalCase_leaving_PB;
  wire  cyc_C2;
  wire  cyc_C1;
  wire  cyc_E4;
  wire  cyc_E3;
  wire  cyc_E2;
  wire  cyc_E1;
  wire [45:0] zSigma1_B4;
  wire [57:0] sigXNU_B3_CX;
  wire [53:0] zComplSigT_C1_sqrt;
  wire [53:0] zComplSigT_C1;
  wire  T_113;
  wire  T_114;
  wire  T_116;
  wire  T_117;
  wire  T_119;
  wire  T_120;
  wire  T_122;
  wire  T_123;
  wire  T_125;
  wire  T_126;
  wire  T_128;
  wire  T_129;
  wire  T_131;
  wire  T_132;
  wire  T_134;
  wire  T_135;
  wire  T_137;
  wire  T_138;
  wire  T_141;
  wire  T_144;
  wire  T_147;
  wire  T_149;
  wire  T_150;
  wire  T_153;
  wire  T_154;
  wire  T_156;
  wire  cyc_S_div;
  wire  T_157;
  wire  cyc_S_sqrt;
  wire  cyc_S;
  wire  signA_S;
  wire [11:0] expA_S;
  wire [51:0] fractA_S;
  wire [2:0] specialCodeA_S;
  wire  isZeroA_S;
  wire [1:0] T_159;
  wire  isSpecialA_S;
  wire  signB_S;
  wire [11:0] expB_S;
  wire [51:0] fractB_S;
  wire [2:0] specialCodeB_S;
  wire  isZeroB_S;
  wire [1:0] T_162;
  wire  isSpecialB_S;
  wire  T_164;
  wire  sign_S;
  wire  T_166;
  wire  T_168;
  wire  T_169;
  wire  T_171;
  wire  T_172;
  wire  T_174;
  wire  normalCase_S_div;
  wire  T_179;
  wire  T_181;
  wire  normalCase_S_sqrt;
  wire  normalCase_S;
  wire  entering_PA_normalCase_div;
  wire  entering_PA_normalCase_sqrt;
  wire  entering_PA_normalCase;
  wire  T_183;
  wire  T_184;
  wire  T_185;
  wire  entering_PA;
  wire  T_187;
  wire  T_188;
  wire  T_190;
  wire  T_191;
  wire  T_193;
  wire  T_195;
  wire  T_196;
  wire  T_197;
  wire  entering_PB_S;
  wire  T_206;
  wire  entering_PC_S;
  wire  T_207;
  wire  GEN_0;
  wire  T_208;
  wire  GEN_1;
  wire  GEN_2;
  wire [2:0] GEN_3;
  wire  GEN_4;
  wire [1:0] GEN_5;
  wire  T_211;
  wire  T_212;
  wire [2:0] GEN_6;
  wire  GEN_7;
  wire  T_213;
  wire [2:0] T_217;
  wire [10:0] T_218;
  wire [10:0] T_219;
  wire [13:0] T_220;
  wire [13:0] GEN_53;
  wire [14:0] T_221;
  wire [13:0] T_222;
  wire [13:0] T_223;
  wire [50:0] T_224;
  wire [13:0] GEN_8;
  wire [50:0] GEN_9;
  wire [50:0] T_225;
  wire [50:0] GEN_10;
  wire  isZeroA_PA;
  wire [1:0] T_227;
  wire  isSpecialA_PA;
  wire [1:0] T_230;
  wire [52:0] sigA_PA;
  wire  isZeroB_PA;
  wire [1:0] T_232;
  wire  isSpecialB_PA;
  wire [1:0] T_235;
  wire [52:0] sigB_PA;
  wire  T_237;
  wire  T_239;
  wire  T_240;
  wire  T_242;
  wire  T_243;
  wire  T_245;
  wire  T_248;
  wire  T_250;
  wire  T_251;
  wire  T_254;
  wire  normalCase_PA;
  wire  valid_normalCase_leaving_PA;
  wire  valid_leaving_PA;
  wire  T_255;
  wire  T_258;
  wire  T_259;
  wire  entering_PB_normalCase;
  wire  entering_PB;
  wire  T_260;
  wire  GEN_11;
  wire  T_261;
  wire  T_262;
  wire [2:0] T_263;
  wire  T_265;
  wire [2:0] T_266;
  wire  T_268;
  wire [1:0] T_269;
  wire  GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire  GEN_15;
  wire [2:0] GEN_16;
  wire  GEN_17;
  wire [1:0] GEN_18;
  wire  T_270;
  wire [13:0] GEN_19;
  wire  GEN_20;
  wire [50:0] GEN_21;
  wire  isZeroA_PB;
  wire [1:0] T_272;
  wire  isSpecialA_PB;
  wire  isZeroB_PB;
  wire [1:0] T_275;
  wire  isSpecialB_PB;
  wire  T_278;
  wire  T_280;
  wire  T_281;
  wire  T_283;
  wire  T_284;
  wire  T_286;
  wire  T_289;
  wire  T_291;
  wire  T_292;
  wire  T_295;
  wire  normalCase_PB;
  wire  valid_leaving_PB;
  wire  T_296;
  wire  T_299;
  wire  T_300;
  wire  entering_PC_normalCase;
  wire  entering_PC;
  wire  T_301;
  wire  GEN_22;
  wire  T_302;
  wire  T_303;
  wire [2:0] T_304;
  wire  T_306;
  wire [2:0] T_307;
  wire  T_309;
  wire [1:0] T_310;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [1:0] GEN_29;
  wire [13:0] GEN_30;
  wire  GEN_31;
  wire [50:0] GEN_32;
  wire  isZeroA_PC;
  wire [1:0] T_312;
  wire  isSpecialA_PC;
  wire  T_314;
  wire  T_316;
  wire  isInfA_PC;
  wire  isNaNA_PC;
  wire  T_319;
  wire  isSigNaNA_PC;
  wire  isZeroB_PC;
  wire [1:0] T_321;
  wire  isSpecialB_PC;
  wire  T_323;
  wire  T_325;
  wire  isInfB_PC;
  wire  isNaNB_PC;
  wire  T_328;
  wire  isSigNaNB_PC;
  wire [1:0] T_330;
  wire [52:0] sigB_PC;
  wire  T_332;
  wire  T_334;
  wire  T_335;
  wire  T_337;
  wire  T_338;
  wire  T_340;
  wire  T_343;
  wire  T_345;
  wire  T_346;
  wire  T_349;
  wire  normalCase_PC;
  wire [14:0] T_351;
  wire [13:0] expP2_PC;
  wire  T_352;
  wire [12:0] T_353;
  wire [13:0] T_355;
  wire [12:0] T_356;
  wire [13:0] T_358;
  wire [13:0] expP1_PC;
  wire  roundingMode_near_even_PC;
  wire  roundingMode_min_PC;
  wire  roundingMode_max_PC;
  wire  roundMagUp_PC;
  wire  overflowY_roundMagUp_PC;
  wire  T_360;
  wire  T_362;
  wire  roundMagDown_PC;
  wire  T_364;
  wire  valid_leaving_PC;
  wire  T_365;
  wire  T_367;
  wire  T_368;
  wire  T_370;
  wire  T_371;
  wire  T_372;
  wire  T_374;
  wire  T_375;
  wire [1:0] T_378;
  wire [2:0] T_381;
  wire [2:0] GEN_54;
  wire [2:0] T_382;
  wire  T_384;
  wire [3:0] T_386;
  wire [2:0] T_387;
  wire [2:0] T_389;
  wire [2:0] T_390;
  wire [2:0] GEN_33;
  wire  cyc_A6_sqrt;
  wire  cyc_A5_sqrt;
  wire  cyc_A4_sqrt;
  wire  cyc_A4;
  wire  cyc_A3;
  wire  cyc_A2;
  wire  cyc_A1;
  wire  T_398;
  wire  cyc_A3_div;
  wire  cyc_A2_div;
  wire  cyc_A1_div;
  wire  cyc_A3_sqrt;
  wire  cyc_A1_sqrt;
  wire  T_404;
  wire  T_405;
  wire [3:0] T_408;
  wire [4:0] T_410;
  wire [3:0] T_411;
  wire [3:0] T_412;
  wire [3:0] GEN_34;
  wire  T_414;
  wire  T_416;
  wire  T_418;
  wire  T_420;
  wire  T_422;
  wire  T_424;
  wire  T_426;
  wire  T_428;
  wire  T_430;
  wire  T_432;
  wire  T_433;
  wire  T_436;
  wire  T_437;
  wire  T_440;
  wire  T_441;
  wire  T_444;
  wire  T_446;
  wire  T_447;
  wire  T_450;
  wire  T_453;
  wire  T_454;
  wire  T_455;
  wire  T_456;
  wire  T_457;
  wire  T_458;
  wire  T_459;
  wire  T_460;
  wire  T_461;
  wire  T_462;
  wire  T_464;
  wire  T_465;
  wire [2:0] T_468;
  wire [3:0] T_470;
  wire [2:0] T_471;
  wire [2:0] T_472;
  wire [2:0] GEN_35;
  wire  cyc_C6_sqrt;
  wire  T_475;
  wire  T_477;
  wire  T_479;
  wire  T_481;
  wire  T_483;
  wire  cyc_C5_div;
  wire  cyc_C4_div;
  wire  cyc_C1_div;
  wire  cyc_C5_sqrt;
  wire  cyc_C4_sqrt;
  wire  cyc_C3_sqrt;
  wire  cyc_C1_sqrt;
  wire  T_495;
  wire  T_496;
  wire [3:0] T_499;
  wire [2:0] T_500;
  wire [2:0] T_501;
  wire [2:0] GEN_36;
  wire  T_503;
  wire  T_505;
  wire  T_507;
  wire  T_509;
  wire  cyc_E3_div;
  wire  cyc_E3_sqrt;
  wire [51:0] zFractB_A4_div;
  wire [2:0] T_519;
  wire  T_521;
  wire  zLinPiece_0_A4_div;
  wire  T_524;
  wire  zLinPiece_1_A4_div;
  wire  T_527;
  wire  zLinPiece_2_A4_div;
  wire  T_530;
  wire  zLinPiece_3_A4_div;
  wire  T_533;
  wire  zLinPiece_4_A4_div;
  wire  T_536;
  wire  zLinPiece_5_A4_div;
  wire  T_539;
  wire  zLinPiece_6_A4_div;
  wire  T_542;
  wire  zLinPiece_7_A4_div;
  wire [8:0] T_545;
  wire [8:0] T_548;
  wire [8:0] T_549;
  wire [8:0] T_552;
  wire [8:0] T_553;
  wire [8:0] T_556;
  wire [8:0] T_557;
  wire [8:0] T_560;
  wire [8:0] T_561;
  wire [8:0] T_564;
  wire [8:0] T_565;
  wire [8:0] T_568;
  wire [8:0] T_569;
  wire [8:0] T_572;
  wire [8:0] zK1_A4_div;
  wire [11:0] T_576;
  wire [11:0] T_580;
  wire [11:0] T_581;
  wire [11:0] T_585;
  wire [11:0] T_586;
  wire [11:0] T_590;
  wire [11:0] T_591;
  wire [11:0] T_595;
  wire [11:0] T_596;
  wire [11:0] T_600;
  wire [11:0] T_601;
  wire [11:0] T_605;
  wire [11:0] T_606;
  wire [11:0] T_610;
  wire [11:0] zComplFractK0_A4_div;
  wire [51:0] zFractB_A7_sqrt;
  wire  T_612;
  wire  T_614;
  wire  T_615;
  wire  T_618;
  wire  zQuadPiece_0_A7_sqrt;
  wire  zQuadPiece_1_A7_sqrt;
  wire  T_625;
  wire  zQuadPiece_2_A7_sqrt;
  wire  zQuadPiece_3_A7_sqrt;
  wire [8:0] T_634;
  wire [8:0] T_637;
  wire [8:0] T_638;
  wire [8:0] T_641;
  wire [8:0] T_642;
  wire [8:0] T_645;
  wire [8:0] zK2_A7_sqrt;
  wire [9:0] T_649;
  wire [9:0] T_653;
  wire [9:0] T_654;
  wire [9:0] T_658;
  wire [9:0] T_659;
  wire [9:0] T_663;
  wire [9:0] zComplK1_A7_sqrt;
  wire  T_664;
  wire  T_666;
  wire  T_667;
  wire  T_668;
  wire  T_670;
  wire  zQuadPiece_0_A6_sqrt;
  wire  zQuadPiece_1_A6_sqrt;
  wire  T_677;
  wire  zQuadPiece_2_A6_sqrt;
  wire  zQuadPiece_3_A6_sqrt;
  wire [12:0] T_687;
  wire [12:0] T_691;
  wire [12:0] T_692;
  wire [12:0] T_696;
  wire [12:0] T_697;
  wire [12:0] T_701;
  wire [12:0] zComplFractK0_A6_sqrt;
  wire [8:0] T_702;
  wire [8:0] T_703;
  wire  T_705;
  wire [8:0] T_707;
  wire [8:0] mulAdd9A_A;
  wire [8:0] T_708;
  wire [8:0] T_709;
  wire [8:0] T_713;
  wire [8:0] mulAdd9B_A;
  wire [9:0] T_717;
  wire [19:0] T_718;
  wire [5:0] T_722;
  wire [13:0] T_723;
  wire [19:0] T_724;
  wire [19:0] T_725;
  wire [7:0] T_729;
  wire [12:0] T_730;
  wire [20:0] T_731;
  wire [20:0] GEN_55;
  wire [20:0] T_732;
  wire [18:0] GEN_56;
  wire [18:0] T_734;
  wire [19:0] GEN_57;
  wire [20:0] T_735;
  wire [19:0] T_736;
  wire [19:0] T_738;
  wire [20:0] GEN_58;
  wire [20:0] T_739;
  wire  T_740;
  wire  T_742;
  wire  T_743;
  wire [10:0] T_746;
  wire [20:0] GEN_59;
  wire [20:0] T_747;
  wire  T_749;
  wire  T_750;
  wire [20:0] T_751;
  wire [21:0] T_753;
  wire [20:0] T_754;
  wire [20:0] T_756;
  wire [20:0] T_757;
  wire  T_758;
  wire [20:0] T_760;
  wire [20:0] T_761;
  wire [24:0] GEN_60;
  wire [24:0] T_762;
  wire [24:0] T_764;
  wire [24:0] GEN_61;
  wire [24:0] T_765;
  wire [23:0] GEN_62;
  wire [23:0] T_766;
  wire [23:0] T_768;
  wire [24:0] GEN_63;
  wire [24:0] mulAdd9C_A;
  wire [17:0] T_769;
  wire [17:0] T_771;
  wire [18:0] T_772;
  wire [18:0] GEN_64;
  wire [19:0] T_773;
  wire [18:0] loMulAdd9Out_A;
  wire  T_774;
  wire [6:0] T_775;
  wire [7:0] T_777;
  wire [6:0] T_778;
  wire [6:0] T_780;
  wire [17:0] T_781;
  wire [24:0] mulAdd9Out_A;
  wire  T_782;
  wire  T_783;
  wire [24:0] T_784;
  wire [14:0] T_785;
  wire [14:0] T_787;
  wire [8:0] zFractR0_A6_sqrt;
  wire [25:0] GEN_65;
  wire [25:0] T_789;
  wire [25:0] sqrR0_A5_sqrt;
  wire  T_790;
  wire  T_791;
  wire [13:0] T_793;
  wire [13:0] T_795;
  wire [8:0] zFractR0_A4_div;
  wire  T_796;
  wire  T_797;
  wire [22:0] T_799;
  wire [22:0] T_801;
  wire [8:0] zSigma0_A2;
  wire [14:0] T_802;
  wire [15:0] T_803;
  wire [15:0] T_804;
  wire [14:0] fractR1_A1;
  wire [15:0] r1_A1;
  wire [16:0] GEN_66;
  wire [16:0] T_807;
  wire [16:0] ER1_A1_sqrt;
  wire  T_808;
  wire [8:0] T_809;
  wire [8:0] GEN_37;
  wire [15:0] T_810;
  wire [15:0] GEN_38;
  wire  T_811;
  wire [24:0] T_813;
  wire [20:0] T_814;
  wire [20:0] GEN_39;
  wire  T_815;
  wire  T_816;
  wire  T_817;
  wire  T_818;
  wire  T_819;
  wire [13:0] T_823;
  wire [13:0] GEN_67;
  wire [13:0] T_824;
  wire [8:0] T_825;
  wire [8:0] T_827;
  wire [13:0] GEN_68;
  wire [13:0] T_828;
  wire [8:0] T_829;
  wire [13:0] GEN_69;
  wire [13:0] T_830;
  wire  T_831;
  wire [8:0] T_832;
  wire [8:0] T_834;
  wire [13:0] GEN_70;
  wire [13:0] T_835;
  wire [13:0] GEN_71;
  wire [13:0] T_836;
  wire [13:0] GEN_40;
  wire  T_840;
  wire [8:0] T_842;
  wire [8:0] T_843;
  wire [8:0] T_845;
  wire [8:0] T_846;
  wire [8:0] T_847;
  wire [8:0] T_848;
  wire [8:0] T_850;
  wire [8:0] T_851;
  wire [7:0] T_853;
  wire [8:0] T_854;
  wire [8:0] T_856;
  wire [8:0] T_857;
  wire [8:0] GEN_41;
  wire [16:0] GEN_42;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire  T_861;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire [52:0] GEN_72;
  wire [52:0] T_865;
  wire [52:0] T_867;
  wire  T_868;
  wire [52:0] T_870;
  wire [52:0] T_871;
  wire [52:0] T_873;
  wire [52:0] T_874;
  wire [33:0] T_875;
  wire [52:0] GEN_73;
  wire [52:0] T_876;
  wire  T_877;
  wire [45:0] T_878;
  wire [45:0] T_880;
  wire [52:0] GEN_74;
  wire [52:0] T_881;
  wire [32:0] T_882;
  wire [45:0] GEN_75;
  wire [45:0] T_883;
  wire [45:0] T_885;
  wire [52:0] GEN_76;
  wire [52:0] T_886;
  wire [45:0] GEN_77;
  wire [45:0] T_887;
  wire [45:0] T_889;
  wire [52:0] GEN_78;
  wire [52:0] T_890;
  wire [52:0] T_892;
  wire [52:0] T_893;
  wire [53:0] GEN_79;
  wire [53:0] T_894;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire  T_900;
  wire [51:0] GEN_80;
  wire [51:0] T_901;
  wire [51:0] T_903;
  wire [50:0] GEN_81;
  wire [50:0] T_904;
  wire [50:0] T_906;
  wire [51:0] GEN_82;
  wire [51:0] T_907;
  wire [52:0] GEN_83;
  wire [52:0] T_908;
  wire [52:0] T_910;
  wire [52:0] GEN_84;
  wire [52:0] T_911;
  wire [52:0] GEN_85;
  wire [52:0] T_912;
  wire [29:0] T_913;
  wire [29:0] T_915;
  wire [52:0] GEN_86;
  wire [52:0] T_916;
  wire [32:0] T_918;
  wire [52:0] GEN_87;
  wire [52:0] T_919;
  wire [53:0] GEN_88;
  wire [53:0] T_920;
  wire  T_921;
  wire  T_922;
  wire  T_923;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire  T_927;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  T_931;
  wire  T_932;
  wire  T_933;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire  T_949;
  wire  T_950;
  wire  T_951;
  wire  T_952;
  wire [1:0] T_953;
  wire [1:0] T_954;
  wire [3:0] T_955;
  wire [104:0] GEN_89;
  wire [104:0] T_956;
  wire [104:0] T_958;
  wire [103:0] GEN_90;
  wire [103:0] T_959;
  wire [103:0] T_961;
  wire [104:0] GEN_91;
  wire [104:0] T_962;
  wire  T_963;
  wire [104:0] GEN_92;
  wire [104:0] T_964;
  wire [104:0] T_966;
  wire [104:0] T_967;
  wire  T_969;
  wire  T_970;
  wire [53:0] GEN_93;
  wire [53:0] T_971;
  wire [53:0] T_973;
  wire [104:0] GEN_94;
  wire [104:0] T_974;
  wire  T_976;
  wire [1:0] T_978;
  wire  T_979;
  wire  T_981;
  wire [1:0] T_983;
  wire [1:0] T_984;
  wire  T_986;
  wire [1:0] T_988;
  wire [1:0] T_989;
  wire [55:0] GEN_95;
  wire [55:0] T_990;
  wire [55:0] T_992;
  wire [104:0] GEN_96;
  wire [104:0] T_993;
  wire [31:0] ESqrR1_B8_sqrt;
  wire [45:0] T_994;
  wire [45:0] T_995;
  wire [45:0] T_997;
  wire [32:0] sqrSigma1_B1;
  wire [57:0] T_998;
  wire  T_999;
  wire  E_C1_div;
  wire  T_1002;
  wire  T_1003;
  wire  T_1004;
  wire [53:0] T_1005;
  wire [53:0] T_1006;
  wire [53:0] T_1008;
  wire  T_1009;
  wire [52:0] T_1011;
  wire [52:0] T_1012;
  wire [53:0] T_1013;
  wire [53:0] T_1015;
  wire [53:0] T_1016;
  wire [53:0] T_1020;
  wire [53:0] sigT_C1;
  wire [55:0] remT_E2;
  wire [31:0] GEN_43;
  wire [57:0] GEN_44;
  wire [32:0] GEN_45;
  wire  T_1021;
  wire  T_1022;
  wire [57:0] GEN_46;
  wire [30:0] T_1023;
  wire [30:0] GEN_47;
  wire [52:0] T_1024;
  wire  T_1025;
  wire  GEN_48;
  wire [52:0] GEN_49;
  wire  GEN_50;
  wire  T_1026;
  wire  T_1027;
  wire  T_1028;
  wire [53:0] T_1029;
  wire  T_1031;
  wire [1:0] T_1034;
  wire  T_1036;
  wire  T_1037;
  wire  T_1038;
  wire  GEN_51;
  wire  GEN_52;
  wire  T_1041;
  wire [13:0] T_1043;
  wire  T_1048;
  wire [13:0] T_1050;
  wire [13:0] T_1051;
  wire [12:0] T_1052;
  wire [13:0] T_1054;
  wire [12:0] T_1055;
  wire [12:0] T_1057;
  wire [13:0] GEN_97;
  wire [13:0] sExpX_E;
  wire [12:0] posExpX_E;
  wire [12:0] T_1058;
  wire  T_1059;
  wire [11:0] T_1060;
  wire  T_1061;
  wire [10:0] T_1062;
  wire  T_1063;
  wire [9:0] T_1064;
  wire  T_1065;
  wire [8:0] T_1066;
  wire  T_1068;
  wire [7:0] T_1069;
  wire  T_1071;
  wire [6:0] T_1072;
  wire  T_1074;
  wire [5:0] T_1075;
  wire [64:0] T_1078;
  wire [49:0] T_1079;
  wire [31:0] T_1080;
  wire [15:0] T_1085;
  wire [31:0] T_1086;
  wire [15:0] T_1087;
  wire [31:0] GEN_98;
  wire [31:0] T_1088;
  wire [31:0] T_1090;
  wire [31:0] T_1091;
  wire [23:0] T_1095;
  wire [31:0] GEN_99;
  wire [31:0] T_1096;
  wire [23:0] T_1097;
  wire [31:0] GEN_100;
  wire [31:0] T_1098;
  wire [31:0] T_1100;
  wire [31:0] T_1101;
  wire [27:0] T_1105;
  wire [31:0] GEN_101;
  wire [31:0] T_1106;
  wire [27:0] T_1107;
  wire [31:0] GEN_102;
  wire [31:0] T_1108;
  wire [31:0] T_1110;
  wire [31:0] T_1111;
  wire [29:0] T_1115;
  wire [31:0] GEN_103;
  wire [31:0] T_1116;
  wire [29:0] T_1117;
  wire [31:0] GEN_104;
  wire [31:0] T_1118;
  wire [31:0] T_1120;
  wire [31:0] T_1121;
  wire [30:0] T_1125;
  wire [31:0] GEN_105;
  wire [31:0] T_1126;
  wire [30:0] T_1127;
  wire [31:0] GEN_106;
  wire [31:0] T_1128;
  wire [31:0] T_1130;
  wire [31:0] T_1131;
  wire [17:0] T_1132;
  wire [15:0] T_1133;
  wire [7:0] T_1138;
  wire [15:0] T_1139;
  wire [7:0] T_1140;
  wire [15:0] GEN_107;
  wire [15:0] T_1141;
  wire [15:0] T_1143;
  wire [15:0] T_1144;
  wire [11:0] T_1148;
  wire [15:0] GEN_108;
  wire [15:0] T_1149;
  wire [11:0] T_1150;
  wire [15:0] GEN_109;
  wire [15:0] T_1151;
  wire [15:0] T_1153;
  wire [15:0] T_1154;
  wire [13:0] T_1158;
  wire [15:0] GEN_110;
  wire [15:0] T_1159;
  wire [13:0] T_1160;
  wire [15:0] GEN_111;
  wire [15:0] T_1161;
  wire [15:0] T_1163;
  wire [15:0] T_1164;
  wire [14:0] T_1168;
  wire [15:0] GEN_112;
  wire [15:0] T_1169;
  wire [14:0] T_1170;
  wire [15:0] GEN_113;
  wire [15:0] T_1171;
  wire [15:0] T_1173;
  wire [15:0] T_1174;
  wire [1:0] T_1175;
  wire  T_1176;
  wire  T_1177;
  wire [1:0] T_1178;
  wire [17:0] T_1179;
  wire [49:0] T_1180;
  wire [49:0] T_1181;
  wire [49:0] T_1182;
  wire [49:0] T_1183;
  wire [49:0] T_1184;
  wire [49:0] T_1185;
  wire [49:0] T_1186;
  wire [49:0] T_1187;
  wire [49:0] T_1188;
  wire [49:0] T_1189;
  wire [49:0] T_1190;
  wire [49:0] T_1191;
  wire [49:0] T_1192;
  wire [52:0] T_1194;
  wire [2:0] T_1205;
  wire [1:0] T_1206;
  wire  T_1207;
  wire  T_1208;
  wire [1:0] T_1209;
  wire  T_1210;
  wire [2:0] T_1211;
  wire [2:0] T_1213;
  wire [2:0] T_1215;
  wire [2:0] T_1217;
  wire [2:0] T_1219;
  wire [52:0] T_1220;
  wire [52:0] T_1222;
  wire [52:0] roundMask_E;
  wire [53:0] T_1225;
  wire [53:0] T_1226;
  wire [53:0] T_1228;
  wire [53:0] incrPosMask_E;
  wire [52:0] T_1229;
  wire [52:0] T_1230;
  wire  hiRoundPosBitT_E;
  wire [51:0] T_1232;
  wire [52:0] GEN_114;
  wire [52:0] T_1235;
  wire [52:0] T_1237;
  wire  all1sHiRoundExtraT_E;
  wire  T_1239;
  wire  T_1241;
  wire  T_1242;
  wire  all1sHiRoundT_E;
  wire [53:0] GEN_116;
  wire [54:0] T_1244;
  wire [53:0] T_1245;
  wire [53:0] GEN_117;
  wire [54:0] T_1246;
  wire [53:0] sigAdjT_E;
  wire [52:0] T_1248;
  wire [53:0] T_1249;
  wire [53:0] sigY0_E;
  wire [53:0] T_1252;
  wire [54:0] T_1254;
  wire [53:0] sigY1_E;
  wire  T_1256;
  wire  T_1258;
  wire  T_1259;
  wire  trueLtX_E1;
  wire  T_1262;
  wire  T_1263;
  wire  T_1264;
  wire  T_1265;
  wire  hiRoundPosBit_E1;
  wire  T_1270;
  wire  T_1272;
  wire  anyRoundExtra_E1;
  wire  T_1273;
  wire  T_1275;
  wire  T_1276;
  wire [53:0] roundEvenMask_E1;
  wire  T_1278;
  wire  T_1281;
  wire  T_1282;
  wire  T_1285;
  wire  T_1288;
  wire  T_1290;
  wire  T_1291;
  wire  T_1292;
  wire  T_1293;
  wire  T_1296;
  wire  T_1300;
  wire  T_1301;
  wire  T_1305;
  wire  T_1306;
  wire  T_1307;
  wire  T_1308;
  wire [53:0] T_1309;
  wire [53:0] T_1310;
  wire [53:0] sigY_E1;
  wire [51:0] fractY_E1;
  wire  inexactY_E1;
  wire  T_1311;
  wire  T_1313;
  wire [13:0] T_1315;
  wire  T_1319;
  wire  T_1320;
  wire [13:0] T_1322;
  wire [13:0] T_1323;
  wire  T_1330;
  wire [13:0] T_1332;
  wire [13:0] T_1333;
  wire  T_1335;
  wire [12:0] T_1336;
  wire [13:0] T_1338;
  wire [12:0] T_1339;
  wire [12:0] T_1341;
  wire [13:0] GEN_118;
  wire [13:0] sExpY_E1;
  wire [11:0] expY_E1;
  wire  T_1342;
  wire  T_1344;
  wire [2:0] T_1346;
  wire  T_1347;
  wire  overflowY_E1;
  wire [12:0] T_1349;
  wire  T_1351;
  wire  totalUnderflowY_E1;
  wire  T_1353;
  wire  T_1354;
  wire  underflowY_E1;
  wire  T_1356;
  wire  T_1359;
  wire  T_1360;
  wire  T_1361;
  wire  T_1362;
  wire  T_1363;
  wire  notSigNaN_invalid_PC;
  wire  T_1366;
  wire  T_1367;
  wire  invalid_PC;
  wire  T_1372;
  wire  T_1375;
  wire  infinity_PC;
  wire  overflow_E1;
  wire  underflow_E1;
  wire  T_1376;
  wire  T_1377;
  wire  inexact_E1;
  wire  T_1378;
  wire  T_1381;
  wire  T_1382;
  wire  notSpecial_isZeroOut_E1;
  wire  T_1383;
  wire  pegMinFiniteMagOut_E1;
  wire  T_1385;
  wire  pegMaxFiniteMagOut_E1;
  wire  T_1386;
  wire  T_1387;
  wire  T_1388;
  wire  notNaN_isInfOut_E1;
  wire  T_1391;
  wire  T_1392;
  wire  isNaNOut_PC;
  wire  T_1394;
  wire  T_1395;
  wire  T_1396;
  wire  signOut_PC;
  wire [11:0] T_1400;
  wire [11:0] T_1401;
  wire [11:0] T_1402;
  wire [11:0] T_1406;
  wire [11:0] T_1407;
  wire [11:0] T_1408;
  wire [11:0] T_1412;
  wire [11:0] T_1413;
  wire [11:0] T_1414;
  wire [11:0] T_1418;
  wire [11:0] T_1419;
  wire [11:0] T_1420;
  wire [11:0] T_1423;
  wire [11:0] T_1424;
  wire [11:0] T_1427;
  wire [11:0] T_1428;
  wire [11:0] T_1431;
  wire [11:0] T_1432;
  wire [11:0] T_1435;
  wire [11:0] expOut_E1;
  wire  T_1436;
  wire  T_1437;
  wire [51:0] T_1441;
  wire [51:0] T_1442;
  wire [51:0] T_1446;
  wire [51:0] fractOut_E1;
  wire [12:0] T_1447;
  wire [64:0] T_1448;
  wire [1:0] T_1449;
  wire [1:0] T_1450;
  wire [2:0] T_1451;
  wire [4:0] T_1452;
  assign io_inReady_div = T_138;
  assign io_inReady_sqrt = T_153;
  assign io_outValid_div = T_371;
  assign io_outValid_sqrt = T_372;
  assign io_out = T_1448;
  assign io_exceptionFlags = T_1452;
  assign io_usingMulAdd = T_955;
  assign io_latchMulAddA_0 = T_864;
  assign io_mulAddA_0 = T_894;
  assign io_latchMulAddB_0 = T_900;
  assign io_mulAddB_0 = T_920;
  assign io_mulAddC_2 = T_993;
  assign ready_PA = T_258;
  assign ready_PB = T_299;
  assign ready_PC = T_368;
  assign leaving_PA = T_255;
  assign leaving_PB = T_296;
  assign leaving_PC = T_365;
  assign cyc_B10_sqrt = T_414;
  assign cyc_B9_sqrt = T_416;
  assign cyc_B8_sqrt = T_418;
  assign cyc_B7_sqrt = T_420;
  assign cyc_B6 = T_422;
  assign cyc_B5 = T_424;
  assign cyc_B4 = T_426;
  assign cyc_B3 = T_428;
  assign cyc_B2 = T_430;
  assign cyc_B1 = T_432;
  assign cyc_B6_div = T_436;
  assign cyc_B5_div = T_440;
  assign cyc_B4_div = T_444;
  assign cyc_B3_div = T_447;
  assign cyc_B2_div = T_450;
  assign cyc_B1_div = T_453;
  assign cyc_B6_sqrt = T_455;
  assign cyc_B5_sqrt = T_457;
  assign cyc_B4_sqrt = T_459;
  assign cyc_B3_sqrt = T_460;
  assign cyc_B2_sqrt = T_461;
  assign cyc_B1_sqrt = T_462;
  assign cyc_C5 = T_475;
  assign cyc_C4 = T_477;
  assign valid_normalCase_leaving_PB = T_479;
  assign cyc_C2 = T_481;
  assign cyc_C1 = T_483;
  assign cyc_E4 = T_503;
  assign cyc_E3 = T_505;
  assign cyc_E2 = T_507;
  assign cyc_E1 = T_509;
  assign zSigma1_B4 = T_997;
  assign sigXNU_B3_CX = T_998;
  assign zComplSigT_C1_sqrt = T_1020;
  assign zComplSigT_C1 = T_1016;
  assign T_113 = cyc_B7_sqrt == 1'h0;
  assign T_114 = ready_PA & T_113;
  assign T_116 = cyc_B6_sqrt == 1'h0;
  assign T_117 = T_114 & T_116;
  assign T_119 = cyc_B5_sqrt == 1'h0;
  assign T_120 = T_117 & T_119;
  assign T_122 = cyc_B4_sqrt == 1'h0;
  assign T_123 = T_120 & T_122;
  assign T_125 = cyc_B3 == 1'h0;
  assign T_126 = T_123 & T_125;
  assign T_128 = cyc_B2 == 1'h0;
  assign T_129 = T_126 & T_128;
  assign T_131 = cyc_B1_sqrt == 1'h0;
  assign T_132 = T_129 & T_131;
  assign T_134 = cyc_C5 == 1'h0;
  assign T_135 = T_132 & T_134;
  assign T_137 = cyc_C4 == 1'h0;
  assign T_138 = T_135 & T_137;
  assign T_141 = ready_PA & T_116;
  assign T_144 = T_141 & T_119;
  assign T_147 = T_144 & T_122;
  assign T_149 = cyc_B2_div == 1'h0;
  assign T_150 = T_147 & T_149;
  assign T_153 = T_150 & T_131;
  assign T_154 = io_inReady_div & io_inValid;
  assign T_156 = io_sqrtOp == 1'h0;
  assign cyc_S_div = T_154 & T_156;
  assign T_157 = io_inReady_sqrt & io_inValid;
  assign cyc_S_sqrt = T_157 & io_sqrtOp;
  assign cyc_S = cyc_S_div | cyc_S_sqrt;
  assign signA_S = io_a[64];
  assign expA_S = io_a[63:52];
  assign fractA_S = io_a[51:0];
  assign specialCodeA_S = expA_S[11:9];
  assign isZeroA_S = specialCodeA_S == 3'h0;
  assign T_159 = specialCodeA_S[2:1];
  assign isSpecialA_S = T_159 == 2'h3;
  assign signB_S = io_b[64];
  assign expB_S = io_b[63:52];
  assign fractB_S = io_b[51:0];
  assign specialCodeB_S = expB_S[11:9];
  assign isZeroB_S = specialCodeB_S == 3'h0;
  assign T_162 = specialCodeB_S[2:1];
  assign isSpecialB_S = T_162 == 2'h3;
  assign T_164 = signA_S ^ signB_S;
  assign sign_S = io_sqrtOp ? signB_S : T_164;
  assign T_166 = isSpecialA_S == 1'h0;
  assign T_168 = isSpecialB_S == 1'h0;
  assign T_169 = T_166 & T_168;
  assign T_171 = isZeroA_S == 1'h0;
  assign T_172 = T_169 & T_171;
  assign T_174 = isZeroB_S == 1'h0;
  assign normalCase_S_div = T_172 & T_174;
  assign T_179 = T_168 & T_174;
  assign T_181 = signB_S == 1'h0;
  assign normalCase_S_sqrt = T_179 & T_181;
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div;
  assign entering_PA_normalCase_div = cyc_S_div & normalCase_S_div;
  assign entering_PA_normalCase_sqrt = cyc_S_sqrt & normalCase_S_sqrt;
  assign entering_PA_normalCase = entering_PA_normalCase_div | entering_PA_normalCase_sqrt;
  assign T_183 = ready_PB == 1'h0;
  assign T_184 = valid_PA | T_183;
  assign T_185 = cyc_S & T_184;
  assign entering_PA = entering_PA_normalCase | T_185;
  assign T_187 = normalCase_S == 1'h0;
  assign T_188 = cyc_S & T_187;
  assign T_190 = valid_PA == 1'h0;
  assign T_191 = T_188 & T_190;
  assign T_193 = valid_PB == 1'h0;
  assign T_195 = ready_PC == 1'h0;
  assign T_196 = T_193 & T_195;
  assign T_197 = leaving_PB | T_196;
  assign entering_PB_S = T_191 & T_197;
  assign T_206 = T_191 & T_193;
  assign entering_PC_S = T_206 & ready_PC;
  assign T_207 = entering_PA | leaving_PA;
  assign GEN_0 = T_207 ? entering_PA : valid_PA;
  assign T_208 = fractB_S[51];
  assign GEN_1 = entering_PA ? io_sqrtOp : sqrtOp_PA;
  assign GEN_2 = entering_PA ? sign_S : sign_PA;
  assign GEN_3 = entering_PA ? specialCodeB_S : specialCodeB_PA;
  assign GEN_4 = entering_PA ? T_208 : fractB_51_PA;
  assign GEN_5 = entering_PA ? io_roundingMode : roundingMode_PA;
  assign T_211 = entering_PA & T_156;
  assign T_212 = fractA_S[51];
  assign GEN_6 = T_211 ? specialCodeA_S : specialCodeA_PA;
  assign GEN_7 = T_211 ? T_212 : fractA_51_PA;
  assign T_213 = expB_S[11];
  assign T_217 = T_213 ? 3'h7 : 3'h0;
  assign T_218 = expB_S[10:0];
  assign T_219 = ~ T_218;
  assign T_220 = {T_217,T_219};
  assign GEN_53 = {{2'd0}, expA_S};
  assign T_221 = GEN_53 + T_220;
  assign T_222 = T_221[13:0];
  assign T_223 = io_sqrtOp ? {{2'd0}, expB_S} : T_222;
  assign T_224 = fractB_S[50:0];
  assign GEN_8 = entering_PA_normalCase ? T_223 : exp_PA;
  assign GEN_9 = entering_PA_normalCase ? T_224 : fractB_other_PA;
  assign T_225 = fractA_S[50:0];
  assign GEN_10 = entering_PA_normalCase_div ? T_225 : fractA_other_PA;
  assign isZeroA_PA = specialCodeA_PA == 3'h0;
  assign T_227 = specialCodeA_PA[2:1];
  assign isSpecialA_PA = T_227 == 2'h3;
  assign T_230 = {1'h1,fractA_51_PA};
  assign sigA_PA = {T_230,fractA_other_PA};
  assign isZeroB_PA = specialCodeB_PA == 3'h0;
  assign T_232 = specialCodeB_PA[2:1];
  assign isSpecialB_PA = T_232 == 2'h3;
  assign T_235 = {1'h1,fractB_51_PA};
  assign sigB_PA = {T_235,fractB_other_PA};
  assign T_237 = isSpecialB_PA == 1'h0;
  assign T_239 = isZeroB_PA == 1'h0;
  assign T_240 = T_237 & T_239;
  assign T_242 = sign_PA == 1'h0;
  assign T_243 = T_240 & T_242;
  assign T_245 = isSpecialA_PA == 1'h0;
  assign T_248 = T_245 & T_237;
  assign T_250 = isZeroA_PA == 1'h0;
  assign T_251 = T_248 & T_250;
  assign T_254 = T_251 & T_239;
  assign normalCase_PA = sqrtOp_PA ? T_243 : T_254;
  assign valid_normalCase_leaving_PA = cyc_B4_div | cyc_B7_sqrt;
  assign valid_leaving_PA = normalCase_PA ? valid_normalCase_leaving_PA : ready_PB;
  assign T_255 = valid_PA & valid_leaving_PA;
  assign T_258 = T_190 | valid_leaving_PA;
  assign T_259 = valid_PA & normalCase_PA;
  assign entering_PB_normalCase = T_259 & valid_normalCase_leaving_PA;
  assign entering_PB = entering_PB_S | leaving_PA;
  assign T_260 = entering_PB | leaving_PB;
  assign GEN_11 = T_260 ? entering_PB : valid_PB;
  assign T_261 = valid_PA ? sqrtOp_PA : io_sqrtOp;
  assign T_262 = valid_PA ? sign_PA : sign_S;
  assign T_263 = valid_PA ? specialCodeA_PA : specialCodeA_S;
  assign T_265 = valid_PA ? fractA_51_PA : T_212;
  assign T_266 = valid_PA ? specialCodeB_PA : specialCodeB_S;
  assign T_268 = valid_PA ? fractB_51_PA : T_208;
  assign T_269 = valid_PA ? roundingMode_PA : io_roundingMode;
  assign GEN_12 = entering_PB ? T_261 : sqrtOp_PB;
  assign GEN_13 = entering_PB ? T_262 : sign_PB;
  assign GEN_14 = entering_PB ? T_263 : specialCodeA_PB;
  assign GEN_15 = entering_PB ? T_265 : fractA_51_PB;
  assign GEN_16 = entering_PB ? T_266 : specialCodeB_PB;
  assign GEN_17 = entering_PB ? T_268 : fractB_51_PB;
  assign GEN_18 = entering_PB ? T_269 : roundingMode_PB;
  assign T_270 = fractA_other_PA[0];
  assign GEN_19 = entering_PB_normalCase ? exp_PA : exp_PB;
  assign GEN_20 = entering_PB_normalCase ? T_270 : fractA_0_PB;
  assign GEN_21 = entering_PB_normalCase ? fractB_other_PA : fractB_other_PB;
  assign isZeroA_PB = specialCodeA_PB == 3'h0;
  assign T_272 = specialCodeA_PB[2:1];
  assign isSpecialA_PB = T_272 == 2'h3;
  assign isZeroB_PB = specialCodeB_PB == 3'h0;
  assign T_275 = specialCodeB_PB[2:1];
  assign isSpecialB_PB = T_275 == 2'h3;
  assign T_278 = isSpecialB_PB == 1'h0;
  assign T_280 = isZeroB_PB == 1'h0;
  assign T_281 = T_278 & T_280;
  assign T_283 = sign_PB == 1'h0;
  assign T_284 = T_281 & T_283;
  assign T_286 = isSpecialA_PB == 1'h0;
  assign T_289 = T_286 & T_278;
  assign T_291 = isZeroA_PB == 1'h0;
  assign T_292 = T_289 & T_291;
  assign T_295 = T_292 & T_280;
  assign normalCase_PB = sqrtOp_PB ? T_284 : T_295;
  assign valid_leaving_PB = normalCase_PB ? valid_normalCase_leaving_PB : ready_PC;
  assign T_296 = valid_PB & valid_leaving_PB;
  assign T_299 = T_193 | valid_leaving_PB;
  assign T_300 = valid_PB & normalCase_PB;
  assign entering_PC_normalCase = T_300 & valid_normalCase_leaving_PB;
  assign entering_PC = entering_PC_S | leaving_PB;
  assign T_301 = entering_PC | leaving_PC;
  assign GEN_22 = T_301 ? entering_PC : valid_PC;
  assign T_302 = valid_PB ? sqrtOp_PB : io_sqrtOp;
  assign T_303 = valid_PB ? sign_PB : sign_S;
  assign T_304 = valid_PB ? specialCodeA_PB : specialCodeA_S;
  assign T_306 = valid_PB ? fractA_51_PB : T_212;
  assign T_307 = valid_PB ? specialCodeB_PB : specialCodeB_S;
  assign T_309 = valid_PB ? fractB_51_PB : T_208;
  assign T_310 = valid_PB ? roundingMode_PB : io_roundingMode;
  assign GEN_23 = entering_PC ? T_302 : sqrtOp_PC;
  assign GEN_24 = entering_PC ? T_303 : sign_PC;
  assign GEN_25 = entering_PC ? T_304 : specialCodeA_PC;
  assign GEN_26 = entering_PC ? T_306 : fractA_51_PC;
  assign GEN_27 = entering_PC ? T_307 : specialCodeB_PC;
  assign GEN_28 = entering_PC ? T_309 : fractB_51_PC;
  assign GEN_29 = entering_PC ? T_310 : roundingMode_PC;
  assign GEN_30 = entering_PC_normalCase ? exp_PB : exp_PC;
  assign GEN_31 = entering_PC_normalCase ? fractA_0_PB : fractA_0_PC;
  assign GEN_32 = entering_PC_normalCase ? fractB_other_PB : fractB_other_PC;
  assign isZeroA_PC = specialCodeA_PC == 3'h0;
  assign T_312 = specialCodeA_PC[2:1];
  assign isSpecialA_PC = T_312 == 2'h3;
  assign T_314 = specialCodeA_PC[0];
  assign T_316 = T_314 == 1'h0;
  assign isInfA_PC = isSpecialA_PC & T_316;
  assign isNaNA_PC = isSpecialA_PC & T_314;
  assign T_319 = fractA_51_PC == 1'h0;
  assign isSigNaNA_PC = isNaNA_PC & T_319;
  assign isZeroB_PC = specialCodeB_PC == 3'h0;
  assign T_321 = specialCodeB_PC[2:1];
  assign isSpecialB_PC = T_321 == 2'h3;
  assign T_323 = specialCodeB_PC[0];
  assign T_325 = T_323 == 1'h0;
  assign isInfB_PC = isSpecialB_PC & T_325;
  assign isNaNB_PC = isSpecialB_PC & T_323;
  assign T_328 = fractB_51_PC == 1'h0;
  assign isSigNaNB_PC = isNaNB_PC & T_328;
  assign T_330 = {1'h1,fractB_51_PC};
  assign sigB_PC = {T_330,fractB_other_PC};
  assign T_332 = isSpecialB_PC == 1'h0;
  assign T_334 = isZeroB_PC == 1'h0;
  assign T_335 = T_332 & T_334;
  assign T_337 = sign_PC == 1'h0;
  assign T_338 = T_335 & T_337;
  assign T_340 = isSpecialA_PC == 1'h0;
  assign T_343 = T_340 & T_332;
  assign T_345 = isZeroA_PC == 1'h0;
  assign T_346 = T_343 & T_345;
  assign T_349 = T_346 & T_334;
  assign normalCase_PC = sqrtOp_PC ? T_338 : T_349;
  assign T_351 = exp_PC + 14'h2;
  assign expP2_PC = T_351[13:0];
  assign T_352 = exp_PC[0];
  assign T_353 = expP2_PC[13:1];
  assign T_355 = {T_353,1'h0};
  assign T_356 = exp_PC[13:1];
  assign T_358 = {T_356,1'h1};
  assign expP1_PC = T_352 ? T_355 : T_358;
  assign roundingMode_near_even_PC = roundingMode_PC == 2'h0;
  assign roundingMode_min_PC = roundingMode_PC == 2'h2;
  assign roundingMode_max_PC = roundingMode_PC == 2'h3;
  assign roundMagUp_PC = sign_PC ? roundingMode_min_PC : roundingMode_max_PC;
  assign overflowY_roundMagUp_PC = roundingMode_near_even_PC | roundMagUp_PC;
  assign T_360 = roundMagUp_PC == 1'h0;
  assign T_362 = roundingMode_near_even_PC == 1'h0;
  assign roundMagDown_PC = T_360 & T_362;
  assign T_364 = normalCase_PC == 1'h0;
  assign valid_leaving_PC = T_364 | cyc_E1;
  assign T_365 = valid_PC & valid_leaving_PC;
  assign T_367 = valid_PC == 1'h0;
  assign T_368 = T_367 | valid_leaving_PC;
  assign T_370 = sqrtOp_PC == 1'h0;
  assign T_371 = leaving_PC & T_370;
  assign T_372 = leaving_PC & sqrtOp_PC;
  assign T_374 = cycleNum_A != 3'h0;
  assign T_375 = entering_PA_normalCase | T_374;
  assign T_378 = entering_PA_normalCase_div ? 2'h3 : 2'h0;
  assign T_381 = entering_PA_normalCase_sqrt ? 3'h6 : 3'h0;
  assign GEN_54 = {{1'd0}, T_378};
  assign T_382 = GEN_54 | T_381;
  assign T_384 = entering_PA_normalCase == 1'h0;
  assign T_386 = cycleNum_A - 3'h1;
  assign T_387 = T_386[2:0];
  assign T_389 = T_384 ? T_387 : 3'h0;
  assign T_390 = T_382 | T_389;
  assign GEN_33 = T_375 ? T_390 : cycleNum_A;
  assign cyc_A6_sqrt = cycleNum_A == 3'h6;
  assign cyc_A5_sqrt = cycleNum_A == 3'h5;
  assign cyc_A4_sqrt = cycleNum_A == 3'h4;
  assign cyc_A4 = cyc_A4_sqrt | entering_PA_normalCase_div;
  assign cyc_A3 = cycleNum_A == 3'h3;
  assign cyc_A2 = cycleNum_A == 3'h2;
  assign cyc_A1 = cycleNum_A == 3'h1;
  assign T_398 = sqrtOp_PA == 1'h0;
  assign cyc_A3_div = cyc_A3 & T_398;
  assign cyc_A2_div = cyc_A2 & T_398;
  assign cyc_A1_div = cyc_A1 & T_398;
  assign cyc_A3_sqrt = cyc_A3 & sqrtOp_PA;
  assign cyc_A1_sqrt = cyc_A1 & sqrtOp_PA;
  assign T_404 = cycleNum_B != 4'h0;
  assign T_405 = cyc_A1 | T_404;
  assign T_408 = sqrtOp_PA ? 4'ha : 4'h6;
  assign T_410 = cycleNum_B - 4'h1;
  assign T_411 = T_410[3:0];
  assign T_412 = cyc_A1 ? T_408 : T_411;
  assign GEN_34 = T_405 ? T_412 : cycleNum_B;
  assign T_414 = cycleNum_B == 4'ha;
  assign T_416 = cycleNum_B == 4'h9;
  assign T_418 = cycleNum_B == 4'h8;
  assign T_420 = cycleNum_B == 4'h7;
  assign T_422 = cycleNum_B == 4'h6;
  assign T_424 = cycleNum_B == 4'h5;
  assign T_426 = cycleNum_B == 4'h4;
  assign T_428 = cycleNum_B == 4'h3;
  assign T_430 = cycleNum_B == 4'h2;
  assign T_432 = cycleNum_B == 4'h1;
  assign T_433 = cyc_B6 & valid_PA;
  assign T_436 = T_433 & T_398;
  assign T_437 = cyc_B5 & valid_PA;
  assign T_440 = T_437 & T_398;
  assign T_441 = cyc_B4 & valid_PA;
  assign T_444 = T_441 & T_398;
  assign T_446 = sqrtOp_PB == 1'h0;
  assign T_447 = cyc_B3 & T_446;
  assign T_450 = cyc_B2 & T_446;
  assign T_453 = cyc_B1 & T_446;
  assign T_454 = cyc_B6 & valid_PB;
  assign T_455 = T_454 & sqrtOp_PB;
  assign T_456 = cyc_B5 & valid_PB;
  assign T_457 = T_456 & sqrtOp_PB;
  assign T_458 = cyc_B4 & valid_PB;
  assign T_459 = T_458 & sqrtOp_PB;
  assign T_460 = cyc_B3 & sqrtOp_PB;
  assign T_461 = cyc_B2 & sqrtOp_PB;
  assign T_462 = cyc_B1 & sqrtOp_PB;
  assign T_464 = cycleNum_C != 3'h0;
  assign T_465 = cyc_B1 | T_464;
  assign T_468 = sqrtOp_PB ? 3'h6 : 3'h5;
  assign T_470 = cycleNum_C - 3'h1;
  assign T_471 = T_470[2:0];
  assign T_472 = cyc_B1 ? T_468 : T_471;
  assign GEN_35 = T_465 ? T_472 : cycleNum_C;
  assign cyc_C6_sqrt = cycleNum_C == 3'h6;
  assign T_475 = cycleNum_C == 3'h5;
  assign T_477 = cycleNum_C == 3'h4;
  assign T_479 = cycleNum_C == 3'h3;
  assign T_481 = cycleNum_C == 3'h2;
  assign T_483 = cycleNum_C == 3'h1;
  assign cyc_C5_div = cyc_C5 & T_446;
  assign cyc_C4_div = cyc_C4 & T_446;
  assign cyc_C1_div = cyc_C1 & T_370;
  assign cyc_C5_sqrt = cyc_C5 & sqrtOp_PB;
  assign cyc_C4_sqrt = cyc_C4 & sqrtOp_PB;
  assign cyc_C3_sqrt = valid_normalCase_leaving_PB & sqrtOp_PB;
  assign cyc_C1_sqrt = cyc_C1 & sqrtOp_PC;
  assign T_495 = cycleNum_E != 3'h0;
  assign T_496 = cyc_C1 | T_495;
  assign T_499 = cycleNum_E - 3'h1;
  assign T_500 = T_499[2:0];
  assign T_501 = cyc_C1 ? 3'h4 : T_500;
  assign GEN_36 = T_496 ? T_501 : cycleNum_E;
  assign T_503 = cycleNum_E == 3'h4;
  assign T_505 = cycleNum_E == 3'h3;
  assign T_507 = cycleNum_E == 3'h2;
  assign T_509 = cycleNum_E == 3'h1;
  assign cyc_E3_div = cyc_E3 & T_370;
  assign cyc_E3_sqrt = cyc_E3 & sqrtOp_PC;
  assign zFractB_A4_div = entering_PA_normalCase_div ? fractB_S : 52'h0;
  assign T_519 = fractB_S[51:49];
  assign T_521 = T_519 == 3'h0;
  assign zLinPiece_0_A4_div = entering_PA_normalCase_div & T_521;
  assign T_524 = T_519 == 3'h1;
  assign zLinPiece_1_A4_div = entering_PA_normalCase_div & T_524;
  assign T_527 = T_519 == 3'h2;
  assign zLinPiece_2_A4_div = entering_PA_normalCase_div & T_527;
  assign T_530 = T_519 == 3'h3;
  assign zLinPiece_3_A4_div = entering_PA_normalCase_div & T_530;
  assign T_533 = T_519 == 3'h4;
  assign zLinPiece_4_A4_div = entering_PA_normalCase_div & T_533;
  assign T_536 = T_519 == 3'h5;
  assign zLinPiece_5_A4_div = entering_PA_normalCase_div & T_536;
  assign T_539 = T_519 == 3'h6;
  assign zLinPiece_6_A4_div = entering_PA_normalCase_div & T_539;
  assign T_542 = T_519 == 3'h7;
  assign zLinPiece_7_A4_div = entering_PA_normalCase_div & T_542;
  assign T_545 = zLinPiece_0_A4_div ? 9'h1c7 : 9'h0;
  assign T_548 = zLinPiece_1_A4_div ? 9'h16c : 9'h0;
  assign T_549 = T_545 | T_548;
  assign T_552 = zLinPiece_2_A4_div ? 9'h12a : 9'h0;
  assign T_553 = T_549 | T_552;
  assign T_556 = zLinPiece_3_A4_div ? 9'hf8 : 9'h0;
  assign T_557 = T_553 | T_556;
  assign T_560 = zLinPiece_4_A4_div ? 9'hd2 : 9'h0;
  assign T_561 = T_557 | T_560;
  assign T_564 = zLinPiece_5_A4_div ? 9'hb4 : 9'h0;
  assign T_565 = T_561 | T_564;
  assign T_568 = zLinPiece_6_A4_div ? 9'h9c : 9'h0;
  assign T_569 = T_565 | T_568;
  assign T_572 = zLinPiece_7_A4_div ? 9'h89 : 9'h0;
  assign zK1_A4_div = T_569 | T_572;
  assign T_576 = zLinPiece_0_A4_div ? 12'h1c : 12'h0;
  assign T_580 = zLinPiece_1_A4_div ? 12'h3a2 : 12'h0;
  assign T_581 = T_576 | T_580;
  assign T_585 = zLinPiece_2_A4_div ? 12'h675 : 12'h0;
  assign T_586 = T_581 | T_585;
  assign T_590 = zLinPiece_3_A4_div ? 12'h8c6 : 12'h0;
  assign T_591 = T_586 | T_590;
  assign T_595 = zLinPiece_4_A4_div ? 12'hab4 : 12'h0;
  assign T_596 = T_591 | T_595;
  assign T_600 = zLinPiece_5_A4_div ? 12'hc56 : 12'h0;
  assign T_601 = T_596 | T_600;
  assign T_605 = zLinPiece_6_A4_div ? 12'hdbd : 12'h0;
  assign T_606 = T_601 | T_605;
  assign T_610 = zLinPiece_7_A4_div ? 12'hef4 : 12'h0;
  assign zComplFractK0_A4_div = T_606 | T_610;
  assign zFractB_A7_sqrt = entering_PA_normalCase_sqrt ? fractB_S : 52'h0;
  assign T_612 = expB_S[0];
  assign T_614 = T_612 == 1'h0;
  assign T_615 = entering_PA_normalCase_sqrt & T_614;
  assign T_618 = T_208 == 1'h0;
  assign zQuadPiece_0_A7_sqrt = T_615 & T_618;
  assign zQuadPiece_1_A7_sqrt = T_615 & T_208;
  assign T_625 = entering_PA_normalCase_sqrt & T_612;
  assign zQuadPiece_2_A7_sqrt = T_625 & T_618;
  assign zQuadPiece_3_A7_sqrt = T_625 & T_208;
  assign T_634 = zQuadPiece_0_A7_sqrt ? 9'h1c8 : 9'h0;
  assign T_637 = zQuadPiece_1_A7_sqrt ? 9'hc1 : 9'h0;
  assign T_638 = T_634 | T_637;
  assign T_641 = zQuadPiece_2_A7_sqrt ? 9'h143 : 9'h0;
  assign T_642 = T_638 | T_641;
  assign T_645 = zQuadPiece_3_A7_sqrt ? 9'h89 : 9'h0;
  assign zK2_A7_sqrt = T_642 | T_645;
  assign T_649 = zQuadPiece_0_A7_sqrt ? 10'h2f : 10'h0;
  assign T_653 = zQuadPiece_1_A7_sqrt ? 10'h1df : 10'h0;
  assign T_654 = T_649 | T_653;
  assign T_658 = zQuadPiece_2_A7_sqrt ? 10'h14d : 10'h0;
  assign T_659 = T_654 | T_658;
  assign T_663 = zQuadPiece_3_A7_sqrt ? 10'h27e : 10'h0;
  assign zComplK1_A7_sqrt = T_659 | T_663;
  assign T_664 = exp_PA[0];
  assign T_666 = T_664 == 1'h0;
  assign T_667 = cyc_A6_sqrt & T_666;
  assign T_668 = sigB_PA[51];
  assign T_670 = T_668 == 1'h0;
  assign zQuadPiece_0_A6_sqrt = T_667 & T_670;
  assign zQuadPiece_1_A6_sqrt = T_667 & T_668;
  assign T_677 = cyc_A6_sqrt & T_664;
  assign zQuadPiece_2_A6_sqrt = T_677 & T_670;
  assign zQuadPiece_3_A6_sqrt = T_677 & T_668;
  assign T_687 = zQuadPiece_0_A6_sqrt ? 13'h1a : 13'h0;
  assign T_691 = zQuadPiece_1_A6_sqrt ? 13'hbca : 13'h0;
  assign T_692 = T_687 | T_691;
  assign T_696 = zQuadPiece_2_A6_sqrt ? 13'h12d3 : 13'h0;
  assign T_697 = T_692 | T_696;
  assign T_701 = zQuadPiece_3_A6_sqrt ? 13'h1b17 : 13'h0;
  assign zComplFractK0_A6_sqrt = T_697 | T_701;
  assign T_702 = zFractB_A4_div[48:40];
  assign T_703 = T_702 | zK2_A7_sqrt;
  assign T_705 = cyc_S == 1'h0;
  assign T_707 = T_705 ? nextMulAdd9A_A : 9'h0;
  assign mulAdd9A_A = T_703 | T_707;
  assign T_708 = zFractB_A7_sqrt[50:42];
  assign T_709 = zK1_A4_div | T_708;
  assign T_713 = T_705 ? nextMulAdd9B_A : 9'h0;
  assign mulAdd9B_A = T_709 | T_713;
  assign T_717 = entering_PA_normalCase_sqrt ? 10'h3ff : 10'h0;
  assign T_718 = {zComplK1_A7_sqrt,T_717};
  assign T_722 = cyc_A6_sqrt ? 6'h3f : 6'h0;
  assign T_723 = {cyc_A6_sqrt,zComplFractK0_A6_sqrt};
  assign T_724 = {T_723,T_722};
  assign T_725 = T_718 | T_724;
  assign T_729 = entering_PA_normalCase_div ? 8'hff : 8'h0;
  assign T_730 = {entering_PA_normalCase_div,zComplFractK0_A4_div};
  assign T_731 = {T_730,T_729};
  assign GEN_55 = {{1'd0}, T_725};
  assign T_732 = GEN_55 | T_731;
  assign GEN_56 = {{10'd0}, fractR0_A};
  assign T_734 = GEN_56 << 10;
  assign GEN_57 = {{1'd0}, T_734};
  assign T_735 = 20'h40000 + GEN_57;
  assign T_736 = T_735[19:0];
  assign T_738 = cyc_A5_sqrt ? T_736 : 20'h0;
  assign GEN_58 = {{1'd0}, T_738};
  assign T_739 = T_732 | GEN_58;
  assign T_740 = hiSqrR0_A_sqrt[9];
  assign T_742 = T_740 == 1'h0;
  assign T_743 = cyc_A4_sqrt & T_742;
  assign T_746 = T_743 ? 11'h400 : 11'h0;
  assign GEN_59 = {{10'd0}, T_746};
  assign T_747 = T_739 | GEN_59;
  assign T_749 = cyc_A4_sqrt & T_740;
  assign T_750 = T_749 | cyc_A3_div;
  assign T_751 = sigB_PA[46:26];
  assign T_753 = T_751 + 21'h400;
  assign T_754 = T_753[20:0];
  assign T_756 = T_750 ? T_754 : 21'h0;
  assign T_757 = T_747 | T_756;
  assign T_758 = cyc_A3_sqrt | cyc_A2;
  assign T_760 = T_758 ? partNegSigma0_A : 21'h0;
  assign T_761 = T_757 | T_760;
  assign GEN_60 = {{16'd0}, fractR0_A};
  assign T_762 = GEN_60 << 16;
  assign T_764 = cyc_A1_sqrt ? T_762 : 25'h0;
  assign GEN_61 = {{4'd0}, T_761};
  assign T_765 = GEN_61 | T_764;
  assign GEN_62 = {{15'd0}, fractR0_A};
  assign T_766 = GEN_62 << 15;
  assign T_768 = cyc_A1_div ? T_766 : 24'h0;
  assign GEN_63 = {{1'd0}, T_768};
  assign mulAdd9C_A = T_765 | GEN_63;
  assign T_769 = mulAdd9A_A * mulAdd9B_A;
  assign T_771 = mulAdd9C_A[17:0];
  assign T_772 = {1'h0,T_771};
  assign GEN_64 = {{1'd0}, T_769};
  assign T_773 = GEN_64 + T_772;
  assign loMulAdd9Out_A = T_773[18:0];
  assign T_774 = loMulAdd9Out_A[18];
  assign T_775 = mulAdd9C_A[24:18];
  assign T_777 = T_775 + 7'h1;
  assign T_778 = T_777[6:0];
  assign T_780 = T_774 ? T_778 : T_775;
  assign T_781 = loMulAdd9Out_A[17:0];
  assign mulAdd9Out_A = {T_780,T_781};
  assign T_782 = mulAdd9Out_A[19];
  assign T_783 = cyc_A6_sqrt & T_782;
  assign T_784 = ~ mulAdd9Out_A;
  assign T_785 = T_784[24:10];
  assign T_787 = T_783 ? T_785 : 15'h0;
  assign zFractR0_A6_sqrt = T_787[8:0];
  assign GEN_65 = {{1'd0}, mulAdd9Out_A};
  assign T_789 = GEN_65 << 1;
  assign sqrR0_A5_sqrt = T_664 ? T_789 : {{1'd0}, mulAdd9Out_A};
  assign T_790 = mulAdd9Out_A[20];
  assign T_791 = entering_PA_normalCase_div & T_790;
  assign T_793 = T_784[24:11];
  assign T_795 = T_791 ? T_793 : 14'h0;
  assign zFractR0_A4_div = T_795[8:0];
  assign T_796 = mulAdd9Out_A[11];
  assign T_797 = cyc_A2 & T_796;
  assign T_799 = T_784[24:2];
  assign T_801 = T_797 ? T_799 : 23'h0;
  assign zSigma0_A2 = T_801[8:0];
  assign T_802 = mulAdd9Out_A[24:10];
  assign T_803 = mulAdd9Out_A[24:9];
  assign T_804 = sqrtOp_PA ? {{1'd0}, T_802} : T_803;
  assign fractR1_A1 = T_804[14:0];
  assign r1_A1 = {1'h1,fractR1_A1};
  assign GEN_66 = {{1'd0}, r1_A1};
  assign T_807 = GEN_66 << 1;
  assign ER1_A1_sqrt = T_664 ? T_807 : {{1'd0}, r1_A1};
  assign T_808 = cyc_A6_sqrt | entering_PA_normalCase_div;
  assign T_809 = zFractR0_A6_sqrt | zFractR0_A4_div;
  assign GEN_37 = T_808 ? T_809 : fractR0_A;
  assign T_810 = sqrR0_A5_sqrt[25:10];
  assign GEN_38 = cyc_A5_sqrt ? T_810 : {{6'd0}, hiSqrR0_A_sqrt};
  assign T_811 = cyc_A4_sqrt | cyc_A3;
  assign T_813 = cyc_A4_sqrt ? mulAdd9Out_A : {{9'd0}, T_803};
  assign T_814 = T_813[20:0];
  assign GEN_39 = T_811 ? T_814 : partNegSigma0_A;
  assign T_815 = entering_PA_normalCase_sqrt | cyc_A6_sqrt;
  assign T_816 = T_815 | cyc_A5_sqrt;
  assign T_817 = T_816 | cyc_A4;
  assign T_818 = T_817 | cyc_A3;
  assign T_819 = T_818 | cyc_A2;
  assign T_823 = entering_PA_normalCase_sqrt ? T_793 : 14'h0;
  assign GEN_67 = {{5'd0}, zFractR0_A6_sqrt};
  assign T_824 = T_823 | GEN_67;
  assign T_825 = sigB_PA[43:35];
  assign T_827 = cyc_A4_sqrt ? T_825 : 9'h0;
  assign GEN_68 = {{5'd0}, T_827};
  assign T_828 = T_824 | GEN_68;
  assign T_829 = zFractB_A4_div[43:35];
  assign GEN_69 = {{5'd0}, T_829};
  assign T_830 = T_828 | GEN_69;
  assign T_831 = cyc_A5_sqrt | cyc_A3;
  assign T_832 = sigB_PA[52:44];
  assign T_834 = T_831 ? T_832 : 9'h0;
  assign GEN_70 = {{5'd0}, T_834};
  assign T_835 = T_830 | GEN_70;
  assign GEN_71 = {{5'd0}, zSigma0_A2};
  assign T_836 = T_835 | GEN_71;
  assign GEN_40 = T_819 ? T_836 : {{5'd0}, nextMulAdd9A_A};
  assign T_840 = T_817 | cyc_A2;
  assign T_842 = T_708 | zFractR0_A6_sqrt;
  assign T_843 = sqrR0_A5_sqrt[9:1];
  assign T_845 = cyc_A5_sqrt ? T_843 : 9'h0;
  assign T_846 = T_842 | T_845;
  assign T_847 = T_846 | zFractR0_A4_div;
  assign T_848 = hiSqrR0_A_sqrt[8:0];
  assign T_850 = cyc_A4_sqrt ? T_848 : 9'h0;
  assign T_851 = T_847 | T_850;
  assign T_853 = fractR0_A[8:1];
  assign T_854 = {1'h1,T_853};
  assign T_856 = cyc_A2 ? T_854 : 9'h0;
  assign T_857 = T_851 | T_856;
  assign GEN_41 = T_840 ? T_857 : nextMulAdd9B_A;
  assign GEN_42 = cyc_A1_sqrt ? ER1_A1_sqrt : ER1_B_sqrt;
  assign T_858 = cyc_A1 | cyc_B7_sqrt;
  assign T_859 = T_858 | cyc_B6_div;
  assign T_860 = T_859 | cyc_B4;
  assign T_861 = T_860 | cyc_B3;
  assign T_862 = T_861 | cyc_C6_sqrt;
  assign T_863 = T_862 | cyc_C4;
  assign T_864 = T_863 | cyc_C1;
  assign GEN_72 = {{36'd0}, ER1_A1_sqrt};
  assign T_865 = GEN_72 << 36;
  assign T_867 = cyc_A1_sqrt ? T_865 : 53'h0;
  assign T_868 = cyc_B7_sqrt | cyc_A1_div;
  assign T_870 = T_868 ? sigB_PA : 53'h0;
  assign T_871 = T_867 | T_870;
  assign T_873 = cyc_B6_div ? sigA_PA : 53'h0;
  assign T_874 = T_871 | T_873;
  assign T_875 = zSigma1_B4[45:12];
  assign GEN_73 = {{19'd0}, T_875};
  assign T_876 = T_874 | GEN_73;
  assign T_877 = cyc_B3 | cyc_C6_sqrt;
  assign T_878 = sigXNU_B3_CX[57:12];
  assign T_880 = T_877 ? T_878 : 46'h0;
  assign GEN_74 = {{7'd0}, T_880};
  assign T_881 = T_876 | GEN_74;
  assign T_882 = sigXN_C[57:25];
  assign GEN_75 = {{13'd0}, T_882};
  assign T_883 = GEN_75 << 13;
  assign T_885 = cyc_C4_div ? T_883 : 46'h0;
  assign GEN_76 = {{7'd0}, T_885};
  assign T_886 = T_881 | GEN_76;
  assign GEN_77 = {{15'd0}, u_C_sqrt};
  assign T_887 = GEN_77 << 15;
  assign T_889 = cyc_C4_sqrt ? T_887 : 46'h0;
  assign GEN_78 = {{7'd0}, T_889};
  assign T_890 = T_886 | GEN_78;
  assign T_892 = cyc_C1_div ? sigB_PC : 53'h0;
  assign T_893 = T_890 | T_892;
  assign GEN_79 = {{1'd0}, T_893};
  assign T_894 = GEN_79 | zComplSigT_C1_sqrt;
  assign T_896 = T_858 | cyc_B6_sqrt;
  assign T_897 = T_896 | cyc_B4;
  assign T_898 = T_897 | cyc_C6_sqrt;
  assign T_899 = T_898 | cyc_C4;
  assign T_900 = T_899 | cyc_C1;
  assign GEN_80 = {{36'd0}, r1_A1};
  assign T_901 = GEN_80 << 36;
  assign T_903 = cyc_A1 ? T_901 : 52'h0;
  assign GEN_81 = {{19'd0}, ESqrR1_B_sqrt};
  assign T_904 = GEN_81 << 19;
  assign T_906 = cyc_B7_sqrt ? T_904 : 51'h0;
  assign GEN_82 = {{1'd0}, T_906};
  assign T_907 = T_903 | GEN_82;
  assign GEN_83 = {{36'd0}, ER1_B_sqrt};
  assign T_908 = GEN_83 << 36;
  assign T_910 = cyc_B6_sqrt ? T_908 : 53'h0;
  assign GEN_84 = {{1'd0}, T_907};
  assign T_911 = GEN_84 | T_910;
  assign GEN_85 = {{7'd0}, zSigma1_B4};
  assign T_912 = T_911 | GEN_85;
  assign T_913 = sqrSigma1_C[30:1];
  assign T_915 = cyc_C6_sqrt ? T_913 : 30'h0;
  assign GEN_86 = {{23'd0}, T_915};
  assign T_916 = T_912 | GEN_86;
  assign T_918 = cyc_C4 ? sqrSigma1_C : 33'h0;
  assign GEN_87 = {{20'd0}, T_918};
  assign T_919 = T_916 | GEN_87;
  assign GEN_88 = {{1'd0}, T_919};
  assign T_920 = GEN_88 | zComplSigT_C1;
  assign T_921 = cyc_A4 | cyc_A3_div;
  assign T_922 = T_921 | cyc_A1_div;
  assign T_923 = T_922 | cyc_B10_sqrt;
  assign T_924 = T_923 | cyc_B9_sqrt;
  assign T_925 = T_924 | cyc_B7_sqrt;
  assign T_926 = T_925 | cyc_B6;
  assign T_927 = T_926 | cyc_B5_sqrt;
  assign T_928 = T_927 | cyc_B3_sqrt;
  assign T_929 = T_928 | cyc_B2_div;
  assign T_930 = T_929 | cyc_B1_sqrt;
  assign T_931 = T_930 | cyc_C4;
  assign T_932 = cyc_A3 | cyc_A2_div;
  assign T_933 = T_932 | cyc_B9_sqrt;
  assign T_934 = T_933 | cyc_B8_sqrt;
  assign T_935 = T_934 | cyc_B6;
  assign T_936 = T_935 | cyc_B5;
  assign T_937 = T_936 | cyc_B4_sqrt;
  assign T_938 = T_937 | cyc_B2_sqrt;
  assign T_939 = T_938 | cyc_B1_div;
  assign T_940 = T_939 | cyc_C6_sqrt;
  assign T_941 = T_940 | valid_normalCase_leaving_PB;
  assign T_942 = cyc_A2 | cyc_A1_div;
  assign T_943 = T_942 | cyc_B8_sqrt;
  assign T_944 = T_943 | cyc_B7_sqrt;
  assign T_945 = T_944 | cyc_B5;
  assign T_946 = T_945 | cyc_B4;
  assign T_947 = T_946 | cyc_B3_sqrt;
  assign T_948 = T_947 | cyc_B1_sqrt;
  assign T_949 = T_948 | cyc_C5;
  assign T_950 = T_949 | cyc_C2;
  assign T_951 = io_latchMulAddA_0 | cyc_B6;
  assign T_952 = T_951 | cyc_B2_sqrt;
  assign T_953 = {T_950,T_952};
  assign T_954 = {T_931,T_941};
  assign T_955 = {T_954,T_953};
  assign GEN_89 = {{47'd0}, sigX1_B};
  assign T_956 = GEN_89 << 47;
  assign T_958 = cyc_B1 ? T_956 : 105'h0;
  assign GEN_90 = {{46'd0}, sigX1_B};
  assign T_959 = GEN_90 << 46;
  assign T_961 = cyc_C6_sqrt ? T_959 : 104'h0;
  assign GEN_91 = {{1'd0}, T_961};
  assign T_962 = T_958 | GEN_91;
  assign T_963 = cyc_C4_sqrt | cyc_C2;
  assign GEN_92 = {{47'd0}, sigXN_C};
  assign T_964 = GEN_92 << 47;
  assign T_966 = T_963 ? T_964 : 105'h0;
  assign T_967 = T_962 | T_966;
  assign T_969 = E_E_div == 1'h0;
  assign T_970 = cyc_E3_div & T_969;
  assign GEN_93 = {{53'd0}, fractA_0_PC};
  assign T_971 = GEN_93 << 53;
  assign T_973 = T_970 ? T_971 : 54'h0;
  assign GEN_94 = {{51'd0}, T_973};
  assign T_974 = T_967 | GEN_94;
  assign T_976 = sigB_PC[0];
  assign T_978 = {T_976,1'h0};
  assign T_979 = sigB_PC[1];
  assign T_981 = T_979 ^ T_976;
  assign T_983 = {T_981,T_976};
  assign T_984 = T_352 ? T_978 : T_983;
  assign T_986 = extraT_E == 1'h0;
  assign T_988 = {T_986,1'h0};
  assign T_989 = T_984 ^ T_988;
  assign GEN_95 = {{54'd0}, T_989};
  assign T_990 = GEN_95 << 54;
  assign T_992 = cyc_E3_sqrt ? T_990 : 56'h0;
  assign GEN_96 = {{49'd0}, T_992};
  assign T_993 = T_974 | GEN_96;
  assign ESqrR1_B8_sqrt = io_mulAddResult_3[103:72];
  assign T_994 = io_mulAddResult_3[90:45];
  assign T_995 = ~ T_994;
  assign T_997 = cyc_B4 ? T_995 : 46'h0;
  assign sqrSigma1_B1 = io_mulAddResult_3[79:47];
  assign T_998 = io_mulAddResult_3[104:47];
  assign T_999 = io_mulAddResult_3[104];
  assign E_C1_div = T_999 == 1'h0;
  assign T_1002 = E_C1_div == 1'h0;
  assign T_1003 = cyc_C1_div & T_1002;
  assign T_1004 = T_1003 | cyc_C1_sqrt;
  assign T_1005 = io_mulAddResult_3[104:51];
  assign T_1006 = ~ T_1005;
  assign T_1008 = T_1004 ? T_1006 : 54'h0;
  assign T_1009 = cyc_C1_div & E_C1_div;
  assign T_1011 = io_mulAddResult_3[102:50];
  assign T_1012 = ~ T_1011;
  assign T_1013 = {1'h0,T_1012};
  assign T_1015 = T_1009 ? T_1013 : 54'h0;
  assign T_1016 = T_1008 | T_1015;
  assign T_1020 = cyc_C1_sqrt ? T_1006 : 54'h0;
  assign sigT_C1 = ~ zComplSigT_C1;
  assign remT_E2 = io_mulAddResult_3[55:0];
  assign GEN_43 = cyc_B8_sqrt ? ESqrR1_B8_sqrt : ESqrR1_B_sqrt;
  assign GEN_44 = cyc_B3 ? sigXNU_B3_CX : sigX1_B;
  assign GEN_45 = cyc_B1 ? sqrSigma1_B1 : sqrSigma1_C;
  assign T_1021 = cyc_C6_sqrt | cyc_C5_div;
  assign T_1022 = T_1021 | cyc_C3_sqrt;
  assign GEN_46 = T_1022 ? sigXNU_B3_CX : sigXN_C;
  assign T_1023 = sigXNU_B3_CX[56:26];
  assign GEN_47 = cyc_C5_sqrt ? T_1023 : u_C_sqrt;
  assign T_1024 = sigT_C1[53:1];
  assign T_1025 = sigT_C1[0];
  assign GEN_48 = cyc_C1 ? E_C1_div : E_E_div;
  assign GEN_49 = cyc_C1 ? T_1024 : sigT_E;
  assign GEN_50 = cyc_C1 ? T_1025 : extraT_E;
  assign T_1026 = remT_E2[55];
  assign T_1027 = remT_E2[53];
  assign T_1028 = sqrtOp_PC ? T_1026 : T_1027;
  assign T_1029 = remT_E2[53:0];
  assign T_1031 = T_1029 == 54'h0;
  assign T_1034 = remT_E2[55:54];
  assign T_1036 = T_1034 == 2'h0;
  assign T_1037 = T_370 | T_1036;
  assign T_1038 = T_1031 & T_1037;
  assign GEN_51 = cyc_E2 ? T_1028 : isNegRemT_E;
  assign GEN_52 = cyc_E2 ? T_1038 : trueEqX_E1;
  assign T_1041 = T_370 & E_E_div;
  assign T_1043 = T_1041 ? exp_PC : 14'h0;
  assign T_1048 = T_370 & T_969;
  assign T_1050 = T_1048 ? expP1_PC : 14'h0;
  assign T_1051 = T_1043 | T_1050;
  assign T_1052 = exp_PC[13:1];
  assign T_1054 = T_1052 + 13'h400;
  assign T_1055 = T_1054[12:0];
  assign T_1057 = sqrtOp_PC ? T_1055 : 13'h0;
  assign GEN_97 = {{1'd0}, T_1057};
  assign sExpX_E = T_1051 | GEN_97;
  assign posExpX_E = sExpX_E[12:0];
  assign T_1058 = ~ posExpX_E;
  assign T_1059 = T_1058[12];
  assign T_1060 = T_1058[11:0];
  assign T_1061 = T_1060[11];
  assign T_1062 = T_1060[10:0];
  assign T_1063 = T_1062[10];
  assign T_1064 = T_1062[9:0];
  assign T_1065 = T_1064[9];
  assign T_1066 = T_1064[8:0];
  assign T_1068 = T_1066[8];
  assign T_1069 = T_1066[7:0];
  assign T_1071 = T_1069[7];
  assign T_1072 = T_1069[6:0];
  assign T_1074 = T_1072[6];
  assign T_1075 = T_1072[5:0];
  assign T_1078 = $signed(65'sh10000000000000000) >>> T_1075;
  assign T_1079 = T_1078[63:14];
  assign T_1080 = T_1079[31:0];
  assign T_1085 = T_1080[31:16];
  assign T_1086 = {{16'd0}, T_1085};
  assign T_1087 = T_1080[15:0];
  assign GEN_98 = {{16'd0}, T_1087};
  assign T_1088 = GEN_98 << 16;
  assign T_1090 = T_1088 & 32'hffff0000;
  assign T_1091 = T_1086 | T_1090;
  assign T_1095 = T_1091[31:8];
  assign GEN_99 = {{8'd0}, T_1095};
  assign T_1096 = GEN_99 & 32'hff00ff;
  assign T_1097 = T_1091[23:0];
  assign GEN_100 = {{8'd0}, T_1097};
  assign T_1098 = GEN_100 << 8;
  assign T_1100 = T_1098 & 32'hff00ff00;
  assign T_1101 = T_1096 | T_1100;
  assign T_1105 = T_1101[31:4];
  assign GEN_101 = {{4'd0}, T_1105};
  assign T_1106 = GEN_101 & 32'hf0f0f0f;
  assign T_1107 = T_1101[27:0];
  assign GEN_102 = {{4'd0}, T_1107};
  assign T_1108 = GEN_102 << 4;
  assign T_1110 = T_1108 & 32'hf0f0f0f0;
  assign T_1111 = T_1106 | T_1110;
  assign T_1115 = T_1111[31:2];
  assign GEN_103 = {{2'd0}, T_1115};
  assign T_1116 = GEN_103 & 32'h33333333;
  assign T_1117 = T_1111[29:0];
  assign GEN_104 = {{2'd0}, T_1117};
  assign T_1118 = GEN_104 << 2;
  assign T_1120 = T_1118 & 32'hcccccccc;
  assign T_1121 = T_1116 | T_1120;
  assign T_1125 = T_1121[31:1];
  assign GEN_105 = {{1'd0}, T_1125};
  assign T_1126 = GEN_105 & 32'h55555555;
  assign T_1127 = T_1121[30:0];
  assign GEN_106 = {{1'd0}, T_1127};
  assign T_1128 = GEN_106 << 1;
  assign T_1130 = T_1128 & 32'haaaaaaaa;
  assign T_1131 = T_1126 | T_1130;
  assign T_1132 = T_1079[49:32];
  assign T_1133 = T_1132[15:0];
  assign T_1138 = T_1133[15:8];
  assign T_1139 = {{8'd0}, T_1138};
  assign T_1140 = T_1133[7:0];
  assign GEN_107 = {{8'd0}, T_1140};
  assign T_1141 = GEN_107 << 8;
  assign T_1143 = T_1141 & 16'hff00;
  assign T_1144 = T_1139 | T_1143;
  assign T_1148 = T_1144[15:4];
  assign GEN_108 = {{4'd0}, T_1148};
  assign T_1149 = GEN_108 & 16'hf0f;
  assign T_1150 = T_1144[11:0];
  assign GEN_109 = {{4'd0}, T_1150};
  assign T_1151 = GEN_109 << 4;
  assign T_1153 = T_1151 & 16'hf0f0;
  assign T_1154 = T_1149 | T_1153;
  assign T_1158 = T_1154[15:2];
  assign GEN_110 = {{2'd0}, T_1158};
  assign T_1159 = GEN_110 & 16'h3333;
  assign T_1160 = T_1154[13:0];
  assign GEN_111 = {{2'd0}, T_1160};
  assign T_1161 = GEN_111 << 2;
  assign T_1163 = T_1161 & 16'hcccc;
  assign T_1164 = T_1159 | T_1163;
  assign T_1168 = T_1164[15:1];
  assign GEN_112 = {{1'd0}, T_1168};
  assign T_1169 = GEN_112 & 16'h5555;
  assign T_1170 = T_1164[14:0];
  assign GEN_113 = {{1'd0}, T_1170};
  assign T_1171 = GEN_113 << 1;
  assign T_1173 = T_1171 & 16'haaaa;
  assign T_1174 = T_1169 | T_1173;
  assign T_1175 = T_1132[17:16];
  assign T_1176 = T_1175[0];
  assign T_1177 = T_1175[1];
  assign T_1178 = {T_1176,T_1177};
  assign T_1179 = {T_1174,T_1178};
  assign T_1180 = {T_1131,T_1179};
  assign T_1181 = ~ T_1180;
  assign T_1182 = T_1074 ? 50'h0 : T_1181;
  assign T_1183 = ~ T_1182;
  assign T_1184 = ~ T_1183;
  assign T_1185 = T_1071 ? 50'h0 : T_1184;
  assign T_1186 = ~ T_1185;
  assign T_1187 = ~ T_1186;
  assign T_1188 = T_1068 ? 50'h0 : T_1187;
  assign T_1189 = ~ T_1188;
  assign T_1190 = ~ T_1189;
  assign T_1191 = T_1065 ? 50'h0 : T_1190;
  assign T_1192 = ~ T_1191;
  assign T_1194 = {T_1192,3'h7};
  assign T_1205 = T_1078[2:0];
  assign T_1206 = T_1205[1:0];
  assign T_1207 = T_1206[0];
  assign T_1208 = T_1206[1];
  assign T_1209 = {T_1207,T_1208};
  assign T_1210 = T_1205[2];
  assign T_1211 = {T_1209,T_1210};
  assign T_1213 = T_1074 ? T_1211 : 3'h0;
  assign T_1215 = T_1071 ? T_1213 : 3'h0;
  assign T_1217 = T_1068 ? T_1215 : 3'h0;
  assign T_1219 = T_1065 ? T_1217 : 3'h0;
  assign T_1220 = T_1063 ? T_1194 : {{50'd0}, T_1219};
  assign T_1222 = T_1061 ? T_1220 : 53'h0;
  assign roundMask_E = T_1059 ? T_1222 : 53'h0;
  assign T_1225 = {1'h0,roundMask_E};
  assign T_1226 = ~ T_1225;
  assign T_1228 = {roundMask_E,1'h1};
  assign incrPosMask_E = T_1226 & T_1228;
  assign T_1229 = incrPosMask_E[53:1];
  assign T_1230 = sigT_E & T_1229;
  assign hiRoundPosBitT_E = T_1230 != 53'h0;
  assign T_1232 = roundMask_E[52:1];
  assign GEN_114 = {{1'd0}, T_1232};
  assign T_1235 = ~ sigT_E;
  assign T_1237 = T_1235 & GEN_114;
  assign all1sHiRoundExtraT_E = T_1237 == 53'h0;
  assign T_1239 = roundMask_E[0];
  assign T_1241 = T_1239 == 1'h0;
  assign T_1242 = T_1241 | hiRoundPosBitT_E;
  assign all1sHiRoundT_E = T_1242 & all1sHiRoundExtraT_E;
  assign GEN_116 = {{1'd0}, sigT_E};
  assign T_1244 = 54'h0 + GEN_116;
  assign T_1245 = T_1244[53:0];
  assign GEN_117 = {{53'd0}, roundMagUp_PC};
  assign T_1246 = T_1245 + GEN_117;
  assign sigAdjT_E = T_1246[53:0];
  assign T_1248 = ~ roundMask_E;
  assign T_1249 = {1'h1,T_1248};
  assign sigY0_E = sigAdjT_E & T_1249;
  assign T_1252 = sigAdjT_E | T_1225;
  assign T_1254 = T_1252 + 54'h1;
  assign sigY1_E = T_1254[53:0];
  assign T_1256 = isNegRemT_E == 1'h0;
  assign T_1258 = trueEqX_E1 == 1'h0;
  assign T_1259 = T_1256 & T_1258;
  assign trueLtX_E1 = sqrtOp_PC ? T_1259 : isNegRemT_E;
  assign T_1262 = trueLtX_E1 == 1'h0;
  assign T_1263 = T_1239 & T_1262;
  assign T_1264 = T_1263 & all1sHiRoundExtraT_E;
  assign T_1265 = T_1264 & extraT_E;
  assign hiRoundPosBit_E1 = hiRoundPosBitT_E ^ T_1265;
  assign T_1270 = T_1258 | T_986;
  assign T_1272 = all1sHiRoundExtraT_E == 1'h0;
  assign anyRoundExtra_E1 = T_1270 | T_1272;
  assign T_1273 = roundingMode_near_even_PC & hiRoundPosBit_E1;
  assign T_1275 = anyRoundExtra_E1 == 1'h0;
  assign T_1276 = T_1273 & T_1275;
  assign roundEvenMask_E1 = T_1276 ? incrPosMask_E : 54'h0;
  assign T_1278 = roundMagDown_PC & extraT_E;
  assign T_1281 = T_1278 & T_1262;
  assign T_1282 = T_1281 & all1sHiRoundT_E;
  assign T_1285 = extraT_E & T_1262;
  assign T_1288 = T_1285 & T_1258;
  assign T_1290 = all1sHiRoundT_E == 1'h0;
  assign T_1291 = T_1288 | T_1290;
  assign T_1292 = roundMagUp_PC & T_1291;
  assign T_1293 = T_1282 | T_1292;
  assign T_1296 = extraT_E | T_1262;
  assign T_1300 = T_1296 & T_1241;
  assign T_1301 = hiRoundPosBitT_E | T_1300;
  assign T_1305 = T_1285 & all1sHiRoundExtraT_E;
  assign T_1306 = T_1301 | T_1305;
  assign T_1307 = roundingMode_near_even_PC & T_1306;
  assign T_1308 = T_1293 | T_1307;
  assign T_1309 = T_1308 ? sigY1_E : sigY0_E;
  assign T_1310 = ~ roundEvenMask_E1;
  assign sigY_E1 = T_1309 & T_1310;
  assign fractY_E1 = sigY_E1[51:0];
  assign inexactY_E1 = hiRoundPosBit_E1 | anyRoundExtra_E1;
  assign T_1311 = sigY_E1[53];
  assign T_1313 = T_1311 == 1'h0;
  assign T_1315 = T_1313 ? sExpX_E : 14'h0;
  assign T_1319 = T_1311 & T_370;
  assign T_1320 = T_1319 & E_E_div;
  assign T_1322 = T_1320 ? expP1_PC : 14'h0;
  assign T_1323 = T_1315 | T_1322;
  assign T_1330 = T_1319 & T_969;
  assign T_1332 = T_1330 ? expP2_PC : 14'h0;
  assign T_1333 = T_1323 | T_1332;
  assign T_1335 = T_1311 & sqrtOp_PC;
  assign T_1336 = expP2_PC[13:1];
  assign T_1338 = T_1336 + 13'h400;
  assign T_1339 = T_1338[12:0];
  assign T_1341 = T_1335 ? T_1339 : 13'h0;
  assign GEN_118 = {{1'd0}, T_1341};
  assign sExpY_E1 = T_1333 | GEN_118;
  assign expY_E1 = sExpY_E1[11:0];
  assign T_1342 = sExpY_E1[13];
  assign T_1344 = T_1342 == 1'h0;
  assign T_1346 = sExpY_E1[12:10];
  assign T_1347 = 3'h3 <= T_1346;
  assign overflowY_E1 = T_1344 & T_1347;
  assign T_1349 = sExpY_E1[12:0];
  assign T_1351 = T_1349 < 13'h3ce;
  assign totalUnderflowY_E1 = T_1342 | T_1351;
  assign T_1353 = posExpX_E <= 13'h401;
  assign T_1354 = T_1353 & inexactY_E1;
  assign underflowY_E1 = totalUnderflowY_E1 | T_1354;
  assign T_1356 = isNaNB_PC == 1'h0;
  assign T_1359 = T_1356 & T_334;
  assign T_1360 = T_1359 & sign_PC;
  assign T_1361 = isZeroA_PC & isZeroB_PC;
  assign T_1362 = isInfA_PC & isInfB_PC;
  assign T_1363 = T_1361 | T_1362;
  assign notSigNaN_invalid_PC = sqrtOp_PC ? T_1360 : T_1363;
  assign T_1366 = T_370 & isSigNaNA_PC;
  assign T_1367 = T_1366 | isSigNaNB_PC;
  assign invalid_PC = T_1367 | notSigNaN_invalid_PC;
  assign T_1372 = T_370 & T_340;
  assign T_1375 = T_1372 & T_345;
  assign infinity_PC = T_1375 & isZeroB_PC;
  assign overflow_E1 = normalCase_PC & overflowY_E1;
  assign underflow_E1 = normalCase_PC & underflowY_E1;
  assign T_1376 = overflow_E1 | underflow_E1;
  assign T_1377 = normalCase_PC & inexactY_E1;
  assign inexact_E1 = T_1376 | T_1377;
  assign T_1378 = isZeroA_PC | isInfB_PC;
  assign T_1381 = totalUnderflowY_E1 & T_360;
  assign T_1382 = T_1378 | T_1381;
  assign notSpecial_isZeroOut_E1 = sqrtOp_PC ? isZeroB_PC : T_1382;
  assign T_1383 = normalCase_PC & totalUnderflowY_E1;
  assign pegMinFiniteMagOut_E1 = T_1383 & roundMagUp_PC;
  assign T_1385 = overflowY_roundMagUp_PC == 1'h0;
  assign pegMaxFiniteMagOut_E1 = overflow_E1 & T_1385;
  assign T_1386 = isInfA_PC | isZeroB_PC;
  assign T_1387 = overflow_E1 & overflowY_roundMagUp_PC;
  assign T_1388 = T_1386 | T_1387;
  assign notNaN_isInfOut_E1 = sqrtOp_PC ? isInfB_PC : T_1388;
  assign T_1391 = T_370 & isNaNA_PC;
  assign T_1392 = T_1391 | isNaNB_PC;
  assign isNaNOut_PC = T_1392 | notSigNaN_invalid_PC;
  assign T_1394 = isNaNOut_PC == 1'h0;
  assign T_1395 = isZeroB_PC & sign_PC;
  assign T_1396 = sqrtOp_PC ? T_1395 : sign_PC;
  assign signOut_PC = T_1394 & T_1396;
  assign T_1400 = notSpecial_isZeroOut_E1 ? 12'he00 : 12'h0;
  assign T_1401 = ~ T_1400;
  assign T_1402 = expY_E1 & T_1401;
  assign T_1406 = pegMinFiniteMagOut_E1 ? 12'hc31 : 12'h0;
  assign T_1407 = ~ T_1406;
  assign T_1408 = T_1402 & T_1407;
  assign T_1412 = pegMaxFiniteMagOut_E1 ? 12'h400 : 12'h0;
  assign T_1413 = ~ T_1412;
  assign T_1414 = T_1408 & T_1413;
  assign T_1418 = notNaN_isInfOut_E1 ? 12'h200 : 12'h0;
  assign T_1419 = ~ T_1418;
  assign T_1420 = T_1414 & T_1419;
  assign T_1423 = pegMinFiniteMagOut_E1 ? 12'h3ce : 12'h0;
  assign T_1424 = T_1420 | T_1423;
  assign T_1427 = pegMaxFiniteMagOut_E1 ? 12'hbff : 12'h0;
  assign T_1428 = T_1424 | T_1427;
  assign T_1431 = notNaN_isInfOut_E1 ? 12'hc00 : 12'h0;
  assign T_1432 = T_1428 | T_1431;
  assign T_1435 = isNaNOut_PC ? 12'he00 : 12'h0;
  assign expOut_E1 = T_1432 | T_1435;
  assign T_1436 = notSpecial_isZeroOut_E1 | totalUnderflowY_E1;
  assign T_1437 = T_1436 | isNaNOut_PC;
  assign T_1441 = isNaNOut_PC ? 52'h8000000000000 : 52'h0;
  assign T_1442 = T_1437 ? T_1441 : fractY_E1;
  assign T_1446 = pegMaxFiniteMagOut_E1 ? 52'hfffffffffffff : 52'h0;
  assign fractOut_E1 = T_1442 | T_1446;
  assign T_1447 = {signOut_PC,expOut_E1};
  assign T_1448 = {T_1447,fractOut_E1};
  assign T_1449 = {underflow_E1,inexact_E1};
  assign T_1450 = {invalid_PC,infinity_PC};
  assign T_1451 = {T_1450,overflow_E1};
  assign T_1452 = {T_1451,T_1449};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  valid_PA = GEN_115[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  sqrtOp_PA = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  sign_PA = GEN_120[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {1{$random}};
  specialCodeB_PA = GEN_121[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_122 = {1{$random}};
  fractB_51_PA = GEN_122[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_123 = {1{$random}};
  roundingMode_PA = GEN_123[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_124 = {1{$random}};
  specialCodeA_PA = GEN_124[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  fractA_51_PA = GEN_125[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {1{$random}};
  exp_PA = GEN_126[13:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {2{$random}};
  fractB_other_PA = GEN_127[50:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {2{$random}};
  fractA_other_PA = GEN_128[50:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {1{$random}};
  valid_PB = GEN_129[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {1{$random}};
  sqrtOp_PB = GEN_130[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  sign_PB = GEN_131[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  specialCodeA_PB = GEN_132[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  fractA_51_PB = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  specialCodeB_PB = GEN_134[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  fractB_51_PB = GEN_135[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {1{$random}};
  roundingMode_PB = GEN_136[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  exp_PB = GEN_137[13:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  fractA_0_PB = GEN_138[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {2{$random}};
  fractB_other_PB = GEN_139[50:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  valid_PC = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  sqrtOp_PC = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  sign_PC = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  specialCodeA_PC = GEN_143[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  fractA_51_PC = GEN_144[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  specialCodeB_PC = GEN_145[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  fractB_51_PC = GEN_146[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  roundingMode_PC = GEN_147[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {1{$random}};
  exp_PC = GEN_148[13:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  fractA_0_PC = GEN_149[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {2{$random}};
  fractB_other_PC = GEN_150[50:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  cycleNum_A = GEN_151[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  cycleNum_B = GEN_152[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  cycleNum_C = GEN_153[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  cycleNum_E = GEN_154[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  fractR0_A = GEN_155[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  hiSqrR0_A_sqrt = GEN_156[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  partNegSigma0_A = GEN_157[20:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  nextMulAdd9A_A = GEN_158[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  nextMulAdd9B_A = GEN_159[8:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {1{$random}};
  ER1_B_sqrt = GEN_160[16:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  ESqrR1_B_sqrt = GEN_161[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {2{$random}};
  sigX1_B = GEN_162[57:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {2{$random}};
  sqrSigma1_C = GEN_163[32:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {2{$random}};
  sigXN_C = GEN_164[57:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {1{$random}};
  u_C_sqrt = GEN_165[30:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_166 = {1{$random}};
  E_E_div = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_167 = {2{$random}};
  sigT_E = GEN_167[52:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_168 = {1{$random}};
  extraT_E = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_169 = {1{$random}};
  isNegRemT_E = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_170 = {1{$random}};
  trueEqX_E1 = GEN_170[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      valid_PA <= 1'h0;
    end else begin
      if(T_207) begin
        valid_PA <= entering_PA;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA) begin
        sqrtOp_PA <= io_sqrtOp;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA) begin
        if(io_sqrtOp) begin
          sign_PA <= signB_S;
        end else begin
          sign_PA <= T_164;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA) begin
        specialCodeB_PA <= specialCodeB_S;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA) begin
        fractB_51_PA <= T_208;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA) begin
        roundingMode_PA <= io_roundingMode;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_211) begin
        specialCodeA_PA <= specialCodeA_S;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_211) begin
        fractA_51_PA <= T_212;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA_normalCase) begin
        if(io_sqrtOp) begin
          exp_PA <= {{2'd0}, expB_S};
        end else begin
          exp_PA <= T_222;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA_normalCase) begin
        fractB_other_PA <= T_224;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PA_normalCase_div) begin
        fractA_other_PA <= T_225;
      end
    end
    if(reset) begin
      valid_PB <= 1'h0;
    end else begin
      if(T_260) begin
        valid_PB <= entering_PB;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          sqrtOp_PB <= sqrtOp_PA;
        end else begin
          sqrtOp_PB <= io_sqrtOp;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          sign_PB <= sign_PA;
        end else begin
          if(io_sqrtOp) begin
            sign_PB <= signB_S;
          end else begin
            sign_PB <= T_164;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          specialCodeA_PB <= specialCodeA_PA;
        end else begin
          specialCodeA_PB <= specialCodeA_S;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          fractA_51_PB <= fractA_51_PA;
        end else begin
          fractA_51_PB <= T_212;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          specialCodeB_PB <= specialCodeB_PA;
        end else begin
          specialCodeB_PB <= specialCodeB_S;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          fractB_51_PB <= fractB_51_PA;
        end else begin
          fractB_51_PB <= T_208;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB) begin
        if(valid_PA) begin
          roundingMode_PB <= roundingMode_PA;
        end else begin
          roundingMode_PB <= io_roundingMode;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB_normalCase) begin
        exp_PB <= exp_PA;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB_normalCase) begin
        fractA_0_PB <= T_270;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PB_normalCase) begin
        fractB_other_PB <= fractB_other_PA;
      end
    end
    if(reset) begin
      valid_PC <= 1'h0;
    end else begin
      if(T_301) begin
        valid_PC <= entering_PC;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          sqrtOp_PC <= sqrtOp_PB;
        end else begin
          sqrtOp_PC <= io_sqrtOp;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          sign_PC <= sign_PB;
        end else begin
          if(io_sqrtOp) begin
            sign_PC <= signB_S;
          end else begin
            sign_PC <= T_164;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          specialCodeA_PC <= specialCodeA_PB;
        end else begin
          specialCodeA_PC <= specialCodeA_S;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          fractA_51_PC <= fractA_51_PB;
        end else begin
          fractA_51_PC <= T_212;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          specialCodeB_PC <= specialCodeB_PB;
        end else begin
          specialCodeB_PC <= specialCodeB_S;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          fractB_51_PC <= fractB_51_PB;
        end else begin
          fractB_51_PC <= T_208;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC) begin
        if(valid_PB) begin
          roundingMode_PC <= roundingMode_PB;
        end else begin
          roundingMode_PC <= io_roundingMode;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC_normalCase) begin
        exp_PC <= exp_PB;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC_normalCase) begin
        fractA_0_PC <= fractA_0_PB;
      end
    end
    if(1'h0) begin
    end else begin
      if(entering_PC_normalCase) begin
        fractB_other_PC <= fractB_other_PB;
      end
    end
    if(reset) begin
      cycleNum_A <= 3'h0;
    end else begin
      if(T_375) begin
        cycleNum_A <= T_390;
      end
    end
    if(reset) begin
      cycleNum_B <= 4'h0;
    end else begin
      if(T_405) begin
        if(cyc_A1) begin
          if(sqrtOp_PA) begin
            cycleNum_B <= 4'ha;
          end else begin
            cycleNum_B <= 4'h6;
          end
        end else begin
          cycleNum_B <= T_411;
        end
      end
    end
    if(reset) begin
      cycleNum_C <= 3'h0;
    end else begin
      if(T_465) begin
        if(cyc_B1) begin
          if(sqrtOp_PB) begin
            cycleNum_C <= 3'h6;
          end else begin
            cycleNum_C <= 3'h5;
          end
        end else begin
          cycleNum_C <= T_471;
        end
      end
    end
    if(reset) begin
      cycleNum_E <= 3'h0;
    end else begin
      if(T_496) begin
        if(cyc_C1) begin
          cycleNum_E <= 3'h4;
        end else begin
          cycleNum_E <= T_500;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_808) begin
        fractR0_A <= T_809;
      end
    end
    if(1'h0) begin
    end else begin
      hiSqrR0_A_sqrt <= GEN_38[9:0];
    end
    if(1'h0) begin
    end else begin
      if(T_811) begin
        partNegSigma0_A <= T_814;
      end
    end
    if(1'h0) begin
    end else begin
      nextMulAdd9A_A <= GEN_40[8:0];
    end
    if(1'h0) begin
    end else begin
      if(T_840) begin
        nextMulAdd9B_A <= T_857;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_A1_sqrt) begin
        if(T_664) begin
          ER1_B_sqrt <= T_807;
        end else begin
          ER1_B_sqrt <= {{1'd0}, r1_A1};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_B8_sqrt) begin
        ESqrR1_B_sqrt <= ESqrR1_B8_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_B3) begin
        sigX1_B <= sigXNU_B3_CX;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_B1) begin
        sqrSigma1_C <= sqrSigma1_B1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1022) begin
        sigXN_C <= sigXNU_B3_CX;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_C5_sqrt) begin
        u_C_sqrt <= T_1023;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_C1) begin
        E_E_div <= E_C1_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_C1) begin
        sigT_E <= T_1024;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_C1) begin
        extraT_E <= T_1025;
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_E2) begin
        if(sqrtOp_PC) begin
          isNegRemT_E <= T_1026;
        end else begin
          isNegRemT_E <= T_1027;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(cyc_E2) begin
        trueEqX_E1 <= T_1038;
      end
    end
  end
endmodule
module Mul54(
  input   clk,
  input   reset,
  input   io_val_s0,
  input   io_latch_a_s0,
  input  [53:0] io_a_s0,
  input   io_latch_b_s0,
  input  [53:0] io_b_s0,
  input  [104:0] io_c_s2,
  output [104:0] io_result_s3
);
  reg  val_s1;
  reg [31:0] GEN_7;
  reg  val_s2;
  reg [31:0] GEN_8;
  reg [53:0] reg_a_s1;
  reg [63:0] GEN_9;
  reg [53:0] reg_b_s1;
  reg [63:0] GEN_10;
  reg [53:0] reg_a_s2;
  reg [63:0] GEN_11;
  reg [53:0] reg_b_s2;
  reg [63:0] GEN_12;
  reg [104:0] reg_result_s3;
  reg [127:0] GEN_13;
  wire [53:0] GEN_0;
  wire [53:0] GEN_1;
  wire [53:0] GEN_2;
  wire [53:0] GEN_3;
  wire [53:0] GEN_4;
  wire [53:0] GEN_5;
  wire [107:0] T_14;
  wire [104:0] T_15;
  wire [105:0] T_16;
  wire [104:0] T_17;
  wire [104:0] GEN_6;
  assign io_result_s3 = reg_result_s3;
  assign GEN_0 = io_latch_a_s0 ? io_a_s0 : reg_a_s1;
  assign GEN_1 = io_latch_b_s0 ? io_b_s0 : reg_b_s1;
  assign GEN_2 = io_val_s0 ? GEN_0 : reg_a_s1;
  assign GEN_3 = io_val_s0 ? GEN_1 : reg_b_s1;
  assign GEN_4 = val_s1 ? reg_a_s1 : reg_a_s2;
  assign GEN_5 = val_s1 ? reg_b_s1 : reg_b_s2;
  assign T_14 = reg_a_s2 * reg_b_s2;
  assign T_15 = T_14[104:0];
  assign T_16 = T_15 + io_c_s2;
  assign T_17 = T_16[104:0];
  assign GEN_6 = val_s2 ? T_17 : reg_result_s3;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  val_s1 = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  val_s2 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {2{$random}};
  reg_a_s1 = GEN_9[53:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {2{$random}};
  reg_b_s1 = GEN_10[53:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {2{$random}};
  reg_a_s2 = GEN_11[53:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_12 = {2{$random}};
  reg_b_s2 = GEN_12[53:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_13 = {4{$random}};
  reg_result_s3 = GEN_13[104:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      val_s1 <= io_val_s0;
    end
    if(1'h0) begin
    end else begin
      val_s2 <= val_s1;
    end
    if(1'h0) begin
    end else begin
      if(io_val_s0) begin
        if(io_latch_a_s0) begin
          reg_a_s1 <= io_a_s0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_val_s0) begin
        if(io_latch_b_s0) begin
          reg_b_s1 <= io_b_s0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(val_s1) begin
        reg_a_s2 <= reg_a_s1;
      end
    end
    if(1'h0) begin
    end else begin
      if(val_s1) begin
        reg_b_s2 <= reg_b_s1;
      end
    end
    if(1'h0) begin
    end else begin
      if(val_s2) begin
        reg_result_s3 <= T_17;
      end
    end
  end
endmodule
module DivSqrtRecF64(
  input   clk,
  input   reset,
  output  io_inReady_div,
  output  io_inReady_sqrt,
  input   io_inValid,
  input   io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [1:0] io_roundingMode,
  output  io_outValid_div,
  output  io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  ds_clk;
  wire  ds_reset;
  wire  ds_io_inReady_div;
  wire  ds_io_inReady_sqrt;
  wire  ds_io_inValid;
  wire  ds_io_sqrtOp;
  wire [64:0] ds_io_a;
  wire [64:0] ds_io_b;
  wire [1:0] ds_io_roundingMode;
  wire  ds_io_outValid_div;
  wire  ds_io_outValid_sqrt;
  wire [64:0] ds_io_out;
  wire [4:0] ds_io_exceptionFlags;
  wire [3:0] ds_io_usingMulAdd;
  wire  ds_io_latchMulAddA_0;
  wire [53:0] ds_io_mulAddA_0;
  wire  ds_io_latchMulAddB_0;
  wire [53:0] ds_io_mulAddB_0;
  wire [104:0] ds_io_mulAddC_2;
  wire [104:0] ds_io_mulAddResult_3;
  wire  mul_clk;
  wire  mul_reset;
  wire  mul_io_val_s0;
  wire  mul_io_latch_a_s0;
  wire [53:0] mul_io_a_s0;
  wire  mul_io_latch_b_s0;
  wire [53:0] mul_io_b_s0;
  wire [104:0] mul_io_c_s2;
  wire [104:0] mul_io_result_s3;
  wire  T_11;
  DivSqrtRecF64_mulAddZ31 ds (
    .clk(ds_clk),
    .reset(ds_reset),
    .io_inReady_div(ds_io_inReady_div),
    .io_inReady_sqrt(ds_io_inReady_sqrt),
    .io_inValid(ds_io_inValid),
    .io_sqrtOp(ds_io_sqrtOp),
    .io_a(ds_io_a),
    .io_b(ds_io_b),
    .io_roundingMode(ds_io_roundingMode),
    .io_outValid_div(ds_io_outValid_div),
    .io_outValid_sqrt(ds_io_outValid_sqrt),
    .io_out(ds_io_out),
    .io_exceptionFlags(ds_io_exceptionFlags),
    .io_usingMulAdd(ds_io_usingMulAdd),
    .io_latchMulAddA_0(ds_io_latchMulAddA_0),
    .io_mulAddA_0(ds_io_mulAddA_0),
    .io_latchMulAddB_0(ds_io_latchMulAddB_0),
    .io_mulAddB_0(ds_io_mulAddB_0),
    .io_mulAddC_2(ds_io_mulAddC_2),
    .io_mulAddResult_3(ds_io_mulAddResult_3)
  );
  Mul54 mul (
    .clk(mul_clk),
    .reset(mul_reset),
    .io_val_s0(mul_io_val_s0),
    .io_latch_a_s0(mul_io_latch_a_s0),
    .io_a_s0(mul_io_a_s0),
    .io_latch_b_s0(mul_io_latch_b_s0),
    .io_b_s0(mul_io_b_s0),
    .io_c_s2(mul_io_c_s2),
    .io_result_s3(mul_io_result_s3)
  );
  assign io_inReady_div = ds_io_inReady_div;
  assign io_inReady_sqrt = ds_io_inReady_sqrt;
  assign io_outValid_div = ds_io_outValid_div;
  assign io_outValid_sqrt = ds_io_outValid_sqrt;
  assign io_out = ds_io_out;
  assign io_exceptionFlags = ds_io_exceptionFlags;
  assign ds_clk = clk;
  assign ds_reset = reset;
  assign ds_io_inValid = io_inValid;
  assign ds_io_sqrtOp = io_sqrtOp;
  assign ds_io_a = io_a;
  assign ds_io_b = io_b;
  assign ds_io_roundingMode = io_roundingMode;
  assign ds_io_mulAddResult_3 = mul_io_result_s3;
  assign mul_clk = clk;
  assign mul_reset = reset;
  assign mul_io_val_s0 = T_11;
  assign mul_io_latch_a_s0 = ds_io_latchMulAddA_0;
  assign mul_io_a_s0 = ds_io_mulAddA_0;
  assign mul_io_latch_b_s0 = ds_io_latchMulAddB_0;
  assign mul_io_b_s0 = ds_io_mulAddB_0;
  assign mul_io_c_s2 = ds_io_mulAddC_2;
  assign T_11 = ds_io_usingMulAdd[0];
endmodule
module RecFNToRecFN_2(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_4;
  wire [2:0] T_5;
  wire  T_7;
  wire [1:0] T_8;
  wire  T_10;
  wire  T_18_sign;
  wire  T_18_isNaN;
  wire  T_18_isInf;
  wire  T_18_isZero;
  wire [12:0] T_18_sExp;
  wire [55:0] T_18_sig;
  wire  T_25;
  wire  T_26;
  wire  T_27;
  wire  T_30;
  wire  T_31;
  wire [12:0] T_32;
  wire  T_35;
  wire [51:0] T_36;
  wire [53:0] T_38;
  wire [1:0] T_39;
  wire [55:0] T_40;
  wire [13:0] T_42;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [9:0] outRawFloat_sExp;
  wire [26:0] outRawFloat_sig;
  wire  T_57;
  wire [3:0] T_58;
  wire  T_60;
  wire [8:0] T_68;
  wire [8:0] T_69;
  wire [9:0] T_70;
  wire [9:0] T_71;
  wire [25:0] T_72;
  wire [29:0] T_73;
  wire  T_75;
  wire [26:0] T_76;
  wire  T_77;
  wire  T_79;
  wire  invalidExc;
  wire  RoundRawFNToRecFN_1_1_clk;
  wire  RoundRawFNToRecFN_1_1_reset;
  wire  RoundRawFNToRecFN_1_1_io_invalidExc;
  wire  RoundRawFNToRecFN_1_1_io_infiniteExc;
  wire  RoundRawFNToRecFN_1_1_io_in_sign;
  wire  RoundRawFNToRecFN_1_1_io_in_isNaN;
  wire  RoundRawFNToRecFN_1_1_io_in_isInf;
  wire  RoundRawFNToRecFN_1_1_io_in_isZero;
  wire [9:0] RoundRawFNToRecFN_1_1_io_in_sExp;
  wire [26:0] RoundRawFNToRecFN_1_1_io_in_sig;
  wire [1:0] RoundRawFNToRecFN_1_1_io_roundingMode;
  wire [32:0] RoundRawFNToRecFN_1_1_io_out;
  wire [4:0] RoundRawFNToRecFN_1_1_io_exceptionFlags;
  RoundRawFNToRecFN RoundRawFNToRecFN_1_1 (
    .clk(RoundRawFNToRecFN_1_1_clk),
    .reset(RoundRawFNToRecFN_1_1_reset),
    .io_invalidExc(RoundRawFNToRecFN_1_1_io_invalidExc),
    .io_infiniteExc(RoundRawFNToRecFN_1_1_io_infiniteExc),
    .io_in_sign(RoundRawFNToRecFN_1_1_io_in_sign),
    .io_in_isNaN(RoundRawFNToRecFN_1_1_io_in_isNaN),
    .io_in_isInf(RoundRawFNToRecFN_1_1_io_in_isInf),
    .io_in_isZero(RoundRawFNToRecFN_1_1_io_in_isZero),
    .io_in_sExp(RoundRawFNToRecFN_1_1_io_in_sExp),
    .io_in_sig(RoundRawFNToRecFN_1_1_io_in_sig),
    .io_roundingMode(RoundRawFNToRecFN_1_1_io_roundingMode),
    .io_out(RoundRawFNToRecFN_1_1_io_out),
    .io_exceptionFlags(RoundRawFNToRecFN_1_1_io_exceptionFlags)
  );
  assign io_out = RoundRawFNToRecFN_1_1_io_out;
  assign io_exceptionFlags = RoundRawFNToRecFN_1_1_io_exceptionFlags;
  assign T_4 = io_in[63:52];
  assign T_5 = T_4[11:9];
  assign T_7 = T_5 == 3'h0;
  assign T_8 = T_4[11:10];
  assign T_10 = T_8 == 2'h3;
  assign T_18_sign = T_25;
  assign T_18_isNaN = T_27;
  assign T_18_isInf = T_31;
  assign T_18_isZero = T_7;
  assign T_18_sExp = T_32;
  assign T_18_sig = T_40;
  assign T_25 = io_in[64];
  assign T_26 = T_4[9];
  assign T_27 = T_10 & T_26;
  assign T_30 = T_26 == 1'h0;
  assign T_31 = T_10 & T_30;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_35 = T_7 == 1'h0;
  assign T_36 = io_in[51:0];
  assign T_38 = {T_36,2'h0};
  assign T_39 = {1'h0,T_35};
  assign T_40 = {T_39,T_38};
  assign T_42 = $signed(T_18_sExp) + $signed(13'sh1900);
  assign outRawFloat_sign = T_18_sign;
  assign outRawFloat_isNaN = T_18_isNaN;
  assign outRawFloat_isInf = T_18_isInf;
  assign outRawFloat_isZero = T_18_isZero;
  assign outRawFloat_sExp = T_71;
  assign outRawFloat_sig = T_76;
  assign T_57 = $signed(T_42) < $signed(14'sh0);
  assign T_58 = T_42[12:9];
  assign T_60 = T_58 != 4'h0;
  assign T_68 = T_42[8:0];
  assign T_69 = T_60 ? 9'h1fc : T_68;
  assign T_70 = {T_57,T_69};
  assign T_71 = $signed(T_70);
  assign T_72 = T_18_sig[55:30];
  assign T_73 = T_18_sig[29:0];
  assign T_75 = T_73 != 30'h0;
  assign T_76 = {T_72,T_75};
  assign T_77 = outRawFloat_sig[24];
  assign T_79 = T_77 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_79;
  assign RoundRawFNToRecFN_1_1_clk = clk;
  assign RoundRawFNToRecFN_1_1_reset = reset;
  assign RoundRawFNToRecFN_1_1_io_invalidExc = invalidExc;
  assign RoundRawFNToRecFN_1_1_io_infiniteExc = 1'h0;
  assign RoundRawFNToRecFN_1_1_io_in_sign = outRawFloat_sign;
  assign RoundRawFNToRecFN_1_1_io_in_isNaN = outRawFloat_isNaN;
  assign RoundRawFNToRecFN_1_1_io_in_isInf = outRawFloat_isInf;
  assign RoundRawFNToRecFN_1_1_io_in_isZero = outRawFloat_isZero;
  assign RoundRawFNToRecFN_1_1_io_in_sExp = outRawFloat_sExp;
  assign RoundRawFNToRecFN_1_1_io_in_sig = outRawFloat_sig;
  assign RoundRawFNToRecFN_1_1_io_roundingMode = io_roundingMode;
endmodule
module FPU(
  input   clk,
  input   reset,
  input  [31:0] io_inst,
  input  [63:0] io_fromint_data,
  input  [2:0] io_fcsr_rm,
  output  io_fcsr_flags_valid,
  output [4:0] io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input   io_dmem_resp_val,
  input  [2:0] io_dmem_resp_type,
  input  [4:0] io_dmem_resp_tag,
  input  [63:0] io_dmem_resp_data,
  input   io_valid,
  output  io_fcsr_rdy,
  output  io_nack_mem,
  output  io_illegal_rm,
  input   io_killx,
  input   io_killm,
  output [4:0] io_dec_cmd,
  output  io_dec_ldst,
  output  io_dec_wen,
  output  io_dec_ren1,
  output  io_dec_ren2,
  output  io_dec_ren3,
  output  io_dec_swap12,
  output  io_dec_swap23,
  output  io_dec_single,
  output  io_dec_fromint,
  output  io_dec_toint,
  output  io_dec_fastpipe,
  output  io_dec_fma,
  output  io_dec_div,
  output  io_dec_sqrt,
  output  io_dec_round,
  output  io_dec_wflags,
  output  io_sboard_set,
  output  io_sboard_clr,
  output [4:0] io_sboard_clra,
  output  io_cp_req_ready,
  input   io_cp_req_valid,
  input  [4:0] io_cp_req_bits_cmd,
  input   io_cp_req_bits_ldst,
  input   io_cp_req_bits_wen,
  input   io_cp_req_bits_ren1,
  input   io_cp_req_bits_ren2,
  input   io_cp_req_bits_ren3,
  input   io_cp_req_bits_swap12,
  input   io_cp_req_bits_swap23,
  input   io_cp_req_bits_single,
  input   io_cp_req_bits_fromint,
  input   io_cp_req_bits_toint,
  input   io_cp_req_bits_fastpipe,
  input   io_cp_req_bits_fma,
  input   io_cp_req_bits_div,
  input   io_cp_req_bits_sqrt,
  input   io_cp_req_bits_round,
  input   io_cp_req_bits_wflags,
  input  [2:0] io_cp_req_bits_rm,
  input  [1:0] io_cp_req_bits_typ,
  input  [64:0] io_cp_req_bits_in1,
  input  [64:0] io_cp_req_bits_in2,
  input  [64:0] io_cp_req_bits_in3,
  input   io_cp_resp_ready,
  output  io_cp_resp_valid,
  output [64:0] io_cp_resp_bits_data,
  output [4:0] io_cp_resp_bits_exc
);
  reg  ex_reg_valid;
  reg [31:0] GEN_57;
  wire  req_valid;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_58;
  wire [31:0] GEN_0;
  wire  ex_cp_valid;
  wire  T_194;
  wire  T_195;
  wire  T_196;
  reg  mem_reg_valid;
  reg [31:0] GEN_59;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_60;
  wire [31:0] GEN_1;
  reg  mem_cp_valid;
  reg [31:0] GEN_100;
  wire  T_199;
  wire  T_201;
  wire  killm;
  wire  T_203;
  wire  T_204;
  wire  T_205;
  reg  wb_reg_valid;
  reg [31:0] GEN_124;
  reg  wb_cp_valid;
  reg [31:0] GEN_125;
  wire  fp_decoder_clk;
  wire  fp_decoder_reset;
  wire [31:0] fp_decoder_io_inst;
  wire [4:0] fp_decoder_io_sigs_cmd;
  wire  fp_decoder_io_sigs_ldst;
  wire  fp_decoder_io_sigs_wen;
  wire  fp_decoder_io_sigs_ren1;
  wire  fp_decoder_io_sigs_ren2;
  wire  fp_decoder_io_sigs_ren3;
  wire  fp_decoder_io_sigs_swap12;
  wire  fp_decoder_io_sigs_swap23;
  wire  fp_decoder_io_sigs_single;
  wire  fp_decoder_io_sigs_fromint;
  wire  fp_decoder_io_sigs_toint;
  wire  fp_decoder_io_sigs_fastpipe;
  wire  fp_decoder_io_sigs_fma;
  wire  fp_decoder_io_sigs_div;
  wire  fp_decoder_io_sigs_sqrt;
  wire  fp_decoder_io_sigs_round;
  wire  fp_decoder_io_sigs_wflags;
  wire [4:0] cp_ctrl_cmd;
  wire  cp_ctrl_ldst;
  wire  cp_ctrl_wen;
  wire  cp_ctrl_ren1;
  wire  cp_ctrl_ren2;
  wire  cp_ctrl_ren3;
  wire  cp_ctrl_swap12;
  wire  cp_ctrl_swap23;
  wire  cp_ctrl_single;
  wire  cp_ctrl_fromint;
  wire  cp_ctrl_toint;
  wire  cp_ctrl_fastpipe;
  wire  cp_ctrl_fma;
  wire  cp_ctrl_div;
  wire  cp_ctrl_sqrt;
  wire  cp_ctrl_round;
  wire  cp_ctrl_wflags;
  reg [4:0] T_245_cmd;
  reg [31:0] GEN_126;
  reg  T_245_ldst;
  reg [31:0] GEN_127;
  reg  T_245_wen;
  reg [31:0] GEN_128;
  reg  T_245_ren1;
  reg [31:0] GEN_164;
  reg  T_245_ren2;
  reg [31:0] GEN_165;
  reg  T_245_ren3;
  reg [31:0] GEN_166;
  reg  T_245_swap12;
  reg [31:0] GEN_167;
  reg  T_245_swap23;
  reg [31:0] GEN_168;
  reg  T_245_single;
  reg [31:0] GEN_169;
  reg  T_245_fromint;
  reg [31:0] GEN_170;
  reg  T_245_toint;
  reg [31:0] GEN_171;
  reg  T_245_fastpipe;
  reg [31:0] GEN_172;
  reg  T_245_fma;
  reg [31:0] GEN_173;
  reg  T_245_div;
  reg [31:0] GEN_174;
  reg  T_245_sqrt;
  reg [31:0] GEN_175;
  reg  T_245_round;
  reg [31:0] GEN_176;
  reg  T_245_wflags;
  reg [31:0] GEN_177;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [4:0] ex_ctrl_cmd;
  wire  ex_ctrl_ldst;
  wire  ex_ctrl_wen;
  wire  ex_ctrl_ren1;
  wire  ex_ctrl_ren2;
  wire  ex_ctrl_ren3;
  wire  ex_ctrl_swap12;
  wire  ex_ctrl_swap23;
  wire  ex_ctrl_single;
  wire  ex_ctrl_fromint;
  wire  ex_ctrl_toint;
  wire  ex_ctrl_fastpipe;
  wire  ex_ctrl_fma;
  wire  ex_ctrl_div;
  wire  ex_ctrl_sqrt;
  wire  ex_ctrl_round;
  wire  ex_ctrl_wflags;
  reg [4:0] mem_ctrl_cmd;
  reg [31:0] GEN_178;
  reg  mem_ctrl_ldst;
  reg [31:0] GEN_179;
  reg  mem_ctrl_wen;
  reg [31:0] GEN_180;
  reg  mem_ctrl_ren1;
  reg [31:0] GEN_181;
  reg  mem_ctrl_ren2;
  reg [31:0] GEN_182;
  reg  mem_ctrl_ren3;
  reg [31:0] GEN_183;
  reg  mem_ctrl_swap12;
  reg [31:0] GEN_184;
  reg  mem_ctrl_swap23;
  reg [31:0] GEN_185;
  reg  mem_ctrl_single;
  reg [31:0] GEN_186;
  reg  mem_ctrl_fromint;
  reg [31:0] GEN_187;
  reg  mem_ctrl_toint;
  reg [31:0] GEN_188;
  reg  mem_ctrl_fastpipe;
  reg [31:0] GEN_189;
  reg  mem_ctrl_fma;
  reg [31:0] GEN_190;
  reg  mem_ctrl_div;
  reg [31:0] GEN_191;
  reg  mem_ctrl_sqrt;
  reg [31:0] GEN_192;
  reg  mem_ctrl_round;
  reg [31:0] GEN_193;
  reg  mem_ctrl_wflags;
  reg [31:0] GEN_194;
  wire [4:0] GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  reg [4:0] wb_ctrl_cmd;
  reg [31:0] GEN_195;
  reg  wb_ctrl_ldst;
  reg [31:0] GEN_196;
  reg  wb_ctrl_wen;
  reg [31:0] GEN_197;
  reg  wb_ctrl_ren1;
  reg [31:0] GEN_198;
  reg  wb_ctrl_ren2;
  reg [31:0] GEN_199;
  reg  wb_ctrl_ren3;
  reg [31:0] GEN_200;
  reg  wb_ctrl_swap12;
  reg [31:0] GEN_201;
  reg  wb_ctrl_swap23;
  reg [31:0] GEN_202;
  reg  wb_ctrl_single;
  reg [31:0] GEN_203;
  reg  wb_ctrl_fromint;
  reg [31:0] GEN_204;
  reg  wb_ctrl_toint;
  reg [31:0] GEN_205;
  reg  wb_ctrl_fastpipe;
  reg [31:0] GEN_206;
  reg  wb_ctrl_fma;
  reg [31:0] GEN_207;
  reg  wb_ctrl_div;
  reg [31:0] GEN_208;
  reg  wb_ctrl_sqrt;
  reg [31:0] GEN_209;
  reg  wb_ctrl_round;
  reg [31:0] GEN_210;
  reg  wb_ctrl_wflags;
  reg [31:0] GEN_211;
  wire [4:0] GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  reg  load_wb;
  reg [31:0] GEN_212;
  wire  T_314;
  wire  T_316;
  reg  load_wb_single;
  reg [31:0] GEN_213;
  wire  GEN_53;
  reg [63:0] load_wb_data;
  reg [63:0] GEN_214;
  wire [63:0] GEN_54;
  reg [4:0] load_wb_tag;
  reg [31:0] GEN_215;
  wire [4:0] GEN_55;
  wire  T_317;
  wire [7:0] T_318;
  wire [22:0] T_319;
  wire  T_321;
  wire  T_323;
  wire  T_324;
  wire [31:0] GEN_141;
  wire [31:0] T_325;
  wire [15:0] T_326;
  wire [15:0] T_327;
  wire  T_329;
  wire [7:0] T_330;
  wire [7:0] T_331;
  wire  T_333;
  wire [3:0] T_334;
  wire [3:0] T_335;
  wire  T_337;
  wire  T_338;
  wire  T_340;
  wire  T_342;
  wire [1:0] T_344;
  wire [1:0] T_345;
  wire  T_346;
  wire  T_348;
  wire  T_350;
  wire [1:0] T_352;
  wire [1:0] T_353;
  wire [1:0] T_354;
  wire [2:0] T_355;
  wire [3:0] T_356;
  wire [3:0] T_357;
  wire  T_359;
  wire  T_360;
  wire  T_362;
  wire  T_364;
  wire [1:0] T_366;
  wire [1:0] T_367;
  wire  T_368;
  wire  T_370;
  wire  T_372;
  wire [1:0] T_374;
  wire [1:0] T_375;
  wire [1:0] T_376;
  wire [2:0] T_377;
  wire [2:0] T_378;
  wire [3:0] T_379;
  wire [7:0] T_380;
  wire [7:0] T_381;
  wire  T_383;
  wire [3:0] T_384;
  wire [3:0] T_385;
  wire  T_387;
  wire  T_388;
  wire  T_390;
  wire  T_392;
  wire [1:0] T_394;
  wire [1:0] T_395;
  wire  T_396;
  wire  T_398;
  wire  T_400;
  wire [1:0] T_402;
  wire [1:0] T_403;
  wire [1:0] T_404;
  wire [2:0] T_405;
  wire [3:0] T_406;
  wire [3:0] T_407;
  wire  T_409;
  wire  T_410;
  wire  T_412;
  wire  T_414;
  wire [1:0] T_416;
  wire [1:0] T_417;
  wire  T_418;
  wire  T_420;
  wire  T_422;
  wire [1:0] T_424;
  wire [1:0] T_425;
  wire [1:0] T_426;
  wire [2:0] T_427;
  wire [2:0] T_428;
  wire [3:0] T_429;
  wire [3:0] T_430;
  wire [4:0] T_431;
  wire [4:0] T_432;
  wire [53:0] GEN_142;
  wire [53:0] T_433;
  wire [21:0] T_434;
  wire [22:0] T_436;
  wire [8:0] GEN_143;
  wire [8:0] T_442;
  wire [8:0] T_443;
  wire [1:0] T_447;
  wire [7:0] GEN_144;
  wire [7:0] T_448;
  wire [8:0] GEN_145;
  wire [9:0] T_449;
  wire [8:0] T_450;
  wire [1:0] T_451;
  wire  T_453;
  wire  T_455;
  wire  T_456;
  wire [2:0] T_460;
  wire [8:0] GEN_146;
  wire [8:0] T_461;
  wire [8:0] T_462;
  wire [8:0] T_463;
  wire [6:0] GEN_147;
  wire [6:0] T_464;
  wire [8:0] GEN_148;
  wire [8:0] T_465;
  wire [22:0] T_466;
  wire [9:0] T_467;
  wire [32:0] rec_s;
  wire  T_468;
  wire [10:0] T_469;
  wire [51:0] T_470;
  wire  T_472;
  wire  T_474;
  wire  T_475;
  wire [63:0] GEN_149;
  wire [63:0] T_476;
  wire [31:0] T_477;
  wire [31:0] T_478;
  wire  T_480;
  wire [15:0] T_481;
  wire [15:0] T_482;
  wire  T_484;
  wire [7:0] T_485;
  wire [7:0] T_486;
  wire  T_488;
  wire [3:0] T_489;
  wire [3:0] T_490;
  wire  T_492;
  wire  T_493;
  wire  T_495;
  wire  T_497;
  wire [1:0] T_499;
  wire [1:0] T_500;
  wire  T_501;
  wire  T_503;
  wire  T_505;
  wire [1:0] T_507;
  wire [1:0] T_508;
  wire [1:0] T_509;
  wire [2:0] T_510;
  wire [3:0] T_511;
  wire [3:0] T_512;
  wire  T_514;
  wire  T_515;
  wire  T_517;
  wire  T_519;
  wire [1:0] T_521;
  wire [1:0] T_522;
  wire  T_523;
  wire  T_525;
  wire  T_527;
  wire [1:0] T_529;
  wire [1:0] T_530;
  wire [1:0] T_531;
  wire [2:0] T_532;
  wire [2:0] T_533;
  wire [3:0] T_534;
  wire [7:0] T_535;
  wire [7:0] T_536;
  wire  T_538;
  wire [3:0] T_539;
  wire [3:0] T_540;
  wire  T_542;
  wire  T_543;
  wire  T_545;
  wire  T_547;
  wire [1:0] T_549;
  wire [1:0] T_550;
  wire  T_551;
  wire  T_553;
  wire  T_555;
  wire [1:0] T_557;
  wire [1:0] T_558;
  wire [1:0] T_559;
  wire [2:0] T_560;
  wire [3:0] T_561;
  wire [3:0] T_562;
  wire  T_564;
  wire  T_565;
  wire  T_567;
  wire  T_569;
  wire [1:0] T_571;
  wire [1:0] T_572;
  wire  T_573;
  wire  T_575;
  wire  T_577;
  wire [1:0] T_579;
  wire [1:0] T_580;
  wire [1:0] T_581;
  wire [2:0] T_582;
  wire [2:0] T_583;
  wire [3:0] T_584;
  wire [3:0] T_585;
  wire [4:0] T_586;
  wire [15:0] T_587;
  wire [15:0] T_588;
  wire  T_590;
  wire [7:0] T_591;
  wire [7:0] T_592;
  wire  T_594;
  wire [3:0] T_595;
  wire [3:0] T_596;
  wire  T_598;
  wire  T_599;
  wire  T_601;
  wire  T_603;
  wire [1:0] T_605;
  wire [1:0] T_606;
  wire  T_607;
  wire  T_609;
  wire  T_611;
  wire [1:0] T_613;
  wire [1:0] T_614;
  wire [1:0] T_615;
  wire [2:0] T_616;
  wire [3:0] T_617;
  wire [3:0] T_618;
  wire  T_620;
  wire  T_621;
  wire  T_623;
  wire  T_625;
  wire [1:0] T_627;
  wire [1:0] T_628;
  wire  T_629;
  wire  T_631;
  wire  T_633;
  wire [1:0] T_635;
  wire [1:0] T_636;
  wire [1:0] T_637;
  wire [2:0] T_638;
  wire [2:0] T_639;
  wire [3:0] T_640;
  wire [7:0] T_641;
  wire [7:0] T_642;
  wire  T_644;
  wire [3:0] T_645;
  wire [3:0] T_646;
  wire  T_648;
  wire  T_649;
  wire  T_651;
  wire  T_653;
  wire [1:0] T_655;
  wire [1:0] T_656;
  wire  T_657;
  wire  T_659;
  wire  T_661;
  wire [1:0] T_663;
  wire [1:0] T_664;
  wire [1:0] T_665;
  wire [2:0] T_666;
  wire [3:0] T_667;
  wire [3:0] T_668;
  wire  T_670;
  wire  T_671;
  wire  T_673;
  wire  T_675;
  wire [1:0] T_677;
  wire [1:0] T_678;
  wire  T_679;
  wire  T_681;
  wire  T_683;
  wire [1:0] T_685;
  wire [1:0] T_686;
  wire [1:0] T_687;
  wire [2:0] T_688;
  wire [2:0] T_689;
  wire [3:0] T_690;
  wire [3:0] T_691;
  wire [4:0] T_692;
  wire [4:0] T_693;
  wire [5:0] T_694;
  wire [5:0] T_695;
  wire [114:0] GEN_150;
  wire [114:0] T_696;
  wire [50:0] T_697;
  wire [51:0] T_699;
  wire [11:0] GEN_151;
  wire [11:0] T_705;
  wire [11:0] T_706;
  wire [1:0] T_710;
  wire [10:0] GEN_152;
  wire [10:0] T_711;
  wire [11:0] GEN_153;
  wire [12:0] T_712;
  wire [11:0] T_713;
  wire [1:0] T_714;
  wire  T_716;
  wire  T_718;
  wire  T_719;
  wire [2:0] T_723;
  wire [11:0] GEN_154;
  wire [11:0] T_724;
  wire [11:0] T_725;
  wire [11:0] T_726;
  wire [9:0] GEN_155;
  wire [9:0] T_727;
  wire [11:0] GEN_156;
  wire [11:0] T_728;
  wire [51:0] T_729;
  wire [12:0] T_730;
  wire [64:0] T_731;
  wire [64:0] T_733;
  wire [64:0] load_wb_data_recoded;
  reg [64:0] regfile [0:31];
  reg [95:0] GEN_216;
  wire [64:0] regfile_T_802_data;
  wire [4:0] regfile_T_802_addr;
  wire  regfile_T_802_en;
  wire [64:0] regfile_T_803_data;
  wire [4:0] regfile_T_803_addr;
  wire  regfile_T_803_en;
  wire [64:0] regfile_T_804_data;
  wire [4:0] regfile_T_804_addr;
  wire  regfile_T_804_en;
  wire [64:0] regfile_T_736_data;
  wire [4:0] regfile_T_736_addr;
  wire  regfile_T_736_mask;
  wire  regfile_T_736_en;
  wire [64:0] regfile_T_1035_data;
  wire [4:0] regfile_T_1035_addr;
  wire  regfile_T_1035_mask;
  wire  regfile_T_1035_en;
  reg [4:0] ex_ra1;
  reg [31:0] GEN_217;
  reg [4:0] ex_ra2;
  reg [31:0] GEN_218;
  reg [4:0] ex_ra3;
  reg [31:0] GEN_219;
  wire  T_741;
  wire [4:0] T_742;
  wire [4:0] GEN_61;
  wire [4:0] GEN_62;
  wire [4:0] GEN_63;
  wire [4:0] GEN_64;
  wire [4:0] T_744;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire  T_749;
  wire  T_750;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] T_752;
  wire [4:0] GEN_71;
  wire [4:0] GEN_72;
  wire [4:0] GEN_73;
  wire [4:0] GEN_74;
  wire [2:0] T_753;
  wire  T_755;
  wire [2:0] ex_rm;
  wire [4:0] req_cmd;
  wire  req_ldst;
  wire  req_wen;
  wire  req_ren1;
  wire  req_ren2;
  wire  req_ren3;
  wire  req_swap12;
  wire  req_swap23;
  wire  req_single;
  wire  req_fromint;
  wire  req_toint;
  wire  req_fastpipe;
  wire  req_fma;
  wire  req_div;
  wire  req_sqrt;
  wire  req_round;
  wire  req_wflags;
  wire [2:0] req_rm;
  wire [1:0] req_typ;
  wire [64:0] req_in1;
  wire [64:0] req_in2;
  wire [64:0] req_in3;
  wire [1:0] T_805;
  wire [64:0] GEN_75;
  wire [64:0] GEN_76;
  wire [4:0] GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire [2:0] GEN_94;
  wire [1:0] GEN_95;
  wire [64:0] GEN_96;
  wire [64:0] GEN_97;
  wire [64:0] GEN_98;
  wire  sfma_clk;
  wire  sfma_reset;
  wire  sfma_io_in_valid;
  wire [4:0] sfma_io_in_bits_cmd;
  wire  sfma_io_in_bits_ldst;
  wire  sfma_io_in_bits_wen;
  wire  sfma_io_in_bits_ren1;
  wire  sfma_io_in_bits_ren2;
  wire  sfma_io_in_bits_ren3;
  wire  sfma_io_in_bits_swap12;
  wire  sfma_io_in_bits_swap23;
  wire  sfma_io_in_bits_single;
  wire  sfma_io_in_bits_fromint;
  wire  sfma_io_in_bits_toint;
  wire  sfma_io_in_bits_fastpipe;
  wire  sfma_io_in_bits_fma;
  wire  sfma_io_in_bits_div;
  wire  sfma_io_in_bits_sqrt;
  wire  sfma_io_in_bits_round;
  wire  sfma_io_in_bits_wflags;
  wire [2:0] sfma_io_in_bits_rm;
  wire [1:0] sfma_io_in_bits_typ;
  wire [64:0] sfma_io_in_bits_in1;
  wire [64:0] sfma_io_in_bits_in2;
  wire [64:0] sfma_io_in_bits_in3;
  wire  sfma_io_out_valid;
  wire [64:0] sfma_io_out_bits_data;
  wire [4:0] sfma_io_out_bits_exc;
  wire  T_806;
  wire  T_807;
  wire  fpiu_clk;
  wire  fpiu_reset;
  wire  fpiu_io_in_valid;
  wire [4:0] fpiu_io_in_bits_cmd;
  wire  fpiu_io_in_bits_ldst;
  wire  fpiu_io_in_bits_wen;
  wire  fpiu_io_in_bits_ren1;
  wire  fpiu_io_in_bits_ren2;
  wire  fpiu_io_in_bits_ren3;
  wire  fpiu_io_in_bits_swap12;
  wire  fpiu_io_in_bits_swap23;
  wire  fpiu_io_in_bits_single;
  wire  fpiu_io_in_bits_fromint;
  wire  fpiu_io_in_bits_toint;
  wire  fpiu_io_in_bits_fastpipe;
  wire  fpiu_io_in_bits_fma;
  wire  fpiu_io_in_bits_div;
  wire  fpiu_io_in_bits_sqrt;
  wire  fpiu_io_in_bits_round;
  wire  fpiu_io_in_bits_wflags;
  wire [2:0] fpiu_io_in_bits_rm;
  wire [1:0] fpiu_io_in_bits_typ;
  wire [64:0] fpiu_io_in_bits_in1;
  wire [64:0] fpiu_io_in_bits_in2;
  wire [64:0] fpiu_io_in_bits_in3;
  wire [4:0] fpiu_io_as_double_cmd;
  wire  fpiu_io_as_double_ldst;
  wire  fpiu_io_as_double_wen;
  wire  fpiu_io_as_double_ren1;
  wire  fpiu_io_as_double_ren2;
  wire  fpiu_io_as_double_ren3;
  wire  fpiu_io_as_double_swap12;
  wire  fpiu_io_as_double_swap23;
  wire  fpiu_io_as_double_single;
  wire  fpiu_io_as_double_fromint;
  wire  fpiu_io_as_double_toint;
  wire  fpiu_io_as_double_fastpipe;
  wire  fpiu_io_as_double_fma;
  wire  fpiu_io_as_double_div;
  wire  fpiu_io_as_double_sqrt;
  wire  fpiu_io_as_double_round;
  wire  fpiu_io_as_double_wflags;
  wire [2:0] fpiu_io_as_double_rm;
  wire [1:0] fpiu_io_as_double_typ;
  wire [64:0] fpiu_io_as_double_in1;
  wire [64:0] fpiu_io_as_double_in2;
  wire [64:0] fpiu_io_as_double_in3;
  wire  fpiu_io_out_valid;
  wire  fpiu_io_out_bits_lt;
  wire [63:0] fpiu_io_out_bits_store;
  wire [63:0] fpiu_io_out_bits_toint;
  wire [4:0] fpiu_io_out_bits_exc;
  wire  T_808;
  wire  T_809;
  wire [4:0] T_812;
  wire  T_813;
  wire  T_814;
  wire  T_815;
  wire  T_816;
  wire  T_817;
  wire [63:0] GEN_99;
  wire  ifpu_clk;
  wire  ifpu_reset;
  wire  ifpu_io_in_valid;
  wire [4:0] ifpu_io_in_bits_cmd;
  wire  ifpu_io_in_bits_ldst;
  wire  ifpu_io_in_bits_wen;
  wire  ifpu_io_in_bits_ren1;
  wire  ifpu_io_in_bits_ren2;
  wire  ifpu_io_in_bits_ren3;
  wire  ifpu_io_in_bits_swap12;
  wire  ifpu_io_in_bits_swap23;
  wire  ifpu_io_in_bits_single;
  wire  ifpu_io_in_bits_fromint;
  wire  ifpu_io_in_bits_toint;
  wire  ifpu_io_in_bits_fastpipe;
  wire  ifpu_io_in_bits_fma;
  wire  ifpu_io_in_bits_div;
  wire  ifpu_io_in_bits_sqrt;
  wire  ifpu_io_in_bits_round;
  wire  ifpu_io_in_bits_wflags;
  wire [2:0] ifpu_io_in_bits_rm;
  wire [1:0] ifpu_io_in_bits_typ;
  wire [64:0] ifpu_io_in_bits_in1;
  wire [64:0] ifpu_io_in_bits_in2;
  wire [64:0] ifpu_io_in_bits_in3;
  wire  ifpu_io_out_valid;
  wire [64:0] ifpu_io_out_bits_data;
  wire [4:0] ifpu_io_out_bits_exc;
  wire  T_819;
  wire [64:0] T_820;
  wire  fpmu_clk;
  wire  fpmu_reset;
  wire  fpmu_io_in_valid;
  wire [4:0] fpmu_io_in_bits_cmd;
  wire  fpmu_io_in_bits_ldst;
  wire  fpmu_io_in_bits_wen;
  wire  fpmu_io_in_bits_ren1;
  wire  fpmu_io_in_bits_ren2;
  wire  fpmu_io_in_bits_ren3;
  wire  fpmu_io_in_bits_swap12;
  wire  fpmu_io_in_bits_swap23;
  wire  fpmu_io_in_bits_single;
  wire  fpmu_io_in_bits_fromint;
  wire  fpmu_io_in_bits_toint;
  wire  fpmu_io_in_bits_fastpipe;
  wire  fpmu_io_in_bits_fma;
  wire  fpmu_io_in_bits_div;
  wire  fpmu_io_in_bits_sqrt;
  wire  fpmu_io_in_bits_round;
  wire  fpmu_io_in_bits_wflags;
  wire [2:0] fpmu_io_in_bits_rm;
  wire [1:0] fpmu_io_in_bits_typ;
  wire [64:0] fpmu_io_in_bits_in1;
  wire [64:0] fpmu_io_in_bits_in2;
  wire [64:0] fpmu_io_in_bits_in3;
  wire  fpmu_io_out_valid;
  wire [64:0] fpmu_io_out_bits_data;
  wire [4:0] fpmu_io_out_bits_exc;
  wire  fpmu_io_lt;
  wire  T_821;
  reg  divSqrt_wen;
  reg [31:0] GEN_220;
  wire  divSqrt_inReady;
  reg [4:0] divSqrt_waddr;
  reg [31:0] GEN_221;
  wire [64:0] divSqrt_wdata;
  wire [4:0] divSqrt_flags;
  reg  divSqrt_in_flight;
  reg [31:0] GEN_222;
  reg  divSqrt_killed;
  reg [31:0] GEN_223;
  wire  FPUFMAPipe_1_1_clk;
  wire  FPUFMAPipe_1_1_reset;
  wire  FPUFMAPipe_1_1_io_in_valid;
  wire [4:0] FPUFMAPipe_1_1_io_in_bits_cmd;
  wire  FPUFMAPipe_1_1_io_in_bits_ldst;
  wire  FPUFMAPipe_1_1_io_in_bits_wen;
  wire  FPUFMAPipe_1_1_io_in_bits_ren1;
  wire  FPUFMAPipe_1_1_io_in_bits_ren2;
  wire  FPUFMAPipe_1_1_io_in_bits_ren3;
  wire  FPUFMAPipe_1_1_io_in_bits_swap12;
  wire  FPUFMAPipe_1_1_io_in_bits_swap23;
  wire  FPUFMAPipe_1_1_io_in_bits_single;
  wire  FPUFMAPipe_1_1_io_in_bits_fromint;
  wire  FPUFMAPipe_1_1_io_in_bits_toint;
  wire  FPUFMAPipe_1_1_io_in_bits_fastpipe;
  wire  FPUFMAPipe_1_1_io_in_bits_fma;
  wire  FPUFMAPipe_1_1_io_in_bits_div;
  wire  FPUFMAPipe_1_1_io_in_bits_sqrt;
  wire  FPUFMAPipe_1_1_io_in_bits_round;
  wire  FPUFMAPipe_1_1_io_in_bits_wflags;
  wire [2:0] FPUFMAPipe_1_1_io_in_bits_rm;
  wire [1:0] FPUFMAPipe_1_1_io_in_bits_typ;
  wire [64:0] FPUFMAPipe_1_1_io_in_bits_in1;
  wire [64:0] FPUFMAPipe_1_1_io_in_bits_in2;
  wire [64:0] FPUFMAPipe_1_1_io_in_bits_in3;
  wire  FPUFMAPipe_1_1_io_out_valid;
  wire [64:0] FPUFMAPipe_1_1_io_out_bits_data;
  wire [4:0] FPUFMAPipe_1_1_io_out_bits_exc;
  wire  T_831;
  wire  T_832;
  wire  T_839;
  wire  T_844;
  wire  T_845;
  wire [1:0] T_848;
  wire  T_849;
  wire  T_850;
  wire [1:0] GEN_157;
  wire [1:0] memLatencyMask;
  reg [1:0] wen;
  reg [31:0] GEN_224;
  reg [4:0] wbInfo_0_rd;
  reg [31:0] GEN_225;
  reg  wbInfo_0_single;
  reg [31:0] GEN_226;
  reg  wbInfo_0_cp;
  reg [31:0] GEN_227;
  reg [1:0] wbInfo_0_pipeid;
  reg [31:0] GEN_228;
  reg [4:0] wbInfo_1_rd;
  reg [31:0] GEN_229;
  reg  wbInfo_1_single;
  reg [31:0] GEN_230;
  reg  wbInfo_1_cp;
  reg [31:0] GEN_231;
  reg [1:0] wbInfo_1_pipeid;
  reg [31:0] GEN_232;
  wire  T_899;
  wire  T_900;
  wire  mem_wen;
  wire [1:0] T_903;
  wire [1:0] T_906;
  wire  T_907;
  wire [1:0] T_910;
  wire  T_913;
  wire [2:0] T_916;
  wire [1:0] T_917;
  wire [1:0] T_918;
  wire [2:0] GEN_158;
  wire [2:0] T_919;
  wire [2:0] GEN_159;
  wire [2:0] T_920;
  wire  T_922;
  wire  T_923;
  wire [2:0] T_926;
  wire [2:0] T_929;
  wire [2:0] T_933;
  wire [3:0] T_939;
  wire [2:0] T_940;
  wire [2:0] T_941;
  wire [3:0] GEN_160;
  wire [3:0] T_942;
  wire [3:0] GEN_161;
  wire [3:0] T_943;
  wire  T_945;
  wire  T_946;
  reg  write_port_busy;
  reg [31:0] GEN_233;
  wire  GEN_101;
  wire  T_947;
  wire [4:0] GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire [1:0] GEN_105;
  wire  T_948;
  wire [1:0] GEN_162;
  wire [1:0] T_952;
  wire [1:0] GEN_106;
  wire  T_954;
  wire  T_955;
  wire  T_956;
  wire [1:0] T_966;
  wire [1:0] T_972;
  wire [1:0] GEN_163;
  wire [1:0] T_974;
  wire [1:0] T_975;
  wire [4:0] T_976;
  wire  GEN_107;
  wire  GEN_108;
  wire [1:0] GEN_109;
  wire [4:0] GEN_110;
  wire  T_979;
  wire  T_980;
  wire  GEN_111;
  wire  GEN_112;
  wire [1:0] GEN_113;
  wire [4:0] GEN_114;
  wire [1:0] GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire [1:0] GEN_118;
  wire [4:0] GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire [1:0] GEN_122;
  wire [4:0] GEN_123;
  wire [4:0] waddr;
  wire [1:0] T_1002;
  wire  T_1004;
  wire  T_1008;
  wire [64:0] T_1009;
  wire [64:0] T_1014;
  wire [64:0] T_1015;
  wire [64:0] wdata;
  wire [4:0] T_1024;
  wire [4:0] T_1029;
  wire [4:0] wexc;
  wire  T_1031;
  wire  T_1032;
  wire  T_1033;
  wire  T_1034;
  wire  T_1037;
  wire [64:0] GEN_129;
  wire  GEN_130;
  wire  T_1040;
  wire  wb_toint_valid;
  reg [4:0] wb_toint_exc;
  reg [31:0] GEN_234;
  wire [4:0] GEN_131;
  wire  T_1041;
  wire  T_1043;
  wire [4:0] T_1045;
  wire [4:0] T_1047;
  wire [4:0] T_1048;
  wire [4:0] T_1051;
  wire [4:0] T_1052;
  wire  T_1053;
  wire  T_1054;
  wire  T_1056;
  wire  T_1058;
  wire  T_1059;
  wire  units_busy;
  wire  T_1060;
  wire  T_1061;
  wire  T_1062;
  wire  T_1064;
  wire  T_1067;
  wire  T_1068;
  wire  T_1070;
  wire  T_1071;
  wire  T_1072;
  wire  T_1074;
  wire  T_1075;
  reg  T_1079;
  reg [31:0] GEN_235;
  wire  T_1080;
  wire  T_1087;
  wire  T_1088;
  wire  T_1089;
  reg  T_1093;
  reg [31:0] GEN_236;
  reg [1:0] T_1095;
  reg [31:0] GEN_237;
  reg [4:0] T_1097;
  reg [31:0] GEN_238;
  reg [64:0] T_1099;
  reg [95:0] GEN_239;
  wire  DivSqrtRecF64_1_clk;
  wire  DivSqrtRecF64_1_reset;
  wire  DivSqrtRecF64_1_io_inReady_div;
  wire  DivSqrtRecF64_1_io_inReady_sqrt;
  wire  DivSqrtRecF64_1_io_inValid;
  wire  DivSqrtRecF64_1_io_sqrtOp;
  wire [64:0] DivSqrtRecF64_1_io_a;
  wire [64:0] DivSqrtRecF64_1_io_b;
  wire [1:0] DivSqrtRecF64_1_io_roundingMode;
  wire  DivSqrtRecF64_1_io_outValid_div;
  wire  DivSqrtRecF64_1_io_outValid_sqrt;
  wire [64:0] DivSqrtRecF64_1_io_out;
  wire [4:0] DivSqrtRecF64_1_io_exceptionFlags;
  wire  T_1100;
  wire  T_1101;
  wire  T_1105;
  wire  T_1106;
  wire  T_1107;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire [4:0] GEN_135;
  wire [1:0] GEN_136;
  wire  T_1111;
  wire  GEN_137;
  wire [64:0] GEN_138;
  wire  GEN_139;
  wire [4:0] GEN_140;
  wire  RecFNToRecFN_2_1_clk;
  wire  RecFNToRecFN_2_1_reset;
  wire [64:0] RecFNToRecFN_2_1_io_in;
  wire [1:0] RecFNToRecFN_2_1_io_roundingMode;
  wire [32:0] RecFNToRecFN_2_1_io_out;
  wire [4:0] RecFNToRecFN_2_1_io_exceptionFlags;
  wire [64:0] T_1113;
  wire [4:0] T_1115;
  wire [4:0] T_1116;
  wire [4:0] GEN_56;
  reg [31:0] GEN_240;
  FPUDecoder fp_decoder (
    .clk(fp_decoder_clk),
    .reset(fp_decoder_reset),
    .io_inst(fp_decoder_io_inst),
    .io_sigs_cmd(fp_decoder_io_sigs_cmd),
    .io_sigs_ldst(fp_decoder_io_sigs_ldst),
    .io_sigs_wen(fp_decoder_io_sigs_wen),
    .io_sigs_ren1(fp_decoder_io_sigs_ren1),
    .io_sigs_ren2(fp_decoder_io_sigs_ren2),
    .io_sigs_ren3(fp_decoder_io_sigs_ren3),
    .io_sigs_swap12(fp_decoder_io_sigs_swap12),
    .io_sigs_swap23(fp_decoder_io_sigs_swap23),
    .io_sigs_single(fp_decoder_io_sigs_single),
    .io_sigs_fromint(fp_decoder_io_sigs_fromint),
    .io_sigs_toint(fp_decoder_io_sigs_toint),
    .io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),
    .io_sigs_fma(fp_decoder_io_sigs_fma),
    .io_sigs_div(fp_decoder_io_sigs_div),
    .io_sigs_sqrt(fp_decoder_io_sigs_sqrt),
    .io_sigs_round(fp_decoder_io_sigs_round),
    .io_sigs_wflags(fp_decoder_io_sigs_wflags)
  );
  FPUFMAPipe sfma (
    .clk(sfma_clk),
    .reset(sfma_reset),
    .io_in_valid(sfma_io_in_valid),
    .io_in_bits_cmd(sfma_io_in_bits_cmd),
    .io_in_bits_ldst(sfma_io_in_bits_ldst),
    .io_in_bits_wen(sfma_io_in_bits_wen),
    .io_in_bits_ren1(sfma_io_in_bits_ren1),
    .io_in_bits_ren2(sfma_io_in_bits_ren2),
    .io_in_bits_ren3(sfma_io_in_bits_ren3),
    .io_in_bits_swap12(sfma_io_in_bits_swap12),
    .io_in_bits_swap23(sfma_io_in_bits_swap23),
    .io_in_bits_single(sfma_io_in_bits_single),
    .io_in_bits_fromint(sfma_io_in_bits_fromint),
    .io_in_bits_toint(sfma_io_in_bits_toint),
    .io_in_bits_fastpipe(sfma_io_in_bits_fastpipe),
    .io_in_bits_fma(sfma_io_in_bits_fma),
    .io_in_bits_div(sfma_io_in_bits_div),
    .io_in_bits_sqrt(sfma_io_in_bits_sqrt),
    .io_in_bits_round(sfma_io_in_bits_round),
    .io_in_bits_wflags(sfma_io_in_bits_wflags),
    .io_in_bits_rm(sfma_io_in_bits_rm),
    .io_in_bits_typ(sfma_io_in_bits_typ),
    .io_in_bits_in1(sfma_io_in_bits_in1),
    .io_in_bits_in2(sfma_io_in_bits_in2),
    .io_in_bits_in3(sfma_io_in_bits_in3),
    .io_out_valid(sfma_io_out_valid),
    .io_out_bits_data(sfma_io_out_bits_data),
    .io_out_bits_exc(sfma_io_out_bits_exc)
  );
  FPToInt fpiu (
    .clk(fpiu_clk),
    .reset(fpiu_reset),
    .io_in_valid(fpiu_io_in_valid),
    .io_in_bits_cmd(fpiu_io_in_bits_cmd),
    .io_in_bits_ldst(fpiu_io_in_bits_ldst),
    .io_in_bits_wen(fpiu_io_in_bits_wen),
    .io_in_bits_ren1(fpiu_io_in_bits_ren1),
    .io_in_bits_ren2(fpiu_io_in_bits_ren2),
    .io_in_bits_ren3(fpiu_io_in_bits_ren3),
    .io_in_bits_swap12(fpiu_io_in_bits_swap12),
    .io_in_bits_swap23(fpiu_io_in_bits_swap23),
    .io_in_bits_single(fpiu_io_in_bits_single),
    .io_in_bits_fromint(fpiu_io_in_bits_fromint),
    .io_in_bits_toint(fpiu_io_in_bits_toint),
    .io_in_bits_fastpipe(fpiu_io_in_bits_fastpipe),
    .io_in_bits_fma(fpiu_io_in_bits_fma),
    .io_in_bits_div(fpiu_io_in_bits_div),
    .io_in_bits_sqrt(fpiu_io_in_bits_sqrt),
    .io_in_bits_round(fpiu_io_in_bits_round),
    .io_in_bits_wflags(fpiu_io_in_bits_wflags),
    .io_in_bits_rm(fpiu_io_in_bits_rm),
    .io_in_bits_typ(fpiu_io_in_bits_typ),
    .io_in_bits_in1(fpiu_io_in_bits_in1),
    .io_in_bits_in2(fpiu_io_in_bits_in2),
    .io_in_bits_in3(fpiu_io_in_bits_in3),
    .io_as_double_cmd(fpiu_io_as_double_cmd),
    .io_as_double_ldst(fpiu_io_as_double_ldst),
    .io_as_double_wen(fpiu_io_as_double_wen),
    .io_as_double_ren1(fpiu_io_as_double_ren1),
    .io_as_double_ren2(fpiu_io_as_double_ren2),
    .io_as_double_ren3(fpiu_io_as_double_ren3),
    .io_as_double_swap12(fpiu_io_as_double_swap12),
    .io_as_double_swap23(fpiu_io_as_double_swap23),
    .io_as_double_single(fpiu_io_as_double_single),
    .io_as_double_fromint(fpiu_io_as_double_fromint),
    .io_as_double_toint(fpiu_io_as_double_toint),
    .io_as_double_fastpipe(fpiu_io_as_double_fastpipe),
    .io_as_double_fma(fpiu_io_as_double_fma),
    .io_as_double_div(fpiu_io_as_double_div),
    .io_as_double_sqrt(fpiu_io_as_double_sqrt),
    .io_as_double_round(fpiu_io_as_double_round),
    .io_as_double_wflags(fpiu_io_as_double_wflags),
    .io_as_double_rm(fpiu_io_as_double_rm),
    .io_as_double_typ(fpiu_io_as_double_typ),
    .io_as_double_in1(fpiu_io_as_double_in1),
    .io_as_double_in2(fpiu_io_as_double_in2),
    .io_as_double_in3(fpiu_io_as_double_in3),
    .io_out_valid(fpiu_io_out_valid),
    .io_out_bits_lt(fpiu_io_out_bits_lt),
    .io_out_bits_store(fpiu_io_out_bits_store),
    .io_out_bits_toint(fpiu_io_out_bits_toint),
    .io_out_bits_exc(fpiu_io_out_bits_exc)
  );
  IntToFP ifpu (
    .clk(ifpu_clk),
    .reset(ifpu_reset),
    .io_in_valid(ifpu_io_in_valid),
    .io_in_bits_cmd(ifpu_io_in_bits_cmd),
    .io_in_bits_ldst(ifpu_io_in_bits_ldst),
    .io_in_bits_wen(ifpu_io_in_bits_wen),
    .io_in_bits_ren1(ifpu_io_in_bits_ren1),
    .io_in_bits_ren2(ifpu_io_in_bits_ren2),
    .io_in_bits_ren3(ifpu_io_in_bits_ren3),
    .io_in_bits_swap12(ifpu_io_in_bits_swap12),
    .io_in_bits_swap23(ifpu_io_in_bits_swap23),
    .io_in_bits_single(ifpu_io_in_bits_single),
    .io_in_bits_fromint(ifpu_io_in_bits_fromint),
    .io_in_bits_toint(ifpu_io_in_bits_toint),
    .io_in_bits_fastpipe(ifpu_io_in_bits_fastpipe),
    .io_in_bits_fma(ifpu_io_in_bits_fma),
    .io_in_bits_div(ifpu_io_in_bits_div),
    .io_in_bits_sqrt(ifpu_io_in_bits_sqrt),
    .io_in_bits_round(ifpu_io_in_bits_round),
    .io_in_bits_wflags(ifpu_io_in_bits_wflags),
    .io_in_bits_rm(ifpu_io_in_bits_rm),
    .io_in_bits_typ(ifpu_io_in_bits_typ),
    .io_in_bits_in1(ifpu_io_in_bits_in1),
    .io_in_bits_in2(ifpu_io_in_bits_in2),
    .io_in_bits_in3(ifpu_io_in_bits_in3),
    .io_out_valid(ifpu_io_out_valid),
    .io_out_bits_data(ifpu_io_out_bits_data),
    .io_out_bits_exc(ifpu_io_out_bits_exc)
  );
  FPToFP fpmu (
    .clk(fpmu_clk),
    .reset(fpmu_reset),
    .io_in_valid(fpmu_io_in_valid),
    .io_in_bits_cmd(fpmu_io_in_bits_cmd),
    .io_in_bits_ldst(fpmu_io_in_bits_ldst),
    .io_in_bits_wen(fpmu_io_in_bits_wen),
    .io_in_bits_ren1(fpmu_io_in_bits_ren1),
    .io_in_bits_ren2(fpmu_io_in_bits_ren2),
    .io_in_bits_ren3(fpmu_io_in_bits_ren3),
    .io_in_bits_swap12(fpmu_io_in_bits_swap12),
    .io_in_bits_swap23(fpmu_io_in_bits_swap23),
    .io_in_bits_single(fpmu_io_in_bits_single),
    .io_in_bits_fromint(fpmu_io_in_bits_fromint),
    .io_in_bits_toint(fpmu_io_in_bits_toint),
    .io_in_bits_fastpipe(fpmu_io_in_bits_fastpipe),
    .io_in_bits_fma(fpmu_io_in_bits_fma),
    .io_in_bits_div(fpmu_io_in_bits_div),
    .io_in_bits_sqrt(fpmu_io_in_bits_sqrt),
    .io_in_bits_round(fpmu_io_in_bits_round),
    .io_in_bits_wflags(fpmu_io_in_bits_wflags),
    .io_in_bits_rm(fpmu_io_in_bits_rm),
    .io_in_bits_typ(fpmu_io_in_bits_typ),
    .io_in_bits_in1(fpmu_io_in_bits_in1),
    .io_in_bits_in2(fpmu_io_in_bits_in2),
    .io_in_bits_in3(fpmu_io_in_bits_in3),
    .io_out_valid(fpmu_io_out_valid),
    .io_out_bits_data(fpmu_io_out_bits_data),
    .io_out_bits_exc(fpmu_io_out_bits_exc),
    .io_lt(fpmu_io_lt)
  );
  FPUFMAPipe_1 FPUFMAPipe_1_1 (
    .clk(FPUFMAPipe_1_1_clk),
    .reset(FPUFMAPipe_1_1_reset),
    .io_in_valid(FPUFMAPipe_1_1_io_in_valid),
    .io_in_bits_cmd(FPUFMAPipe_1_1_io_in_bits_cmd),
    .io_in_bits_ldst(FPUFMAPipe_1_1_io_in_bits_ldst),
    .io_in_bits_wen(FPUFMAPipe_1_1_io_in_bits_wen),
    .io_in_bits_ren1(FPUFMAPipe_1_1_io_in_bits_ren1),
    .io_in_bits_ren2(FPUFMAPipe_1_1_io_in_bits_ren2),
    .io_in_bits_ren3(FPUFMAPipe_1_1_io_in_bits_ren3),
    .io_in_bits_swap12(FPUFMAPipe_1_1_io_in_bits_swap12),
    .io_in_bits_swap23(FPUFMAPipe_1_1_io_in_bits_swap23),
    .io_in_bits_single(FPUFMAPipe_1_1_io_in_bits_single),
    .io_in_bits_fromint(FPUFMAPipe_1_1_io_in_bits_fromint),
    .io_in_bits_toint(FPUFMAPipe_1_1_io_in_bits_toint),
    .io_in_bits_fastpipe(FPUFMAPipe_1_1_io_in_bits_fastpipe),
    .io_in_bits_fma(FPUFMAPipe_1_1_io_in_bits_fma),
    .io_in_bits_div(FPUFMAPipe_1_1_io_in_bits_div),
    .io_in_bits_sqrt(FPUFMAPipe_1_1_io_in_bits_sqrt),
    .io_in_bits_round(FPUFMAPipe_1_1_io_in_bits_round),
    .io_in_bits_wflags(FPUFMAPipe_1_1_io_in_bits_wflags),
    .io_in_bits_rm(FPUFMAPipe_1_1_io_in_bits_rm),
    .io_in_bits_typ(FPUFMAPipe_1_1_io_in_bits_typ),
    .io_in_bits_in1(FPUFMAPipe_1_1_io_in_bits_in1),
    .io_in_bits_in2(FPUFMAPipe_1_1_io_in_bits_in2),
    .io_in_bits_in3(FPUFMAPipe_1_1_io_in_bits_in3),
    .io_out_valid(FPUFMAPipe_1_1_io_out_valid),
    .io_out_bits_data(FPUFMAPipe_1_1_io_out_bits_data),
    .io_out_bits_exc(FPUFMAPipe_1_1_io_out_bits_exc)
  );
  DivSqrtRecF64 DivSqrtRecF64_1 (
    .clk(DivSqrtRecF64_1_clk),
    .reset(DivSqrtRecF64_1_reset),
    .io_inReady_div(DivSqrtRecF64_1_io_inReady_div),
    .io_inReady_sqrt(DivSqrtRecF64_1_io_inReady_sqrt),
    .io_inValid(DivSqrtRecF64_1_io_inValid),
    .io_sqrtOp(DivSqrtRecF64_1_io_sqrtOp),
    .io_a(DivSqrtRecF64_1_io_a),
    .io_b(DivSqrtRecF64_1_io_b),
    .io_roundingMode(DivSqrtRecF64_1_io_roundingMode),
    .io_outValid_div(DivSqrtRecF64_1_io_outValid_div),
    .io_outValid_sqrt(DivSqrtRecF64_1_io_outValid_sqrt),
    .io_out(DivSqrtRecF64_1_io_out),
    .io_exceptionFlags(DivSqrtRecF64_1_io_exceptionFlags)
  );
  RecFNToRecFN_2 RecFNToRecFN_2_1 (
    .clk(RecFNToRecFN_2_1_clk),
    .reset(RecFNToRecFN_2_1_reset),
    .io_in(RecFNToRecFN_2_1_io_in),
    .io_roundingMode(RecFNToRecFN_2_1_io_roundingMode),
    .io_out(RecFNToRecFN_2_1_io_out),
    .io_exceptionFlags(RecFNToRecFN_2_1_io_exceptionFlags)
  );
  assign io_fcsr_flags_valid = T_1043;
  assign io_fcsr_flags_bits = T_1052;
  assign io_store_data = fpiu_io_out_bits_store;
  assign io_toint_data = fpiu_io_out_bits_toint;
  assign io_fcsr_rdy = T_1070;
  assign io_nack_mem = T_1072;
  assign io_illegal_rm = T_1089;
  assign io_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_dec_wen = fp_decoder_io_sigs_wen;
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_dec_swap12 = fp_decoder_io_sigs_swap12;
  assign io_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_dec_single = fp_decoder_io_sigs_single;
  assign io_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_dec_toint = fp_decoder_io_sigs_toint;
  assign io_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_dec_fma = fp_decoder_io_sigs_fma;
  assign io_dec_div = fp_decoder_io_sigs_div;
  assign io_dec_sqrt = fp_decoder_io_sigs_sqrt;
  assign io_dec_round = fp_decoder_io_sigs_round;
  assign io_dec_wflags = fp_decoder_io_sigs_wflags;
  assign io_sboard_set = T_1080;
  assign io_sboard_clr = T_1087;
  assign io_sboard_clra = waddr;
  assign io_cp_req_ready = T_1040;
  assign io_cp_resp_valid = GEN_130;
  assign io_cp_resp_bits_data = GEN_129;
  assign io_cp_resp_bits_exc = GEN_56;
  assign req_valid = ex_reg_valid | io_cp_req_valid;
  assign GEN_0 = io_valid ? io_inst : ex_reg_inst;
  assign ex_cp_valid = io_cp_req_ready & io_cp_req_valid;
  assign T_194 = io_killx == 1'h0;
  assign T_195 = ex_reg_valid & T_194;
  assign T_196 = T_195 | ex_cp_valid;
  assign GEN_1 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T_199 = io_killm | io_nack_mem;
  assign T_201 = mem_cp_valid == 1'h0;
  assign killm = T_199 & T_201;
  assign T_203 = killm == 1'h0;
  assign T_204 = T_203 | mem_cp_valid;
  assign T_205 = mem_reg_valid & T_204;
  assign fp_decoder_clk = clk;
  assign fp_decoder_reset = reset;
  assign fp_decoder_io_inst = io_inst;
  assign cp_ctrl_cmd = io_cp_req_bits_cmd;
  assign cp_ctrl_ldst = io_cp_req_bits_ldst;
  assign cp_ctrl_wen = io_cp_req_bits_wen;
  assign cp_ctrl_ren1 = io_cp_req_bits_ren1;
  assign cp_ctrl_ren2 = io_cp_req_bits_ren2;
  assign cp_ctrl_ren3 = io_cp_req_bits_ren3;
  assign cp_ctrl_swap12 = io_cp_req_bits_swap12;
  assign cp_ctrl_swap23 = io_cp_req_bits_swap23;
  assign cp_ctrl_single = io_cp_req_bits_single;
  assign cp_ctrl_fromint = io_cp_req_bits_fromint;
  assign cp_ctrl_toint = io_cp_req_bits_toint;
  assign cp_ctrl_fastpipe = io_cp_req_bits_fastpipe;
  assign cp_ctrl_fma = io_cp_req_bits_fma;
  assign cp_ctrl_div = io_cp_req_bits_div;
  assign cp_ctrl_sqrt = io_cp_req_bits_sqrt;
  assign cp_ctrl_round = io_cp_req_bits_round;
  assign cp_ctrl_wflags = io_cp_req_bits_wflags;
  assign GEN_2 = io_valid ? fp_decoder_io_sigs_cmd : T_245_cmd;
  assign GEN_3 = io_valid ? fp_decoder_io_sigs_ldst : T_245_ldst;
  assign GEN_4 = io_valid ? fp_decoder_io_sigs_wen : T_245_wen;
  assign GEN_5 = io_valid ? fp_decoder_io_sigs_ren1 : T_245_ren1;
  assign GEN_6 = io_valid ? fp_decoder_io_sigs_ren2 : T_245_ren2;
  assign GEN_7 = io_valid ? fp_decoder_io_sigs_ren3 : T_245_ren3;
  assign GEN_8 = io_valid ? fp_decoder_io_sigs_swap12 : T_245_swap12;
  assign GEN_9 = io_valid ? fp_decoder_io_sigs_swap23 : T_245_swap23;
  assign GEN_10 = io_valid ? fp_decoder_io_sigs_single : T_245_single;
  assign GEN_11 = io_valid ? fp_decoder_io_sigs_fromint : T_245_fromint;
  assign GEN_12 = io_valid ? fp_decoder_io_sigs_toint : T_245_toint;
  assign GEN_13 = io_valid ? fp_decoder_io_sigs_fastpipe : T_245_fastpipe;
  assign GEN_14 = io_valid ? fp_decoder_io_sigs_fma : T_245_fma;
  assign GEN_15 = io_valid ? fp_decoder_io_sigs_div : T_245_div;
  assign GEN_16 = io_valid ? fp_decoder_io_sigs_sqrt : T_245_sqrt;
  assign GEN_17 = io_valid ? fp_decoder_io_sigs_round : T_245_round;
  assign GEN_18 = io_valid ? fp_decoder_io_sigs_wflags : T_245_wflags;
  assign ex_ctrl_cmd = ex_cp_valid ? cp_ctrl_cmd : T_245_cmd;
  assign ex_ctrl_ldst = ex_cp_valid ? cp_ctrl_ldst : T_245_ldst;
  assign ex_ctrl_wen = ex_cp_valid ? cp_ctrl_wen : T_245_wen;
  assign ex_ctrl_ren1 = ex_cp_valid ? cp_ctrl_ren1 : T_245_ren1;
  assign ex_ctrl_ren2 = ex_cp_valid ? cp_ctrl_ren2 : T_245_ren2;
  assign ex_ctrl_ren3 = ex_cp_valid ? cp_ctrl_ren3 : T_245_ren3;
  assign ex_ctrl_swap12 = ex_cp_valid ? cp_ctrl_swap12 : T_245_swap12;
  assign ex_ctrl_swap23 = ex_cp_valid ? cp_ctrl_swap23 : T_245_swap23;
  assign ex_ctrl_single = ex_cp_valid ? cp_ctrl_single : T_245_single;
  assign ex_ctrl_fromint = ex_cp_valid ? cp_ctrl_fromint : T_245_fromint;
  assign ex_ctrl_toint = ex_cp_valid ? cp_ctrl_toint : T_245_toint;
  assign ex_ctrl_fastpipe = ex_cp_valid ? cp_ctrl_fastpipe : T_245_fastpipe;
  assign ex_ctrl_fma = ex_cp_valid ? cp_ctrl_fma : T_245_fma;
  assign ex_ctrl_div = ex_cp_valid ? cp_ctrl_div : T_245_div;
  assign ex_ctrl_sqrt = ex_cp_valid ? cp_ctrl_sqrt : T_245_sqrt;
  assign ex_ctrl_round = ex_cp_valid ? cp_ctrl_round : T_245_round;
  assign ex_ctrl_wflags = ex_cp_valid ? cp_ctrl_wflags : T_245_wflags;
  assign GEN_19 = req_valid ? ex_ctrl_cmd : mem_ctrl_cmd;
  assign GEN_20 = req_valid ? ex_ctrl_ldst : mem_ctrl_ldst;
  assign GEN_21 = req_valid ? ex_ctrl_wen : mem_ctrl_wen;
  assign GEN_22 = req_valid ? ex_ctrl_ren1 : mem_ctrl_ren1;
  assign GEN_23 = req_valid ? ex_ctrl_ren2 : mem_ctrl_ren2;
  assign GEN_24 = req_valid ? ex_ctrl_ren3 : mem_ctrl_ren3;
  assign GEN_25 = req_valid ? ex_ctrl_swap12 : mem_ctrl_swap12;
  assign GEN_26 = req_valid ? ex_ctrl_swap23 : mem_ctrl_swap23;
  assign GEN_27 = req_valid ? ex_ctrl_single : mem_ctrl_single;
  assign GEN_28 = req_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign GEN_29 = req_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign GEN_30 = req_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign GEN_31 = req_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign GEN_32 = req_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_33 = req_valid ? ex_ctrl_sqrt : mem_ctrl_sqrt;
  assign GEN_34 = req_valid ? ex_ctrl_round : mem_ctrl_round;
  assign GEN_35 = req_valid ? ex_ctrl_wflags : mem_ctrl_wflags;
  assign GEN_36 = mem_reg_valid ? mem_ctrl_cmd : wb_ctrl_cmd;
  assign GEN_37 = mem_reg_valid ? mem_ctrl_ldst : wb_ctrl_ldst;
  assign GEN_38 = mem_reg_valid ? mem_ctrl_wen : wb_ctrl_wen;
  assign GEN_39 = mem_reg_valid ? mem_ctrl_ren1 : wb_ctrl_ren1;
  assign GEN_40 = mem_reg_valid ? mem_ctrl_ren2 : wb_ctrl_ren2;
  assign GEN_41 = mem_reg_valid ? mem_ctrl_ren3 : wb_ctrl_ren3;
  assign GEN_42 = mem_reg_valid ? mem_ctrl_swap12 : wb_ctrl_swap12;
  assign GEN_43 = mem_reg_valid ? mem_ctrl_swap23 : wb_ctrl_swap23;
  assign GEN_44 = mem_reg_valid ? mem_ctrl_single : wb_ctrl_single;
  assign GEN_45 = mem_reg_valid ? mem_ctrl_fromint : wb_ctrl_fromint;
  assign GEN_46 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign GEN_47 = mem_reg_valid ? mem_ctrl_fastpipe : wb_ctrl_fastpipe;
  assign GEN_48 = mem_reg_valid ? mem_ctrl_fma : wb_ctrl_fma;
  assign GEN_49 = mem_reg_valid ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_50 = mem_reg_valid ? mem_ctrl_sqrt : wb_ctrl_sqrt;
  assign GEN_51 = mem_reg_valid ? mem_ctrl_round : wb_ctrl_round;
  assign GEN_52 = mem_reg_valid ? mem_ctrl_wflags : wb_ctrl_wflags;
  assign T_314 = io_dmem_resp_type[0];
  assign T_316 = T_314 == 1'h0;
  assign GEN_53 = io_dmem_resp_val ? T_316 : load_wb_single;
  assign GEN_54 = io_dmem_resp_val ? io_dmem_resp_data : load_wb_data;
  assign GEN_55 = io_dmem_resp_val ? io_dmem_resp_tag : load_wb_tag;
  assign T_317 = load_wb_data[31];
  assign T_318 = load_wb_data[30:23];
  assign T_319 = load_wb_data[22:0];
  assign T_321 = T_318 == 8'h0;
  assign T_323 = T_319 == 23'h0;
  assign T_324 = T_321 & T_323;
  assign GEN_141 = {{9'd0}, T_319};
  assign T_325 = GEN_141 << 9;
  assign T_326 = T_325[31:16];
  assign T_327 = T_325[15:0];
  assign T_329 = T_326 != 16'h0;
  assign T_330 = T_326[15:8];
  assign T_331 = T_326[7:0];
  assign T_333 = T_330 != 8'h0;
  assign T_334 = T_330[7:4];
  assign T_335 = T_330[3:0];
  assign T_337 = T_334 != 4'h0;
  assign T_338 = T_334[3];
  assign T_340 = T_334[2];
  assign T_342 = T_334[1];
  assign T_344 = T_340 ? 2'h2 : {{1'd0}, T_342};
  assign T_345 = T_338 ? 2'h3 : T_344;
  assign T_346 = T_335[3];
  assign T_348 = T_335[2];
  assign T_350 = T_335[1];
  assign T_352 = T_348 ? 2'h2 : {{1'd0}, T_350};
  assign T_353 = T_346 ? 2'h3 : T_352;
  assign T_354 = T_337 ? T_345 : T_353;
  assign T_355 = {T_337,T_354};
  assign T_356 = T_331[7:4];
  assign T_357 = T_331[3:0];
  assign T_359 = T_356 != 4'h0;
  assign T_360 = T_356[3];
  assign T_362 = T_356[2];
  assign T_364 = T_356[1];
  assign T_366 = T_362 ? 2'h2 : {{1'd0}, T_364};
  assign T_367 = T_360 ? 2'h3 : T_366;
  assign T_368 = T_357[3];
  assign T_370 = T_357[2];
  assign T_372 = T_357[1];
  assign T_374 = T_370 ? 2'h2 : {{1'd0}, T_372};
  assign T_375 = T_368 ? 2'h3 : T_374;
  assign T_376 = T_359 ? T_367 : T_375;
  assign T_377 = {T_359,T_376};
  assign T_378 = T_333 ? T_355 : T_377;
  assign T_379 = {T_333,T_378};
  assign T_380 = T_327[15:8];
  assign T_381 = T_327[7:0];
  assign T_383 = T_380 != 8'h0;
  assign T_384 = T_380[7:4];
  assign T_385 = T_380[3:0];
  assign T_387 = T_384 != 4'h0;
  assign T_388 = T_384[3];
  assign T_390 = T_384[2];
  assign T_392 = T_384[1];
  assign T_394 = T_390 ? 2'h2 : {{1'd0}, T_392};
  assign T_395 = T_388 ? 2'h3 : T_394;
  assign T_396 = T_385[3];
  assign T_398 = T_385[2];
  assign T_400 = T_385[1];
  assign T_402 = T_398 ? 2'h2 : {{1'd0}, T_400};
  assign T_403 = T_396 ? 2'h3 : T_402;
  assign T_404 = T_387 ? T_395 : T_403;
  assign T_405 = {T_387,T_404};
  assign T_406 = T_381[7:4];
  assign T_407 = T_381[3:0];
  assign T_409 = T_406 != 4'h0;
  assign T_410 = T_406[3];
  assign T_412 = T_406[2];
  assign T_414 = T_406[1];
  assign T_416 = T_412 ? 2'h2 : {{1'd0}, T_414};
  assign T_417 = T_410 ? 2'h3 : T_416;
  assign T_418 = T_407[3];
  assign T_420 = T_407[2];
  assign T_422 = T_407[1];
  assign T_424 = T_420 ? 2'h2 : {{1'd0}, T_422};
  assign T_425 = T_418 ? 2'h3 : T_424;
  assign T_426 = T_409 ? T_417 : T_425;
  assign T_427 = {T_409,T_426};
  assign T_428 = T_383 ? T_405 : T_427;
  assign T_429 = {T_383,T_428};
  assign T_430 = T_329 ? T_379 : T_429;
  assign T_431 = {T_329,T_430};
  assign T_432 = ~ T_431;
  assign GEN_142 = {{31'd0}, T_319};
  assign T_433 = GEN_142 << T_432;
  assign T_434 = T_433[21:0];
  assign T_436 = {T_434,1'h0};
  assign GEN_143 = {{4'd0}, T_432};
  assign T_442 = GEN_143 ^ 9'h1ff;
  assign T_443 = T_321 ? T_442 : {{1'd0}, T_318};
  assign T_447 = T_321 ? 2'h2 : 2'h1;
  assign GEN_144 = {{6'd0}, T_447};
  assign T_448 = 8'h80 | GEN_144;
  assign GEN_145 = {{1'd0}, T_448};
  assign T_449 = T_443 + GEN_145;
  assign T_450 = T_449[8:0];
  assign T_451 = T_450[8:7];
  assign T_453 = T_451 == 2'h3;
  assign T_455 = T_323 == 1'h0;
  assign T_456 = T_453 & T_455;
  assign T_460 = T_324 ? 3'h7 : 3'h0;
  assign GEN_146 = {{6'd0}, T_460};
  assign T_461 = GEN_146 << 6;
  assign T_462 = ~ T_461;
  assign T_463 = T_450 & T_462;
  assign GEN_147 = {{6'd0}, T_456};
  assign T_464 = GEN_147 << 6;
  assign GEN_148 = {{2'd0}, T_464};
  assign T_465 = T_463 | GEN_148;
  assign T_466 = T_321 ? T_436 : T_319;
  assign T_467 = {T_317,T_465};
  assign rec_s = {T_467,T_466};
  assign T_468 = load_wb_data[63];
  assign T_469 = load_wb_data[62:52];
  assign T_470 = load_wb_data[51:0];
  assign T_472 = T_469 == 11'h0;
  assign T_474 = T_470 == 52'h0;
  assign T_475 = T_472 & T_474;
  assign GEN_149 = {{12'd0}, T_470};
  assign T_476 = GEN_149 << 12;
  assign T_477 = T_476[63:32];
  assign T_478 = T_476[31:0];
  assign T_480 = T_477 != 32'h0;
  assign T_481 = T_477[31:16];
  assign T_482 = T_477[15:0];
  assign T_484 = T_481 != 16'h0;
  assign T_485 = T_481[15:8];
  assign T_486 = T_481[7:0];
  assign T_488 = T_485 != 8'h0;
  assign T_489 = T_485[7:4];
  assign T_490 = T_485[3:0];
  assign T_492 = T_489 != 4'h0;
  assign T_493 = T_489[3];
  assign T_495 = T_489[2];
  assign T_497 = T_489[1];
  assign T_499 = T_495 ? 2'h2 : {{1'd0}, T_497};
  assign T_500 = T_493 ? 2'h3 : T_499;
  assign T_501 = T_490[3];
  assign T_503 = T_490[2];
  assign T_505 = T_490[1];
  assign T_507 = T_503 ? 2'h2 : {{1'd0}, T_505};
  assign T_508 = T_501 ? 2'h3 : T_507;
  assign T_509 = T_492 ? T_500 : T_508;
  assign T_510 = {T_492,T_509};
  assign T_511 = T_486[7:4];
  assign T_512 = T_486[3:0];
  assign T_514 = T_511 != 4'h0;
  assign T_515 = T_511[3];
  assign T_517 = T_511[2];
  assign T_519 = T_511[1];
  assign T_521 = T_517 ? 2'h2 : {{1'd0}, T_519};
  assign T_522 = T_515 ? 2'h3 : T_521;
  assign T_523 = T_512[3];
  assign T_525 = T_512[2];
  assign T_527 = T_512[1];
  assign T_529 = T_525 ? 2'h2 : {{1'd0}, T_527};
  assign T_530 = T_523 ? 2'h3 : T_529;
  assign T_531 = T_514 ? T_522 : T_530;
  assign T_532 = {T_514,T_531};
  assign T_533 = T_488 ? T_510 : T_532;
  assign T_534 = {T_488,T_533};
  assign T_535 = T_482[15:8];
  assign T_536 = T_482[7:0];
  assign T_538 = T_535 != 8'h0;
  assign T_539 = T_535[7:4];
  assign T_540 = T_535[3:0];
  assign T_542 = T_539 != 4'h0;
  assign T_543 = T_539[3];
  assign T_545 = T_539[2];
  assign T_547 = T_539[1];
  assign T_549 = T_545 ? 2'h2 : {{1'd0}, T_547};
  assign T_550 = T_543 ? 2'h3 : T_549;
  assign T_551 = T_540[3];
  assign T_553 = T_540[2];
  assign T_555 = T_540[1];
  assign T_557 = T_553 ? 2'h2 : {{1'd0}, T_555};
  assign T_558 = T_551 ? 2'h3 : T_557;
  assign T_559 = T_542 ? T_550 : T_558;
  assign T_560 = {T_542,T_559};
  assign T_561 = T_536[7:4];
  assign T_562 = T_536[3:0];
  assign T_564 = T_561 != 4'h0;
  assign T_565 = T_561[3];
  assign T_567 = T_561[2];
  assign T_569 = T_561[1];
  assign T_571 = T_567 ? 2'h2 : {{1'd0}, T_569};
  assign T_572 = T_565 ? 2'h3 : T_571;
  assign T_573 = T_562[3];
  assign T_575 = T_562[2];
  assign T_577 = T_562[1];
  assign T_579 = T_575 ? 2'h2 : {{1'd0}, T_577};
  assign T_580 = T_573 ? 2'h3 : T_579;
  assign T_581 = T_564 ? T_572 : T_580;
  assign T_582 = {T_564,T_581};
  assign T_583 = T_538 ? T_560 : T_582;
  assign T_584 = {T_538,T_583};
  assign T_585 = T_484 ? T_534 : T_584;
  assign T_586 = {T_484,T_585};
  assign T_587 = T_478[31:16];
  assign T_588 = T_478[15:0];
  assign T_590 = T_587 != 16'h0;
  assign T_591 = T_587[15:8];
  assign T_592 = T_587[7:0];
  assign T_594 = T_591 != 8'h0;
  assign T_595 = T_591[7:4];
  assign T_596 = T_591[3:0];
  assign T_598 = T_595 != 4'h0;
  assign T_599 = T_595[3];
  assign T_601 = T_595[2];
  assign T_603 = T_595[1];
  assign T_605 = T_601 ? 2'h2 : {{1'd0}, T_603};
  assign T_606 = T_599 ? 2'h3 : T_605;
  assign T_607 = T_596[3];
  assign T_609 = T_596[2];
  assign T_611 = T_596[1];
  assign T_613 = T_609 ? 2'h2 : {{1'd0}, T_611};
  assign T_614 = T_607 ? 2'h3 : T_613;
  assign T_615 = T_598 ? T_606 : T_614;
  assign T_616 = {T_598,T_615};
  assign T_617 = T_592[7:4];
  assign T_618 = T_592[3:0];
  assign T_620 = T_617 != 4'h0;
  assign T_621 = T_617[3];
  assign T_623 = T_617[2];
  assign T_625 = T_617[1];
  assign T_627 = T_623 ? 2'h2 : {{1'd0}, T_625};
  assign T_628 = T_621 ? 2'h3 : T_627;
  assign T_629 = T_618[3];
  assign T_631 = T_618[2];
  assign T_633 = T_618[1];
  assign T_635 = T_631 ? 2'h2 : {{1'd0}, T_633};
  assign T_636 = T_629 ? 2'h3 : T_635;
  assign T_637 = T_620 ? T_628 : T_636;
  assign T_638 = {T_620,T_637};
  assign T_639 = T_594 ? T_616 : T_638;
  assign T_640 = {T_594,T_639};
  assign T_641 = T_588[15:8];
  assign T_642 = T_588[7:0];
  assign T_644 = T_641 != 8'h0;
  assign T_645 = T_641[7:4];
  assign T_646 = T_641[3:0];
  assign T_648 = T_645 != 4'h0;
  assign T_649 = T_645[3];
  assign T_651 = T_645[2];
  assign T_653 = T_645[1];
  assign T_655 = T_651 ? 2'h2 : {{1'd0}, T_653};
  assign T_656 = T_649 ? 2'h3 : T_655;
  assign T_657 = T_646[3];
  assign T_659 = T_646[2];
  assign T_661 = T_646[1];
  assign T_663 = T_659 ? 2'h2 : {{1'd0}, T_661};
  assign T_664 = T_657 ? 2'h3 : T_663;
  assign T_665 = T_648 ? T_656 : T_664;
  assign T_666 = {T_648,T_665};
  assign T_667 = T_642[7:4];
  assign T_668 = T_642[3:0];
  assign T_670 = T_667 != 4'h0;
  assign T_671 = T_667[3];
  assign T_673 = T_667[2];
  assign T_675 = T_667[1];
  assign T_677 = T_673 ? 2'h2 : {{1'd0}, T_675};
  assign T_678 = T_671 ? 2'h3 : T_677;
  assign T_679 = T_668[3];
  assign T_681 = T_668[2];
  assign T_683 = T_668[1];
  assign T_685 = T_681 ? 2'h2 : {{1'd0}, T_683};
  assign T_686 = T_679 ? 2'h3 : T_685;
  assign T_687 = T_670 ? T_678 : T_686;
  assign T_688 = {T_670,T_687};
  assign T_689 = T_644 ? T_666 : T_688;
  assign T_690 = {T_644,T_689};
  assign T_691 = T_590 ? T_640 : T_690;
  assign T_692 = {T_590,T_691};
  assign T_693 = T_480 ? T_586 : T_692;
  assign T_694 = {T_480,T_693};
  assign T_695 = ~ T_694;
  assign GEN_150 = {{63'd0}, T_470};
  assign T_696 = GEN_150 << T_695;
  assign T_697 = T_696[50:0];
  assign T_699 = {T_697,1'h0};
  assign GEN_151 = {{6'd0}, T_695};
  assign T_705 = GEN_151 ^ 12'hfff;
  assign T_706 = T_472 ? T_705 : {{1'd0}, T_469};
  assign T_710 = T_472 ? 2'h2 : 2'h1;
  assign GEN_152 = {{9'd0}, T_710};
  assign T_711 = 11'h400 | GEN_152;
  assign GEN_153 = {{1'd0}, T_711};
  assign T_712 = T_706 + GEN_153;
  assign T_713 = T_712[11:0];
  assign T_714 = T_713[11:10];
  assign T_716 = T_714 == 2'h3;
  assign T_718 = T_474 == 1'h0;
  assign T_719 = T_716 & T_718;
  assign T_723 = T_475 ? 3'h7 : 3'h0;
  assign GEN_154 = {{9'd0}, T_723};
  assign T_724 = GEN_154 << 9;
  assign T_725 = ~ T_724;
  assign T_726 = T_713 & T_725;
  assign GEN_155 = {{9'd0}, T_719};
  assign T_727 = GEN_155 << 9;
  assign GEN_156 = {{2'd0}, T_727};
  assign T_728 = T_726 | GEN_156;
  assign T_729 = T_472 ? T_699 : T_470;
  assign T_730 = {T_468,T_728};
  assign T_731 = {T_730,T_729};
  assign T_733 = {32'hffffffff,rec_s};
  assign load_wb_data_recoded = load_wb_single ? T_733 : T_731;
  assign regfile_T_802_addr = ex_ra1;
  assign regfile_T_802_en = 1'h1;
  assign regfile_T_802_data = regfile[regfile_T_802_addr];
  assign regfile_T_803_addr = ex_ra2;
  assign regfile_T_803_en = 1'h1;
  assign regfile_T_803_data = regfile[regfile_T_803_addr];
  assign regfile_T_804_addr = ex_ra3;
  assign regfile_T_804_en = 1'h1;
  assign regfile_T_804_data = regfile[regfile_T_804_addr];
  assign regfile_T_736_data = load_wb_data_recoded;
  assign regfile_T_736_addr = load_wb_tag;
  assign regfile_T_736_mask = load_wb;
  assign regfile_T_736_en = load_wb;
  assign regfile_T_1035_data = wdata;
  assign regfile_T_1035_addr = waddr;
  assign regfile_T_1035_mask = T_1034;
  assign regfile_T_1035_en = T_1034;
  assign T_741 = fp_decoder_io_sigs_swap12 == 1'h0;
  assign T_742 = io_inst[19:15];
  assign GEN_61 = T_741 ? T_742 : ex_ra1;
  assign GEN_62 = fp_decoder_io_sigs_swap12 ? T_742 : ex_ra2;
  assign GEN_63 = fp_decoder_io_sigs_ren1 ? GEN_61 : ex_ra1;
  assign GEN_64 = fp_decoder_io_sigs_ren1 ? GEN_62 : ex_ra2;
  assign T_744 = io_inst[24:20];
  assign GEN_65 = fp_decoder_io_sigs_swap12 ? T_744 : GEN_63;
  assign GEN_66 = fp_decoder_io_sigs_swap23 ? T_744 : ex_ra3;
  assign T_749 = fp_decoder_io_sigs_swap23 == 1'h0;
  assign T_750 = T_741 & T_749;
  assign GEN_67 = T_750 ? T_744 : GEN_64;
  assign GEN_68 = fp_decoder_io_sigs_ren2 ? GEN_65 : GEN_63;
  assign GEN_69 = fp_decoder_io_sigs_ren2 ? GEN_66 : ex_ra3;
  assign GEN_70 = fp_decoder_io_sigs_ren2 ? GEN_67 : GEN_64;
  assign T_752 = io_inst[31:27];
  assign GEN_71 = fp_decoder_io_sigs_ren3 ? T_752 : GEN_69;
  assign GEN_72 = io_valid ? GEN_68 : ex_ra1;
  assign GEN_73 = io_valid ? GEN_70 : ex_ra2;
  assign GEN_74 = io_valid ? GEN_71 : ex_ra3;
  assign T_753 = ex_reg_inst[14:12];
  assign T_755 = T_753 == 3'h7;
  assign ex_rm = T_755 ? io_fcsr_rm : T_753;
  assign req_cmd = GEN_77;
  assign req_ldst = GEN_78;
  assign req_wen = GEN_79;
  assign req_ren1 = GEN_80;
  assign req_ren2 = GEN_81;
  assign req_ren3 = GEN_82;
  assign req_swap12 = GEN_83;
  assign req_swap23 = GEN_84;
  assign req_single = GEN_85;
  assign req_fromint = GEN_86;
  assign req_toint = GEN_87;
  assign req_fastpipe = GEN_88;
  assign req_fma = GEN_89;
  assign req_div = GEN_90;
  assign req_sqrt = GEN_91;
  assign req_round = GEN_92;
  assign req_wflags = GEN_93;
  assign req_rm = GEN_94;
  assign req_typ = GEN_95;
  assign req_in1 = GEN_96;
  assign req_in2 = GEN_97;
  assign req_in3 = GEN_98;
  assign T_805 = ex_reg_inst[21:20];
  assign GEN_75 = io_cp_req_bits_swap23 ? io_cp_req_bits_in3 : io_cp_req_bits_in2;
  assign GEN_76 = io_cp_req_bits_swap23 ? io_cp_req_bits_in2 : io_cp_req_bits_in3;
  assign GEN_77 = ex_cp_valid ? io_cp_req_bits_cmd : ex_ctrl_cmd;
  assign GEN_78 = ex_cp_valid ? io_cp_req_bits_ldst : ex_ctrl_ldst;
  assign GEN_79 = ex_cp_valid ? io_cp_req_bits_wen : ex_ctrl_wen;
  assign GEN_80 = ex_cp_valid ? io_cp_req_bits_ren1 : ex_ctrl_ren1;
  assign GEN_81 = ex_cp_valid ? io_cp_req_bits_ren2 : ex_ctrl_ren2;
  assign GEN_82 = ex_cp_valid ? io_cp_req_bits_ren3 : ex_ctrl_ren3;
  assign GEN_83 = ex_cp_valid ? io_cp_req_bits_swap12 : ex_ctrl_swap12;
  assign GEN_84 = ex_cp_valid ? io_cp_req_bits_swap23 : ex_ctrl_swap23;
  assign GEN_85 = ex_cp_valid ? io_cp_req_bits_single : ex_ctrl_single;
  assign GEN_86 = ex_cp_valid ? io_cp_req_bits_fromint : ex_ctrl_fromint;
  assign GEN_87 = ex_cp_valid ? io_cp_req_bits_toint : ex_ctrl_toint;
  assign GEN_88 = ex_cp_valid ? io_cp_req_bits_fastpipe : ex_ctrl_fastpipe;
  assign GEN_89 = ex_cp_valid ? io_cp_req_bits_fma : ex_ctrl_fma;
  assign GEN_90 = ex_cp_valid ? io_cp_req_bits_div : ex_ctrl_div;
  assign GEN_91 = ex_cp_valid ? io_cp_req_bits_sqrt : ex_ctrl_sqrt;
  assign GEN_92 = ex_cp_valid ? io_cp_req_bits_round : ex_ctrl_round;
  assign GEN_93 = ex_cp_valid ? io_cp_req_bits_wflags : ex_ctrl_wflags;
  assign GEN_94 = ex_cp_valid ? io_cp_req_bits_rm : ex_rm;
  assign GEN_95 = ex_cp_valid ? io_cp_req_bits_typ : T_805;
  assign GEN_96 = ex_cp_valid ? io_cp_req_bits_in1 : regfile_T_802_data;
  assign GEN_97 = ex_cp_valid ? GEN_75 : regfile_T_803_data;
  assign GEN_98 = ex_cp_valid ? GEN_76 : regfile_T_804_data;
  assign sfma_clk = clk;
  assign sfma_reset = reset;
  assign sfma_io_in_valid = T_807;
  assign sfma_io_in_bits_cmd = req_cmd;
  assign sfma_io_in_bits_ldst = req_ldst;
  assign sfma_io_in_bits_wen = req_wen;
  assign sfma_io_in_bits_ren1 = req_ren1;
  assign sfma_io_in_bits_ren2 = req_ren2;
  assign sfma_io_in_bits_ren3 = req_ren3;
  assign sfma_io_in_bits_swap12 = req_swap12;
  assign sfma_io_in_bits_swap23 = req_swap23;
  assign sfma_io_in_bits_single = req_single;
  assign sfma_io_in_bits_fromint = req_fromint;
  assign sfma_io_in_bits_toint = req_toint;
  assign sfma_io_in_bits_fastpipe = req_fastpipe;
  assign sfma_io_in_bits_fma = req_fma;
  assign sfma_io_in_bits_div = req_div;
  assign sfma_io_in_bits_sqrt = req_sqrt;
  assign sfma_io_in_bits_round = req_round;
  assign sfma_io_in_bits_wflags = req_wflags;
  assign sfma_io_in_bits_rm = req_rm;
  assign sfma_io_in_bits_typ = req_typ;
  assign sfma_io_in_bits_in1 = req_in1;
  assign sfma_io_in_bits_in2 = req_in2;
  assign sfma_io_in_bits_in3 = req_in3;
  assign T_806 = req_valid & ex_ctrl_fma;
  assign T_807 = T_806 & ex_ctrl_single;
  assign fpiu_clk = clk;
  assign fpiu_reset = reset;
  assign fpiu_io_in_valid = T_815;
  assign fpiu_io_in_bits_cmd = req_cmd;
  assign fpiu_io_in_bits_ldst = req_ldst;
  assign fpiu_io_in_bits_wen = req_wen;
  assign fpiu_io_in_bits_ren1 = req_ren1;
  assign fpiu_io_in_bits_ren2 = req_ren2;
  assign fpiu_io_in_bits_ren3 = req_ren3;
  assign fpiu_io_in_bits_swap12 = req_swap12;
  assign fpiu_io_in_bits_swap23 = req_swap23;
  assign fpiu_io_in_bits_single = req_single;
  assign fpiu_io_in_bits_fromint = req_fromint;
  assign fpiu_io_in_bits_toint = req_toint;
  assign fpiu_io_in_bits_fastpipe = req_fastpipe;
  assign fpiu_io_in_bits_fma = req_fma;
  assign fpiu_io_in_bits_div = req_div;
  assign fpiu_io_in_bits_sqrt = req_sqrt;
  assign fpiu_io_in_bits_round = req_round;
  assign fpiu_io_in_bits_wflags = req_wflags;
  assign fpiu_io_in_bits_rm = req_rm;
  assign fpiu_io_in_bits_typ = req_typ;
  assign fpiu_io_in_bits_in1 = req_in1;
  assign fpiu_io_in_bits_in2 = req_in2;
  assign fpiu_io_in_bits_in3 = req_in3;
  assign T_808 = ex_ctrl_toint | ex_ctrl_div;
  assign T_809 = T_808 | ex_ctrl_sqrt;
  assign T_812 = ex_ctrl_cmd & 5'hd;
  assign T_813 = 5'h5 == T_812;
  assign T_814 = T_809 | T_813;
  assign T_815 = req_valid & T_814;
  assign T_816 = fpiu_io_out_valid & mem_cp_valid;
  assign T_817 = T_816 & mem_ctrl_toint;
  assign GEN_99 = T_817 ? fpiu_io_out_bits_toint : 64'h0;
  assign ifpu_clk = clk;
  assign ifpu_reset = reset;
  assign ifpu_io_in_valid = T_819;
  assign ifpu_io_in_bits_cmd = req_cmd;
  assign ifpu_io_in_bits_ldst = req_ldst;
  assign ifpu_io_in_bits_wen = req_wen;
  assign ifpu_io_in_bits_ren1 = req_ren1;
  assign ifpu_io_in_bits_ren2 = req_ren2;
  assign ifpu_io_in_bits_ren3 = req_ren3;
  assign ifpu_io_in_bits_swap12 = req_swap12;
  assign ifpu_io_in_bits_swap23 = req_swap23;
  assign ifpu_io_in_bits_single = req_single;
  assign ifpu_io_in_bits_fromint = req_fromint;
  assign ifpu_io_in_bits_toint = req_toint;
  assign ifpu_io_in_bits_fastpipe = req_fastpipe;
  assign ifpu_io_in_bits_fma = req_fma;
  assign ifpu_io_in_bits_div = req_div;
  assign ifpu_io_in_bits_sqrt = req_sqrt;
  assign ifpu_io_in_bits_round = req_round;
  assign ifpu_io_in_bits_wflags = req_wflags;
  assign ifpu_io_in_bits_rm = req_rm;
  assign ifpu_io_in_bits_typ = req_typ;
  assign ifpu_io_in_bits_in1 = T_820;
  assign ifpu_io_in_bits_in2 = req_in2;
  assign ifpu_io_in_bits_in3 = req_in3;
  assign T_819 = req_valid & ex_ctrl_fromint;
  assign T_820 = ex_cp_valid ? io_cp_req_bits_in1 : {{1'd0}, io_fromint_data};
  assign fpmu_clk = clk;
  assign fpmu_reset = reset;
  assign fpmu_io_in_valid = T_821;
  assign fpmu_io_in_bits_cmd = req_cmd;
  assign fpmu_io_in_bits_ldst = req_ldst;
  assign fpmu_io_in_bits_wen = req_wen;
  assign fpmu_io_in_bits_ren1 = req_ren1;
  assign fpmu_io_in_bits_ren2 = req_ren2;
  assign fpmu_io_in_bits_ren3 = req_ren3;
  assign fpmu_io_in_bits_swap12 = req_swap12;
  assign fpmu_io_in_bits_swap23 = req_swap23;
  assign fpmu_io_in_bits_single = req_single;
  assign fpmu_io_in_bits_fromint = req_fromint;
  assign fpmu_io_in_bits_toint = req_toint;
  assign fpmu_io_in_bits_fastpipe = req_fastpipe;
  assign fpmu_io_in_bits_fma = req_fma;
  assign fpmu_io_in_bits_div = req_div;
  assign fpmu_io_in_bits_sqrt = req_sqrt;
  assign fpmu_io_in_bits_round = req_round;
  assign fpmu_io_in_bits_wflags = req_wflags;
  assign fpmu_io_in_bits_rm = req_rm;
  assign fpmu_io_in_bits_typ = req_typ;
  assign fpmu_io_in_bits_in1 = req_in1;
  assign fpmu_io_in_bits_in2 = req_in2;
  assign fpmu_io_in_bits_in3 = req_in3;
  assign fpmu_io_lt = fpiu_io_out_bits_lt;
  assign T_821 = req_valid & ex_ctrl_fastpipe;
  assign divSqrt_inReady = T_1100;
  assign divSqrt_wdata = T_1113;
  assign divSqrt_flags = T_1116;
  assign FPUFMAPipe_1_1_clk = clk;
  assign FPUFMAPipe_1_1_reset = reset;
  assign FPUFMAPipe_1_1_io_in_valid = T_832;
  assign FPUFMAPipe_1_1_io_in_bits_cmd = req_cmd;
  assign FPUFMAPipe_1_1_io_in_bits_ldst = req_ldst;
  assign FPUFMAPipe_1_1_io_in_bits_wen = req_wen;
  assign FPUFMAPipe_1_1_io_in_bits_ren1 = req_ren1;
  assign FPUFMAPipe_1_1_io_in_bits_ren2 = req_ren2;
  assign FPUFMAPipe_1_1_io_in_bits_ren3 = req_ren3;
  assign FPUFMAPipe_1_1_io_in_bits_swap12 = req_swap12;
  assign FPUFMAPipe_1_1_io_in_bits_swap23 = req_swap23;
  assign FPUFMAPipe_1_1_io_in_bits_single = req_single;
  assign FPUFMAPipe_1_1_io_in_bits_fromint = req_fromint;
  assign FPUFMAPipe_1_1_io_in_bits_toint = req_toint;
  assign FPUFMAPipe_1_1_io_in_bits_fastpipe = req_fastpipe;
  assign FPUFMAPipe_1_1_io_in_bits_fma = req_fma;
  assign FPUFMAPipe_1_1_io_in_bits_div = req_div;
  assign FPUFMAPipe_1_1_io_in_bits_sqrt = req_sqrt;
  assign FPUFMAPipe_1_1_io_in_bits_round = req_round;
  assign FPUFMAPipe_1_1_io_in_bits_wflags = req_wflags;
  assign FPUFMAPipe_1_1_io_in_bits_rm = req_rm;
  assign FPUFMAPipe_1_1_io_in_bits_typ = req_typ;
  assign FPUFMAPipe_1_1_io_in_bits_in1 = req_in1;
  assign FPUFMAPipe_1_1_io_in_bits_in2 = req_in2;
  assign FPUFMAPipe_1_1_io_in_bits_in3 = req_in3;
  assign T_831 = ex_ctrl_single == 1'h0;
  assign T_832 = T_806 & T_831;
  assign T_839 = mem_ctrl_fma & mem_ctrl_single;
  assign T_844 = mem_ctrl_single == 1'h0;
  assign T_845 = mem_ctrl_fma & T_844;
  assign T_848 = T_845 ? 2'h2 : 2'h0;
  assign T_849 = mem_ctrl_fastpipe | mem_ctrl_fromint;
  assign T_850 = T_849 | T_839;
  assign GEN_157 = {{1'd0}, T_850};
  assign memLatencyMask = GEN_157 | T_848;
  assign T_899 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T_900 = T_899 | mem_ctrl_fromint;
  assign mem_wen = mem_reg_valid & T_900;
  assign T_903 = ex_ctrl_fastpipe ? 2'h2 : 2'h0;
  assign T_906 = ex_ctrl_fromint ? 2'h2 : 2'h0;
  assign T_907 = ex_ctrl_fma & ex_ctrl_single;
  assign T_910 = T_907 ? 2'h2 : 2'h0;
  assign T_913 = ex_ctrl_fma & T_831;
  assign T_916 = T_913 ? 3'h4 : 3'h0;
  assign T_917 = T_903 | T_906;
  assign T_918 = T_917 | T_910;
  assign GEN_158 = {{1'd0}, T_918};
  assign T_919 = GEN_158 | T_916;
  assign GEN_159 = {{1'd0}, memLatencyMask};
  assign T_920 = GEN_159 & T_919;
  assign T_922 = T_920 != 3'h0;
  assign T_923 = mem_wen & T_922;
  assign T_926 = ex_ctrl_fastpipe ? 3'h4 : 3'h0;
  assign T_929 = ex_ctrl_fromint ? 3'h4 : 3'h0;
  assign T_933 = T_907 ? 3'h4 : 3'h0;
  assign T_939 = T_913 ? 4'h8 : 4'h0;
  assign T_940 = T_926 | T_929;
  assign T_941 = T_940 | T_933;
  assign GEN_160 = {{1'd0}, T_941};
  assign T_942 = GEN_160 | T_939;
  assign GEN_161 = {{2'd0}, wen};
  assign T_943 = GEN_161 & T_942;
  assign T_945 = T_943 != 4'h0;
  assign T_946 = T_923 | T_945;
  assign GEN_101 = req_valid ? T_946 : write_port_busy;
  assign T_947 = wen[1];
  assign GEN_102 = T_947 ? wbInfo_1_rd : wbInfo_0_rd;
  assign GEN_103 = T_947 ? wbInfo_1_single : wbInfo_0_single;
  assign GEN_104 = T_947 ? wbInfo_1_cp : wbInfo_0_cp;
  assign GEN_105 = T_947 ? wbInfo_1_pipeid : wbInfo_0_pipeid;
  assign T_948 = wen[1:1];
  assign GEN_162 = {{1'd0}, T_948};
  assign T_952 = GEN_162 | memLatencyMask;
  assign GEN_106 = T_203 ? T_952 : {{1'd0}, T_948};
  assign T_954 = write_port_busy == 1'h0;
  assign T_955 = memLatencyMask[0];
  assign T_956 = T_954 & T_955;
  assign T_966 = T_839 ? 2'h2 : 2'h0;
  assign T_972 = T_845 ? 2'h3 : 2'h0;
  assign GEN_163 = {{1'd0}, mem_ctrl_fromint};
  assign T_974 = GEN_163 | T_966;
  assign T_975 = T_974 | T_972;
  assign T_976 = mem_reg_inst[11:7];
  assign GEN_107 = T_956 ? mem_cp_valid : GEN_104;
  assign GEN_108 = T_956 ? mem_ctrl_single : GEN_103;
  assign GEN_109 = T_956 ? T_975 : GEN_105;
  assign GEN_110 = T_956 ? T_976 : GEN_102;
  assign T_979 = memLatencyMask[1];
  assign T_980 = T_954 & T_979;
  assign GEN_111 = T_980 ? mem_cp_valid : wbInfo_1_cp;
  assign GEN_112 = T_980 ? mem_ctrl_single : wbInfo_1_single;
  assign GEN_113 = T_980 ? T_975 : wbInfo_1_pipeid;
  assign GEN_114 = T_980 ? T_976 : wbInfo_1_rd;
  assign GEN_115 = mem_wen ? GEN_106 : {{1'd0}, T_948};
  assign GEN_116 = mem_wen ? GEN_107 : GEN_104;
  assign GEN_117 = mem_wen ? GEN_108 : GEN_103;
  assign GEN_118 = mem_wen ? GEN_109 : GEN_105;
  assign GEN_119 = mem_wen ? GEN_110 : GEN_102;
  assign GEN_120 = mem_wen ? GEN_111 : wbInfo_1_cp;
  assign GEN_121 = mem_wen ? GEN_112 : wbInfo_1_single;
  assign GEN_122 = mem_wen ? GEN_113 : wbInfo_1_pipeid;
  assign GEN_123 = mem_wen ? GEN_114 : wbInfo_1_rd;
  assign waddr = divSqrt_wen ? divSqrt_waddr : wbInfo_0_rd;
  assign T_1002 = wbInfo_0_pipeid & 2'h1;
  assign T_1004 = wbInfo_0_pipeid >= 2'h2;
  assign T_1008 = T_1002 >= 2'h1;
  assign T_1009 = T_1008 ? FPUFMAPipe_1_1_io_out_bits_data : sfma_io_out_bits_data;
  assign T_1014 = T_1008 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T_1015 = T_1004 ? T_1009 : T_1014;
  assign wdata = divSqrt_wen ? divSqrt_wdata : T_1015;
  assign T_1024 = T_1008 ? FPUFMAPipe_1_1_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T_1029 = T_1008 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign wexc = T_1004 ? T_1024 : T_1029;
  assign T_1031 = wbInfo_0_cp == 1'h0;
  assign T_1032 = wen[0];
  assign T_1033 = T_1031 & T_1032;
  assign T_1034 = T_1033 | divSqrt_wen;
  assign T_1037 = wbInfo_0_cp & T_1032;
  assign GEN_129 = T_1037 ? wdata : {{1'd0}, GEN_99};
  assign GEN_130 = T_1037 ? 1'h1 : T_817;
  assign T_1040 = ex_reg_valid == 1'h0;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign GEN_131 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T_1041 = wb_toint_valid | divSqrt_wen;
  assign T_1043 = T_1041 | T_1032;
  assign T_1045 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T_1047 = divSqrt_wen ? divSqrt_flags : 5'h0;
  assign T_1048 = T_1045 | T_1047;
  assign T_1051 = T_1032 ? wexc : 5'h0;
  assign T_1052 = T_1048 | T_1051;
  assign T_1053 = mem_ctrl_div | mem_ctrl_sqrt;
  assign T_1054 = mem_reg_valid & T_1053;
  assign T_1056 = divSqrt_inReady == 1'h0;
  assign T_1058 = wen != 2'h0;
  assign T_1059 = T_1056 | T_1058;
  assign units_busy = T_1054 & T_1059;
  assign T_1060 = ex_reg_valid & ex_ctrl_wflags;
  assign T_1061 = mem_reg_valid & mem_ctrl_wflags;
  assign T_1062 = T_1060 | T_1061;
  assign T_1064 = T_1062 | wb_toint_valid;
  assign T_1067 = T_1064 | T_1058;
  assign T_1068 = T_1067 | divSqrt_in_flight;
  assign T_1070 = T_1068 == 1'h0;
  assign T_1071 = units_busy | write_port_busy;
  assign T_1072 = T_1071 | divSqrt_in_flight;
  assign T_1074 = wb_cp_valid == 1'h0;
  assign T_1075 = wb_reg_valid & T_1074;
  assign T_1080 = T_1075 & T_1079;
  assign T_1087 = T_1074 & divSqrt_wen;
  assign T_1088 = ex_rm[2];
  assign T_1089 = T_1088 & ex_ctrl_round;
  assign DivSqrtRecF64_1_clk = clk;
  assign DivSqrtRecF64_1_reset = reset;
  assign DivSqrtRecF64_1_io_inValid = T_1106;
  assign DivSqrtRecF64_1_io_sqrtOp = mem_ctrl_sqrt;
  assign DivSqrtRecF64_1_io_a = fpiu_io_as_double_in1;
  assign DivSqrtRecF64_1_io_b = fpiu_io_as_double_in2;
  assign DivSqrtRecF64_1_io_roundingMode = fpiu_io_as_double_rm[1:0];
  assign T_1100 = DivSqrtRecF64_1_io_sqrtOp ? DivSqrtRecF64_1_io_inReady_sqrt : DivSqrtRecF64_1_io_inReady_div;
  assign T_1101 = DivSqrtRecF64_1_io_outValid_div | DivSqrtRecF64_1_io_outValid_sqrt;
  assign T_1105 = divSqrt_in_flight == 1'h0;
  assign T_1106 = T_1054 & T_1105;
  assign T_1107 = DivSqrtRecF64_1_io_inValid & divSqrt_inReady;
  assign GEN_132 = T_1107 ? 1'h1 : divSqrt_in_flight;
  assign GEN_133 = T_1107 ? killm : divSqrt_killed;
  assign GEN_134 = T_1107 ? mem_ctrl_single : T_1093;
  assign GEN_135 = T_1107 ? T_976 : divSqrt_waddr;
  assign GEN_136 = T_1107 ? DivSqrtRecF64_1_io_roundingMode : T_1095;
  assign T_1111 = divSqrt_killed == 1'h0;
  assign GEN_137 = T_1101 ? T_1111 : 1'h0;
  assign GEN_138 = T_1101 ? DivSqrtRecF64_1_io_out : T_1099;
  assign GEN_139 = T_1101 ? 1'h0 : GEN_132;
  assign GEN_140 = T_1101 ? DivSqrtRecF64_1_io_exceptionFlags : T_1097;
  assign RecFNToRecFN_2_1_clk = clk;
  assign RecFNToRecFN_2_1_reset = reset;
  assign RecFNToRecFN_2_1_io_in = T_1099;
  assign RecFNToRecFN_2_1_io_roundingMode = T_1095;
  assign T_1113 = T_1093 ? {{32'd0}, RecFNToRecFN_2_1_io_out} : T_1099;
  assign T_1115 = T_1093 ? RecFNToRecFN_2_1_io_exceptionFlags : 5'h0;
  assign T_1116 = T_1097 | T_1115;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_56 = GEN_240[4:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  ex_reg_valid = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  ex_reg_inst = GEN_58[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  mem_reg_valid = GEN_59[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {1{$random}};
  mem_reg_inst = GEN_60[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  mem_cp_valid = GEN_100[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_124 = {1{$random}};
  wb_reg_valid = GEN_124[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  wb_cp_valid = GEN_125[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {1{$random}};
  T_245_cmd = GEN_126[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {1{$random}};
  T_245_ldst = GEN_127[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {1{$random}};
  T_245_wen = GEN_128[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {1{$random}};
  T_245_ren1 = GEN_164[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {1{$random}};
  T_245_ren2 = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_166 = {1{$random}};
  T_245_ren3 = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_167 = {1{$random}};
  T_245_swap12 = GEN_167[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_168 = {1{$random}};
  T_245_swap23 = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_169 = {1{$random}};
  T_245_single = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_170 = {1{$random}};
  T_245_fromint = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_171 = {1{$random}};
  T_245_toint = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_172 = {1{$random}};
  T_245_fastpipe = GEN_172[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_173 = {1{$random}};
  T_245_fma = GEN_173[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_174 = {1{$random}};
  T_245_div = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_175 = {1{$random}};
  T_245_sqrt = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_176 = {1{$random}};
  T_245_round = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_177 = {1{$random}};
  T_245_wflags = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_178 = {1{$random}};
  mem_ctrl_cmd = GEN_178[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_179 = {1{$random}};
  mem_ctrl_ldst = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_180 = {1{$random}};
  mem_ctrl_wen = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_181 = {1{$random}};
  mem_ctrl_ren1 = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_182 = {1{$random}};
  mem_ctrl_ren2 = GEN_182[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_183 = {1{$random}};
  mem_ctrl_ren3 = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_184 = {1{$random}};
  mem_ctrl_swap12 = GEN_184[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_185 = {1{$random}};
  mem_ctrl_swap23 = GEN_185[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_186 = {1{$random}};
  mem_ctrl_single = GEN_186[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_187 = {1{$random}};
  mem_ctrl_fromint = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_188 = {1{$random}};
  mem_ctrl_toint = GEN_188[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_189 = {1{$random}};
  mem_ctrl_fastpipe = GEN_189[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_190 = {1{$random}};
  mem_ctrl_fma = GEN_190[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_191 = {1{$random}};
  mem_ctrl_div = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_192 = {1{$random}};
  mem_ctrl_sqrt = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_193 = {1{$random}};
  mem_ctrl_round = GEN_193[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_194 = {1{$random}};
  mem_ctrl_wflags = GEN_194[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_195 = {1{$random}};
  wb_ctrl_cmd = GEN_195[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_196 = {1{$random}};
  wb_ctrl_ldst = GEN_196[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_197 = {1{$random}};
  wb_ctrl_wen = GEN_197[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_198 = {1{$random}};
  wb_ctrl_ren1 = GEN_198[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_199 = {1{$random}};
  wb_ctrl_ren2 = GEN_199[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_200 = {1{$random}};
  wb_ctrl_ren3 = GEN_200[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_201 = {1{$random}};
  wb_ctrl_swap12 = GEN_201[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_202 = {1{$random}};
  wb_ctrl_swap23 = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_203 = {1{$random}};
  wb_ctrl_single = GEN_203[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_204 = {1{$random}};
  wb_ctrl_fromint = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_205 = {1{$random}};
  wb_ctrl_toint = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_206 = {1{$random}};
  wb_ctrl_fastpipe = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_207 = {1{$random}};
  wb_ctrl_fma = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_208 = {1{$random}};
  wb_ctrl_div = GEN_208[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_209 = {1{$random}};
  wb_ctrl_sqrt = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_210 = {1{$random}};
  wb_ctrl_round = GEN_210[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_211 = {1{$random}};
  wb_ctrl_wflags = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_212 = {1{$random}};
  load_wb = GEN_212[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_213 = {1{$random}};
  load_wb_single = GEN_213[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_214 = {2{$random}};
  load_wb_data = GEN_214[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_215 = {1{$random}};
  load_wb_tag = GEN_215[4:0];
  `endif
  GEN_216 = {3{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = GEN_216[64:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_217 = {1{$random}};
  ex_ra1 = GEN_217[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_218 = {1{$random}};
  ex_ra2 = GEN_218[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_219 = {1{$random}};
  ex_ra3 = GEN_219[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_220 = {1{$random}};
  divSqrt_wen = GEN_220[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_221 = {1{$random}};
  divSqrt_waddr = GEN_221[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_222 = {1{$random}};
  divSqrt_in_flight = GEN_222[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_223 = {1{$random}};
  divSqrt_killed = GEN_223[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_224 = {1{$random}};
  wen = GEN_224[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_225 = {1{$random}};
  wbInfo_0_rd = GEN_225[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_226 = {1{$random}};
  wbInfo_0_single = GEN_226[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_227 = {1{$random}};
  wbInfo_0_cp = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_228 = {1{$random}};
  wbInfo_0_pipeid = GEN_228[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_229 = {1{$random}};
  wbInfo_1_rd = GEN_229[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_230 = {1{$random}};
  wbInfo_1_single = GEN_230[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_231 = {1{$random}};
  wbInfo_1_cp = GEN_231[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_232 = {1{$random}};
  wbInfo_1_pipeid = GEN_232[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_233 = {1{$random}};
  write_port_busy = GEN_233[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_234 = {1{$random}};
  wb_toint_exc = GEN_234[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_235 = {1{$random}};
  T_1079 = GEN_235[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_236 = {1{$random}};
  T_1093 = GEN_236[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_237 = {1{$random}};
  T_1095 = GEN_237[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_238 = {1{$random}};
  T_1097 = GEN_238[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_239 = {3{$random}};
  T_1099 = GEN_239[64:0];
  `endif
  GEN_240 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        ex_reg_inst <= io_inst;
      end
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T_196;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if(reset) begin
      mem_cp_valid <= 1'h0;
    end else begin
      mem_cp_valid <= ex_cp_valid;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T_205;
    end
    if(reset) begin
      wb_cp_valid <= 1'h0;
    end else begin
      wb_cp_valid <= mem_cp_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_cmd <= fp_decoder_io_sigs_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_ldst <= fp_decoder_io_sigs_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_wen <= fp_decoder_io_sigs_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_ren1 <= fp_decoder_io_sigs_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_ren2 <= fp_decoder_io_sigs_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_ren3 <= fp_decoder_io_sigs_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_swap12 <= fp_decoder_io_sigs_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_swap23 <= fp_decoder_io_sigs_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_single <= fp_decoder_io_sigs_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_fromint <= fp_decoder_io_sigs_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_toint <= fp_decoder_io_sigs_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_fastpipe <= fp_decoder_io_sigs_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_fma <= fp_decoder_io_sigs_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_div <= fp_decoder_io_sigs_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_sqrt <= fp_decoder_io_sigs_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_round <= fp_decoder_io_sigs_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        T_245_wflags <= fp_decoder_io_sigs_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_cmd <= cp_ctrl_cmd;
        end else begin
          mem_ctrl_cmd <= T_245_cmd;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_ldst <= cp_ctrl_ldst;
        end else begin
          mem_ctrl_ldst <= T_245_ldst;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_wen <= cp_ctrl_wen;
        end else begin
          mem_ctrl_wen <= T_245_wen;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_ren1 <= cp_ctrl_ren1;
        end else begin
          mem_ctrl_ren1 <= T_245_ren1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_ren2 <= cp_ctrl_ren2;
        end else begin
          mem_ctrl_ren2 <= T_245_ren2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_ren3 <= cp_ctrl_ren3;
        end else begin
          mem_ctrl_ren3 <= T_245_ren3;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_swap12 <= cp_ctrl_swap12;
        end else begin
          mem_ctrl_swap12 <= T_245_swap12;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_swap23 <= cp_ctrl_swap23;
        end else begin
          mem_ctrl_swap23 <= T_245_swap23;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_single <= cp_ctrl_single;
        end else begin
          mem_ctrl_single <= T_245_single;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_fromint <= cp_ctrl_fromint;
        end else begin
          mem_ctrl_fromint <= T_245_fromint;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_toint <= cp_ctrl_toint;
        end else begin
          mem_ctrl_toint <= T_245_toint;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_fastpipe <= cp_ctrl_fastpipe;
        end else begin
          mem_ctrl_fastpipe <= T_245_fastpipe;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_fma <= cp_ctrl_fma;
        end else begin
          mem_ctrl_fma <= T_245_fma;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_div <= cp_ctrl_div;
        end else begin
          mem_ctrl_div <= T_245_div;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_sqrt <= cp_ctrl_sqrt;
        end else begin
          mem_ctrl_sqrt <= T_245_sqrt;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_round <= cp_ctrl_round;
        end else begin
          mem_ctrl_round <= T_245_round;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        if(ex_cp_valid) begin
          mem_ctrl_wflags <= cp_ctrl_wflags;
        end else begin
          mem_ctrl_wflags <= T_245_wflags;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_cmd <= mem_ctrl_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_ldst <= mem_ctrl_ldst;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_wen <= mem_ctrl_wen;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_ren1 <= mem_ctrl_ren1;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_ren2 <= mem_ctrl_ren2;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_ren3 <= mem_ctrl_ren3;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_swap12 <= mem_ctrl_swap12;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_swap23 <= mem_ctrl_swap23;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_single <= mem_ctrl_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_fromint <= mem_ctrl_fromint;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_toint <= mem_ctrl_toint;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_fastpipe <= mem_ctrl_fastpipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_fma <= mem_ctrl_fma;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_div <= mem_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_sqrt <= mem_ctrl_sqrt;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_round <= mem_ctrl_round;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_reg_valid) begin
        wb_ctrl_wflags <= mem_ctrl_wflags;
      end
    end
    if(1'h0) begin
    end else begin
      load_wb <= io_dmem_resp_val;
    end
    if(1'h0) begin
    end else begin
      if(io_dmem_resp_val) begin
        load_wb_single <= T_316;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_dmem_resp_val) begin
        load_wb_data <= io_dmem_resp_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_dmem_resp_val) begin
        load_wb_tag <= io_dmem_resp_tag;
      end
    end
    if(regfile_T_736_en & regfile_T_736_mask) begin
      regfile[regfile_T_736_addr] <= regfile_T_736_data;
    end
    if(regfile_T_1035_en & regfile_T_1035_mask) begin
      regfile[regfile_T_1035_addr] <= regfile_T_1035_data;
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        if(fp_decoder_io_sigs_ren2) begin
          if(fp_decoder_io_sigs_swap12) begin
            ex_ra1 <= T_744;
          end else begin
            if(fp_decoder_io_sigs_ren1) begin
              if(T_741) begin
                ex_ra1 <= T_742;
              end
            end
          end
        end else begin
          if(fp_decoder_io_sigs_ren1) begin
            if(T_741) begin
              ex_ra1 <= T_742;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        if(fp_decoder_io_sigs_ren2) begin
          if(T_750) begin
            ex_ra2 <= T_744;
          end else begin
            if(fp_decoder_io_sigs_ren1) begin
              if(fp_decoder_io_sigs_swap12) begin
                ex_ra2 <= T_742;
              end
            end
          end
        end else begin
          if(fp_decoder_io_sigs_ren1) begin
            if(fp_decoder_io_sigs_swap12) begin
              ex_ra2 <= T_742;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_valid) begin
        if(fp_decoder_io_sigs_ren3) begin
          ex_ra3 <= T_752;
        end else begin
          if(fp_decoder_io_sigs_ren2) begin
            if(fp_decoder_io_sigs_swap23) begin
              ex_ra3 <= T_744;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1101) begin
        divSqrt_wen <= T_1111;
      end else begin
        divSqrt_wen <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1107) begin
        divSqrt_waddr <= T_976;
      end
    end
    if(reset) begin
      divSqrt_in_flight <= 1'h0;
    end else begin
      if(T_1101) begin
        divSqrt_in_flight <= 1'h0;
      end else begin
        if(T_1107) begin
          divSqrt_in_flight <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1107) begin
        divSqrt_killed <= killm;
      end
    end
    if(reset) begin
      wen <= 2'h0;
    end else begin
      if(mem_wen) begin
        if(T_203) begin
          wen <= T_952;
        end else begin
          wen <= {{1'd0}, T_948};
        end
      end else begin
        wen <= {{1'd0}, T_948};
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_956) begin
          wbInfo_0_rd <= T_976;
        end else begin
          if(T_947) begin
            wbInfo_0_rd <= wbInfo_1_rd;
          end
        end
      end else begin
        if(T_947) begin
          wbInfo_0_rd <= wbInfo_1_rd;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_956) begin
          wbInfo_0_single <= mem_ctrl_single;
        end else begin
          if(T_947) begin
            wbInfo_0_single <= wbInfo_1_single;
          end
        end
      end else begin
        if(T_947) begin
          wbInfo_0_single <= wbInfo_1_single;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_956) begin
          wbInfo_0_cp <= mem_cp_valid;
        end else begin
          if(T_947) begin
            wbInfo_0_cp <= wbInfo_1_cp;
          end
        end
      end else begin
        if(T_947) begin
          wbInfo_0_cp <= wbInfo_1_cp;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_956) begin
          wbInfo_0_pipeid <= T_975;
        end else begin
          if(T_947) begin
            wbInfo_0_pipeid <= wbInfo_1_pipeid;
          end
        end
      end else begin
        if(T_947) begin
          wbInfo_0_pipeid <= wbInfo_1_pipeid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_980) begin
          wbInfo_1_rd <= T_976;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_980) begin
          wbInfo_1_single <= mem_ctrl_single;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_980) begin
          wbInfo_1_cp <= mem_cp_valid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_wen) begin
        if(T_980) begin
          wbInfo_1_pipeid <= T_975;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(req_valid) begin
        write_port_busy <= T_946;
      end
    end
    if(1'h0) begin
    end else begin
      if(mem_ctrl_toint) begin
        wb_toint_exc <= fpiu_io_out_bits_exc;
      end
    end
    if(1'h0) begin
    end else begin
      T_1079 <= T_1053;
    end
    if(1'h0) begin
    end else begin
      if(T_1107) begin
        T_1093 <= mem_ctrl_single;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1107) begin
        T_1095 <= DivSqrtRecF64_1_io_roundingMode;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1101) begin
        T_1097 <= DivSqrtRecF64_1_io_exceptionFlags;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1101) begin
        T_1099 <= DivSqrtRecF64_1_io_out;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output [2:0] io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input  [2:0] io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module RRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_prv,
  input   io_in_0_bits_pum,
  input   io_in_0_bits_mxr,
  input  [26:0] io_in_0_bits_addr,
  input   io_in_0_bits_store,
  input   io_in_0_bits_fetch,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_prv,
  input   io_in_1_bits_pum,
  input   io_in_1_bits_mxr,
  input  [26:0] io_in_1_bits_addr,
  input   io_in_1_bits_store,
  input   io_in_1_bits_fetch,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_prv,
  output  io_out_bits_pum,
  output  io_out_bits_mxr,
  output [26:0] io_out_bits_addr,
  output  io_out_bits_store,
  output  io_out_bits_fetch,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_prv;
  wire  GEN_0_bits_pum;
  wire  GEN_0_bits_mxr;
  wire [26:0] GEN_0_bits_addr;
  wire  GEN_0_bits_store;
  wire  GEN_0_bits_fetch;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [26:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_prv;
  wire  GEN_1_bits_pum;
  wire  GEN_1_bits_mxr;
  wire [26:0] GEN_1_bits_addr;
  wire  GEN_1_bits_store;
  wire  GEN_1_bits_fetch;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_prv;
  wire  GEN_2_bits_pum;
  wire  GEN_2_bits_mxr;
  wire [26:0] GEN_2_bits_addr;
  wire  GEN_2_bits_store;
  wire  GEN_2_bits_fetch;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_prv;
  wire  GEN_3_bits_pum;
  wire  GEN_3_bits_mxr;
  wire [26:0] GEN_3_bits_addr;
  wire  GEN_3_bits_store;
  wire  GEN_3_bits_fetch;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_prv;
  wire  GEN_4_bits_pum;
  wire  GEN_4_bits_mxr;
  wire [26:0] GEN_4_bits_addr;
  wire  GEN_4_bits_store;
  wire  GEN_4_bits_fetch;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_prv;
  wire  GEN_5_bits_pum;
  wire  GEN_5_bits_mxr;
  wire [26:0] GEN_5_bits_addr;
  wire  GEN_5_bits_store;
  wire  GEN_5_bits_fetch;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_prv;
  wire  GEN_6_bits_pum;
  wire  GEN_6_bits_mxr;
  wire [26:0] GEN_6_bits_addr;
  wire  GEN_6_bits_store;
  wire  GEN_6_bits_fetch;
  wire  T_220;
  reg  lastGrant;
  reg [31:0] GEN_0;
  wire  GEN_63;
  wire  grantMask_1;
  wire  validMask_1;
  wire  T_224;
  wire  T_228;
  wire  T_230;
  wire  T_234;
  wire  T_235;
  wire  T_236;
  wire  GEN_64;
  wire  GEN_65;
  assign io_in_0_ready = T_235;
  assign io_in_1_ready = T_236;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_prv = GEN_1_bits_prv;
  assign io_out_bits_pum = GEN_2_bits_pum;
  assign io_out_bits_mxr = GEN_3_bits_mxr;
  assign io_out_bits_addr = GEN_4_bits_addr;
  assign io_out_bits_store = GEN_5_bits_store;
  assign io_out_bits_fetch = GEN_6_bits_fetch;
  assign io_chosen = choice;
  assign choice = GEN_65;
  assign GEN_0_ready = GEN_7;
  assign GEN_0_valid = GEN_8;
  assign GEN_0_bits_prv = GEN_9;
  assign GEN_0_bits_pum = GEN_10;
  assign GEN_0_bits_mxr = GEN_11;
  assign GEN_0_bits_addr = GEN_12;
  assign GEN_0_bits_store = GEN_13;
  assign GEN_0_bits_fetch = GEN_14;
  assign GEN_7 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = io_chosen ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign GEN_10 = io_chosen ? io_in_1_bits_pum : io_in_0_bits_pum;
  assign GEN_11 = io_chosen ? io_in_1_bits_mxr : io_in_0_bits_mxr;
  assign GEN_12 = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign GEN_13 = io_chosen ? io_in_1_bits_store : io_in_0_bits_store;
  assign GEN_14 = io_chosen ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign GEN_1_ready = GEN_7;
  assign GEN_1_valid = GEN_8;
  assign GEN_1_bits_prv = GEN_9;
  assign GEN_1_bits_pum = GEN_10;
  assign GEN_1_bits_mxr = GEN_11;
  assign GEN_1_bits_addr = GEN_12;
  assign GEN_1_bits_store = GEN_13;
  assign GEN_1_bits_fetch = GEN_14;
  assign GEN_2_ready = GEN_7;
  assign GEN_2_valid = GEN_8;
  assign GEN_2_bits_prv = GEN_9;
  assign GEN_2_bits_pum = GEN_10;
  assign GEN_2_bits_mxr = GEN_11;
  assign GEN_2_bits_addr = GEN_12;
  assign GEN_2_bits_store = GEN_13;
  assign GEN_2_bits_fetch = GEN_14;
  assign GEN_3_ready = GEN_7;
  assign GEN_3_valid = GEN_8;
  assign GEN_3_bits_prv = GEN_9;
  assign GEN_3_bits_pum = GEN_10;
  assign GEN_3_bits_mxr = GEN_11;
  assign GEN_3_bits_addr = GEN_12;
  assign GEN_3_bits_store = GEN_13;
  assign GEN_3_bits_fetch = GEN_14;
  assign GEN_4_ready = GEN_7;
  assign GEN_4_valid = GEN_8;
  assign GEN_4_bits_prv = GEN_9;
  assign GEN_4_bits_pum = GEN_10;
  assign GEN_4_bits_mxr = GEN_11;
  assign GEN_4_bits_addr = GEN_12;
  assign GEN_4_bits_store = GEN_13;
  assign GEN_4_bits_fetch = GEN_14;
  assign GEN_5_ready = GEN_7;
  assign GEN_5_valid = GEN_8;
  assign GEN_5_bits_prv = GEN_9;
  assign GEN_5_bits_pum = GEN_10;
  assign GEN_5_bits_mxr = GEN_11;
  assign GEN_5_bits_addr = GEN_12;
  assign GEN_5_bits_store = GEN_13;
  assign GEN_5_bits_fetch = GEN_14;
  assign GEN_6_ready = GEN_7;
  assign GEN_6_valid = GEN_8;
  assign GEN_6_bits_prv = GEN_9;
  assign GEN_6_bits_pum = GEN_10;
  assign GEN_6_bits_mxr = GEN_11;
  assign GEN_6_bits_addr = GEN_12;
  assign GEN_6_bits_store = GEN_13;
  assign GEN_6_bits_fetch = GEN_14;
  assign T_220 = io_out_ready & io_out_valid;
  assign GEN_63 = T_220 ? io_chosen : lastGrant;
  assign grantMask_1 = 1'h1 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign T_224 = validMask_1 | io_in_0_valid;
  assign T_228 = validMask_1 == 1'h0;
  assign T_230 = T_224 == 1'h0;
  assign T_234 = grantMask_1 | T_230;
  assign T_235 = T_228 & io_out_ready;
  assign T_236 = T_234 & io_out_ready;
  assign GEN_64 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_65 = validMask_1 ? 1'h1 : GEN_64;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  lastGrant = GEN_0[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_220) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module PTW(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [1:0] io_requestor_0_req_bits_prv,
  input   io_requestor_0_req_bits_pum,
  input   io_requestor_0_req_bits_mxr,
  input  [26:0] io_requestor_0_req_bits_addr,
  input   io_requestor_0_req_bits_store,
  input   io_requestor_0_req_bits_fetch,
  output  io_requestor_0_resp_valid,
  output [15:0] io_requestor_0_resp_bits_pte_reserved_for_hardware,
  output [37:0] io_requestor_0_resp_bits_pte_ppn,
  output [1:0] io_requestor_0_resp_bits_pte_reserved_for_software,
  output  io_requestor_0_resp_bits_pte_d,
  output  io_requestor_0_resp_bits_pte_a,
  output  io_requestor_0_resp_bits_pte_g,
  output  io_requestor_0_resp_bits_pte_u,
  output  io_requestor_0_resp_bits_pte_x,
  output  io_requestor_0_resp_bits_pte_w,
  output  io_requestor_0_resp_bits_pte_r,
  output  io_requestor_0_resp_bits_pte_v,
  output [6:0] io_requestor_0_ptbr_asid,
  output [37:0] io_requestor_0_ptbr_ppn,
  output  io_requestor_0_invalidate,
  output  io_requestor_0_status_debug,
  output [1:0] io_requestor_0_status_prv,
  output  io_requestor_0_status_sd,
  output [30:0] io_requestor_0_status_zero3,
  output  io_requestor_0_status_sd_rv32,
  output [1:0] io_requestor_0_status_zero2,
  output [4:0] io_requestor_0_status_vm,
  output [3:0] io_requestor_0_status_zero1,
  output  io_requestor_0_status_mxr,
  output  io_requestor_0_status_pum,
  output  io_requestor_0_status_mprv,
  output [1:0] io_requestor_0_status_xs,
  output [1:0] io_requestor_0_status_fs,
  output [1:0] io_requestor_0_status_mpp,
  output [1:0] io_requestor_0_status_hpp,
  output  io_requestor_0_status_spp,
  output  io_requestor_0_status_mpie,
  output  io_requestor_0_status_hpie,
  output  io_requestor_0_status_spie,
  output  io_requestor_0_status_upie,
  output  io_requestor_0_status_mie,
  output  io_requestor_0_status_hie,
  output  io_requestor_0_status_sie,
  output  io_requestor_0_status_uie,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [1:0] io_requestor_1_req_bits_prv,
  input   io_requestor_1_req_bits_pum,
  input   io_requestor_1_req_bits_mxr,
  input  [26:0] io_requestor_1_req_bits_addr,
  input   io_requestor_1_req_bits_store,
  input   io_requestor_1_req_bits_fetch,
  output  io_requestor_1_resp_valid,
  output [15:0] io_requestor_1_resp_bits_pte_reserved_for_hardware,
  output [37:0] io_requestor_1_resp_bits_pte_ppn,
  output [1:0] io_requestor_1_resp_bits_pte_reserved_for_software,
  output  io_requestor_1_resp_bits_pte_d,
  output  io_requestor_1_resp_bits_pte_a,
  output  io_requestor_1_resp_bits_pte_g,
  output  io_requestor_1_resp_bits_pte_u,
  output  io_requestor_1_resp_bits_pte_x,
  output  io_requestor_1_resp_bits_pte_w,
  output  io_requestor_1_resp_bits_pte_r,
  output  io_requestor_1_resp_bits_pte_v,
  output [6:0] io_requestor_1_ptbr_asid,
  output [37:0] io_requestor_1_ptbr_ppn,
  output  io_requestor_1_invalidate,
  output  io_requestor_1_status_debug,
  output [1:0] io_requestor_1_status_prv,
  output  io_requestor_1_status_sd,
  output [30:0] io_requestor_1_status_zero3,
  output  io_requestor_1_status_sd_rv32,
  output [1:0] io_requestor_1_status_zero2,
  output [4:0] io_requestor_1_status_vm,
  output [3:0] io_requestor_1_status_zero1,
  output  io_requestor_1_status_mxr,
  output  io_requestor_1_status_pum,
  output  io_requestor_1_status_mprv,
  output [1:0] io_requestor_1_status_xs,
  output [1:0] io_requestor_1_status_fs,
  output [1:0] io_requestor_1_status_mpp,
  output [1:0] io_requestor_1_status_hpp,
  output  io_requestor_1_status_spp,
  output  io_requestor_1_status_mpie,
  output  io_requestor_1_status_hpie,
  output  io_requestor_1_status_spie,
  output  io_requestor_1_status_upie,
  output  io_requestor_1_status_mie,
  output  io_requestor_1_status_hie,
  output  io_requestor_1_status_sie,
  output  io_requestor_1_status_uie,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [6:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered,
  input  [6:0] io_dpath_ptbr_asid,
  input  [37:0] io_dpath_ptbr_ppn,
  input   io_dpath_invalidate,
  input   io_dpath_status_debug,
  input  [1:0] io_dpath_status_prv,
  input   io_dpath_status_sd,
  input  [30:0] io_dpath_status_zero3,
  input   io_dpath_status_sd_rv32,
  input  [1:0] io_dpath_status_zero2,
  input  [4:0] io_dpath_status_vm,
  input  [3:0] io_dpath_status_zero1,
  input   io_dpath_status_mxr,
  input   io_dpath_status_pum,
  input   io_dpath_status_mprv,
  input  [1:0] io_dpath_status_xs,
  input  [1:0] io_dpath_status_fs,
  input  [1:0] io_dpath_status_mpp,
  input  [1:0] io_dpath_status_hpp,
  input   io_dpath_status_spp,
  input   io_dpath_status_mpie,
  input   io_dpath_status_hpie,
  input   io_dpath_status_spie,
  input   io_dpath_status_upie,
  input   io_dpath_status_mie,
  input   io_dpath_status_hie,
  input   io_dpath_status_sie,
  input   io_dpath_status_uie
);
  reg [2:0] state;
  reg [31:0] GEN_51;
  reg [1:0] count;
  reg [31:0] GEN_125;
  reg  s1_kill;
  reg [31:0] GEN_127;
  reg [1:0] r_req_prv;
  reg [31:0] GEN_128;
  reg  r_req_pum;
  reg [31:0] GEN_129;
  reg  r_req_mxr;
  reg [31:0] GEN_130;
  reg [26:0] r_req_addr;
  reg [31:0] GEN_131;
  reg  r_req_store;
  reg [31:0] GEN_132;
  reg  r_req_fetch;
  reg [31:0] GEN_133;
  reg  r_req_dest;
  reg [31:0] GEN_134;
  reg [15:0] r_pte_reserved_for_hardware;
  reg [31:0] GEN_135;
  reg [37:0] r_pte_ppn;
  reg [63:0] GEN_136;
  reg [1:0] r_pte_reserved_for_software;
  reg [31:0] GEN_137;
  reg  r_pte_d;
  reg [31:0] GEN_138;
  reg  r_pte_a;
  reg [31:0] GEN_139;
  reg  r_pte_g;
  reg [31:0] GEN_140;
  reg  r_pte_u;
  reg [31:0] GEN_141;
  reg  r_pte_x;
  reg [31:0] GEN_142;
  reg  r_pte_w;
  reg [31:0] GEN_143;
  reg  r_pte_r;
  reg [31:0] GEN_144;
  reg  r_pte_v;
  reg [31:0] GEN_145;
  wire [8:0] T_2185;
  wire [17:0] T_2186;
  wire [8:0] vpn_idxs_1;
  wire [8:0] vpn_idxs_2;
  wire [1:0] T_2189;
  wire  T_2191;
  wire  T_2195;
  wire [8:0] T_2196;
  wire [8:0] vpn_idx;
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_prv;
  wire  arb_io_in_0_bits_pum;
  wire  arb_io_in_0_bits_mxr;
  wire [26:0] arb_io_in_0_bits_addr;
  wire  arb_io_in_0_bits_store;
  wire  arb_io_in_0_bits_fetch;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_prv;
  wire  arb_io_in_1_bits_pum;
  wire  arb_io_in_1_bits_mxr;
  wire [26:0] arb_io_in_1_bits_addr;
  wire  arb_io_in_1_bits_store;
  wire  arb_io_in_1_bits_fetch;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_prv;
  wire  arb_io_out_bits_pum;
  wire  arb_io_out_bits_mxr;
  wire [26:0] arb_io_out_bits_addr;
  wire  arb_io_out_bits_store;
  wire  arb_io_out_bits_fetch;
  wire  arb_io_chosen;
  wire  T_2204;
  wire [15:0] T_2229_reserved_for_hardware;
  wire [37:0] T_2229_ppn;
  wire [1:0] T_2229_reserved_for_software;
  wire  T_2229_d;
  wire  T_2229_a;
  wire  T_2229_g;
  wire  T_2229_u;
  wire  T_2229_x;
  wire  T_2229_w;
  wire  T_2229_r;
  wire  T_2229_v;
  wire  T_2241;
  wire  T_2242;
  wire  T_2243;
  wire  T_2244;
  wire  T_2245;
  wire  T_2246;
  wire  T_2247;
  wire  T_2248;
  wire [1:0] T_2249;
  wire [37:0] T_2250;
  wire [15:0] T_2251;
  wire [15:0] T_2276_reserved_for_hardware;
  wire [37:0] T_2276_ppn;
  wire [1:0] T_2276_reserved_for_software;
  wire  T_2276_d;
  wire  T_2276_a;
  wire  T_2276_g;
  wire  T_2276_u;
  wire  T_2276_x;
  wire  T_2276_w;
  wire  T_2276_r;
  wire  T_2276_v;
  wire [15:0] pte_reserved_for_hardware;
  wire [37:0] pte_ppn;
  wire [1:0] pte_reserved_for_software;
  wire  pte_d;
  wire  pte_a;
  wire  pte_g;
  wire  pte_u;
  wire  pte_x;
  wire  pte_w;
  wire  pte_r;
  wire  pte_v;
  wire [19:0] T_2310;
  wire [17:0] T_2311;
  wire  T_2313;
  wire  GEN_2;
  wire [46:0] T_2315;
  wire [49:0] GEN_115;
  wire [49:0] pte_addr;
  wire  T_2316;
  wire [1:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [26:0] GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire [37:0] GEN_10;
  reg [7:0] T_2318;
  reg [31:0] GEN_146;
  reg [7:0] T_2320;
  reg [31:0] GEN_147;
  reg [31:0] T_2327_0;
  reg [31:0] GEN_148;
  reg [31:0] T_2327_1;
  reg [31:0] GEN_149;
  reg [31:0] T_2327_2;
  reg [31:0] GEN_150;
  reg [31:0] T_2327_3;
  reg [31:0] GEN_151;
  reg [31:0] T_2327_4;
  reg [31:0] GEN_152;
  reg [31:0] T_2327_5;
  reg [31:0] GEN_153;
  reg [31:0] T_2327_6;
  reg [31:0] GEN_154;
  reg [31:0] T_2327_7;
  reg [31:0] GEN_155;
  reg [19:0] T_2335_0;
  reg [31:0] GEN_156;
  reg [19:0] T_2335_1;
  reg [31:0] GEN_157;
  reg [19:0] T_2335_2;
  reg [31:0] GEN_158;
  reg [19:0] T_2335_3;
  reg [31:0] GEN_159;
  reg [19:0] T_2335_4;
  reg [31:0] GEN_160;
  reg [19:0] T_2335_5;
  reg [31:0] GEN_161;
  reg [19:0] T_2335_6;
  reg [31:0] GEN_162;
  reg [19:0] T_2335_7;
  reg [31:0] GEN_163;
  wire [49:0] GEN_116;
  wire  T_2337;
  wire [49:0] GEN_117;
  wire  T_2338;
  wire [49:0] GEN_118;
  wire  T_2339;
  wire [49:0] GEN_119;
  wire  T_2340;
  wire [49:0] GEN_120;
  wire  T_2341;
  wire [49:0] GEN_121;
  wire  T_2342;
  wire [49:0] GEN_122;
  wire  T_2343;
  wire [49:0] GEN_123;
  wire  T_2344;
  wire [1:0] T_2345;
  wire [1:0] T_2346;
  wire [3:0] T_2347;
  wire [1:0] T_2348;
  wire [1:0] T_2349;
  wire [3:0] T_2350;
  wire [7:0] T_2351;
  wire [7:0] T_2352;
  wire  T_2354;
  wire  T_2356;
  wire  T_2357;
  wire  T_2359;
  wire  T_2360;
  wire  T_2362;
  wire  T_2363;
  wire  T_2364;
  wire  T_2366;
  wire  T_2367;
  wire [7:0] T_2368;
  wire  T_2370;
  wire [7:0] T_2372;
  wire  T_2373;
  wire [1:0] T_2374;
  wire [7:0] T_2375;
  wire  T_2376;
  wire [2:0] T_2377;
  wire [7:0] T_2378;
  wire  T_2379;
  wire [3:0] T_2380;
  wire [2:0] T_2381;
  wire  T_2383;
  wire  T_2384;
  wire  T_2385;
  wire  T_2386;
  wire  T_2387;
  wire  T_2388;
  wire  T_2389;
  wire [2:0] T_2399;
  wire [2:0] T_2400;
  wire [2:0] T_2401;
  wire [2:0] T_2402;
  wire [2:0] T_2403;
  wire [2:0] T_2404;
  wire [2:0] T_2405;
  wire [2:0] T_2406;
  wire [7:0] T_2408;
  wire [7:0] T_2409;
  wire [31:0] GEN_0;
  wire [31:0] GEN_11;
  wire [31:0] GEN_12;
  wire [31:0] GEN_13;
  wire [31:0] GEN_14;
  wire [31:0] GEN_15;
  wire [31:0] GEN_16;
  wire [31:0] GEN_17;
  wire [31:0] GEN_18;
  wire [19:0] GEN_1;
  wire [19:0] GEN_19;
  wire [19:0] GEN_20;
  wire [19:0] GEN_21;
  wire [19:0] GEN_22;
  wire [19:0] GEN_23;
  wire [19:0] GEN_24;
  wire [19:0] GEN_25;
  wire [19:0] GEN_26;
  wire [7:0] GEN_27;
  wire [31:0] GEN_29;
  wire [31:0] GEN_30;
  wire [31:0] GEN_31;
  wire [31:0] GEN_32;
  wire [31:0] GEN_33;
  wire [31:0] GEN_34;
  wire [31:0] GEN_35;
  wire [31:0] GEN_36;
  wire [19:0] GEN_38;
  wire [19:0] GEN_39;
  wire [19:0] GEN_40;
  wire [19:0] GEN_41;
  wire [19:0] GEN_42;
  wire [19:0] GEN_43;
  wire [19:0] GEN_44;
  wire [19:0] GEN_45;
  wire  T_2410;
  wire  T_2411;
  wire [3:0] T_2412;
  wire [3:0] T_2413;
  wire  T_2415;
  wire [3:0] T_2416;
  wire [1:0] T_2417;
  wire [1:0] T_2418;
  wire  T_2420;
  wire [1:0] T_2421;
  wire  T_2422;
  wire [1:0] T_2423;
  wire [2:0] T_2424;
  wire  T_2426;
  wire  T_2428;
  wire [1:0] T_2430;
  wire [7:0] GEN_124;
  wire [7:0] T_2431;
  wire [7:0] T_2432;
  wire [7:0] T_2433;
  wire [7:0] T_2434;
  wire [7:0] T_2435;
  wire [1:0] T_2436;
  wire  T_2437;
  wire  T_2439;
  wire [3:0] T_2441;
  wire [7:0] GEN_126;
  wire [7:0] T_2442;
  wire [7:0] T_2443;
  wire [7:0] T_2444;
  wire [7:0] T_2445;
  wire [7:0] T_2446;
  wire [2:0] T_2447;
  wire  T_2448;
  wire  T_2450;
  wire [7:0] T_2452;
  wire [7:0] T_2453;
  wire [7:0] T_2454;
  wire [7:0] T_2455;
  wire [7:0] T_2456;
  wire [7:0] T_2457;
  wire [7:0] GEN_46;
  wire [7:0] GEN_47;
  wire  T_2461;
  wire  pte_cache_hit;
  wire  T_2462;
  wire  T_2463;
  wire  T_2464;
  wire  T_2465;
  wire  T_2466;
  wire  T_2467;
  wire  T_2468;
  wire  T_2469;
  wire [19:0] T_2471;
  wire [19:0] T_2473;
  wire [19:0] T_2475;
  wire [19:0] T_2477;
  wire [19:0] T_2479;
  wire [19:0] T_2481;
  wire [19:0] T_2483;
  wire [19:0] T_2485;
  wire [19:0] T_2487;
  wire [19:0] T_2488;
  wire [19:0] T_2489;
  wire [19:0] T_2490;
  wire [19:0] T_2491;
  wire [19:0] T_2492;
  wire [19:0] T_2493;
  wire [19:0] pte_cache_data;
  wire [15:0] T_2519_reserved_for_hardware;
  wire [37:0] T_2519_ppn;
  wire [1:0] T_2519_reserved_for_software;
  wire  T_2519_d;
  wire  T_2519_a;
  wire  T_2519_g;
  wire  T_2519_u;
  wire  T_2519_x;
  wire  T_2519_w;
  wire  T_2519_r;
  wire  T_2519_v;
  wire [63:0] T_2532;
  wire  T_2533;
  wire  T_2534;
  wire  T_2535;
  wire  T_2536;
  wire  T_2537;
  wire  T_2538;
  wire  T_2539;
  wire  T_2540;
  wire [1:0] T_2541;
  wire [37:0] T_2542;
  wire [15:0] T_2543;
  wire [15:0] pte_wdata_reserved_for_hardware;
  wire [37:0] pte_wdata_ppn;
  wire [1:0] pte_wdata_reserved_for_software;
  wire  pte_wdata_d;
  wire  pte_wdata_a;
  wire  pte_wdata_g;
  wire  pte_wdata_u;
  wire  pte_wdata_x;
  wire  pte_wdata_w;
  wire  pte_wdata_r;
  wire  pte_wdata_v;
  wire  T_2557;
  wire  T_2558;
  wire [4:0] T_2561;
  wire [1:0] T_2563;
  wire [1:0] T_2564;
  wire [2:0] T_2565;
  wire [4:0] T_2566;
  wire [1:0] T_2567;
  wire [2:0] T_2568;
  wire [53:0] T_2569;
  wire [55:0] T_2570;
  wire [58:0] T_2571;
  wire [63:0] T_2572;
  wire [19:0] T_2574;
  wire [17:0] T_2575;
  wire [37:0] resp_ppns_0;
  wire [28:0] T_2576;
  wire [37:0] resp_ppns_1;
  wire [37:0] resp_ppns_2;
  wire  T_2578;
  wire  T_2580;
  wire  T_2581;
  wire [37:0] T_2590;
  wire [37:0] T_2591;
  wire  T_2595;
  wire  T_2606;
  wire [2:0] GEN_48;
  wire [2:0] GEN_49;
  wire [1:0] GEN_50;
  wire  T_2608;
  wire [2:0] T_2611;
  wire [1:0] T_2612;
  wire [2:0] GEN_52;
  wire [1:0] GEN_53;
  wire [37:0] GEN_54;
  wire  T_2614;
  wire  T_2615;
  wire [2:0] GEN_55;
  wire  GEN_56;
  wire [2:0] GEN_57;
  wire [1:0] GEN_58;
  wire [37:0] GEN_59;
  wire  T_2616;
  wire  GEN_60;
  wire [2:0] GEN_61;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire  T_2618;
  wire [2:0] GEN_64;
  wire  T_2619;
  wire  T_2620;
  wire  T_2621;
  wire  T_2622;
  wire  T_2624;
  wire  T_2625;
  wire  T_2626;
  wire  T_2629;
  wire  T_2630;
  wire  T_2631;
  wire  T_2632;
  wire  T_2633;
  wire  T_2635;
  wire  T_2637;
  wire  T_2638;
  wire  T_2639;
  wire  T_2640;
  wire [2:0] GEN_65;
  wire  T_2642;
  wire [15:0] GEN_66;
  wire [37:0] GEN_67;
  wire [1:0] GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  T_2654;
  wire [2:0] GEN_77;
  wire [1:0] GEN_78;
  wire [2:0] GEN_79;
  wire [15:0] GEN_80;
  wire [37:0] GEN_81;
  wire [1:0] GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire [1:0] GEN_91;
  wire [2:0] GEN_92;
  wire [15:0] GEN_93;
  wire [37:0] GEN_94;
  wire [1:0] GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire [1:0] GEN_104;
  wire  T_2658;
  wire [2:0] GEN_105;
  wire [2:0] GEN_106;
  wire  T_2659;
  wire  GEN_107;
  wire [2:0] GEN_108;
  wire [2:0] GEN_109;
  wire  GEN_110;
  wire  T_2661;
  wire [2:0] GEN_111;
  wire [2:0] GEN_112;
  wire [2:0] GEN_113;
  wire  T_2662;
  wire [2:0] GEN_114;
  wire [6:0] GEN_28;
  reg [31:0] GEN_164;
  wire [63:0] GEN_37;
  reg [63:0] GEN_165;
  RRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_prv(arb_io_in_0_bits_prv),
    .io_in_0_bits_pum(arb_io_in_0_bits_pum),
    .io_in_0_bits_mxr(arb_io_in_0_bits_mxr),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_store(arb_io_in_0_bits_store),
    .io_in_0_bits_fetch(arb_io_in_0_bits_fetch),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_prv(arb_io_in_1_bits_prv),
    .io_in_1_bits_pum(arb_io_in_1_bits_pum),
    .io_in_1_bits_mxr(arb_io_in_1_bits_mxr),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_store(arb_io_in_1_bits_store),
    .io_in_1_bits_fetch(arb_io_in_1_bits_fetch),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_prv(arb_io_out_bits_prv),
    .io_out_bits_pum(arb_io_out_bits_pum),
    .io_out_bits_mxr(arb_io_out_bits_mxr),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_store(arb_io_out_bits_store),
    .io_out_bits_fetch(arb_io_out_bits_fetch),
    .io_chosen(arb_io_chosen)
  );
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_0_resp_valid = T_2581;
  assign io_requestor_0_resp_bits_pte_reserved_for_hardware = r_pte_reserved_for_hardware;
  assign io_requestor_0_resp_bits_pte_ppn = T_2591;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign io_requestor_0_resp_bits_pte_a = r_pte_a;
  assign io_requestor_0_resp_bits_pte_g = r_pte_g;
  assign io_requestor_0_resp_bits_pte_u = r_pte_u;
  assign io_requestor_0_resp_bits_pte_x = r_pte_x;
  assign io_requestor_0_resp_bits_pte_w = r_pte_w;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign io_requestor_0_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_0_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_debug = io_dpath_status_debug;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_mxr = io_dpath_status_mxr;
  assign io_requestor_0_status_pum = io_dpath_status_pum;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_mpp = io_dpath_status_mpp;
  assign io_requestor_0_status_hpp = io_dpath_status_hpp;
  assign io_requestor_0_status_spp = io_dpath_status_spp;
  assign io_requestor_0_status_mpie = io_dpath_status_mpie;
  assign io_requestor_0_status_hpie = io_dpath_status_hpie;
  assign io_requestor_0_status_spie = io_dpath_status_spie;
  assign io_requestor_0_status_upie = io_dpath_status_upie;
  assign io_requestor_0_status_mie = io_dpath_status_mie;
  assign io_requestor_0_status_hie = io_dpath_status_hie;
  assign io_requestor_0_status_sie = io_dpath_status_sie;
  assign io_requestor_0_status_uie = io_dpath_status_uie;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  assign io_requestor_1_resp_valid = T_2595;
  assign io_requestor_1_resp_bits_pte_reserved_for_hardware = r_pte_reserved_for_hardware;
  assign io_requestor_1_resp_bits_pte_ppn = T_2591;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_a = r_pte_a;
  assign io_requestor_1_resp_bits_pte_g = r_pte_g;
  assign io_requestor_1_resp_bits_pte_u = r_pte_u;
  assign io_requestor_1_resp_bits_pte_x = r_pte_x;
  assign io_requestor_1_resp_bits_pte_w = r_pte_w;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_1_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_debug = io_dpath_status_debug;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_mxr = io_dpath_status_mxr;
  assign io_requestor_1_status_pum = io_dpath_status_pum;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_mpp = io_dpath_status_mpp;
  assign io_requestor_1_status_hpp = io_dpath_status_hpp;
  assign io_requestor_1_status_spp = io_dpath_status_spp;
  assign io_requestor_1_status_mpie = io_dpath_status_mpie;
  assign io_requestor_1_status_hpie = io_dpath_status_hpie;
  assign io_requestor_1_status_spie = io_dpath_status_spie;
  assign io_requestor_1_status_upie = io_dpath_status_upie;
  assign io_requestor_1_status_mie = io_dpath_status_mie;
  assign io_requestor_1_status_hie = io_dpath_status_hie;
  assign io_requestor_1_status_sie = io_dpath_status_sie;
  assign io_requestor_1_status_uie = io_dpath_status_uie;
  assign io_mem_req_valid = T_2558;
  assign io_mem_req_bits_addr = pte_addr[39:0];
  assign io_mem_req_bits_tag = GEN_28;
  assign io_mem_req_bits_cmd = T_2561;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_data = GEN_37;
  assign io_mem_s1_kill = s1_kill;
  assign io_mem_s1_data = T_2572;
  assign io_mem_invalidate_lr = 1'h0;
  assign T_2185 = r_req_addr[26:18];
  assign T_2186 = r_req_addr[26:9];
  assign vpn_idxs_1 = T_2186[8:0];
  assign vpn_idxs_2 = r_req_addr[8:0];
  assign T_2189 = count & 2'h1;
  assign T_2191 = count >= 2'h2;
  assign T_2195 = T_2189 >= 2'h1;
  assign T_2196 = T_2195 ? vpn_idxs_1 : T_2185;
  assign vpn_idx = T_2191 ? vpn_idxs_2 : T_2196;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_requestor_0_req_valid;
  assign arb_io_in_0_bits_prv = io_requestor_0_req_bits_prv;
  assign arb_io_in_0_bits_pum = io_requestor_0_req_bits_pum;
  assign arb_io_in_0_bits_mxr = io_requestor_0_req_bits_mxr;
  assign arb_io_in_0_bits_addr = io_requestor_0_req_bits_addr;
  assign arb_io_in_0_bits_store = io_requestor_0_req_bits_store;
  assign arb_io_in_0_bits_fetch = io_requestor_0_req_bits_fetch;
  assign arb_io_in_1_valid = io_requestor_1_req_valid;
  assign arb_io_in_1_bits_prv = io_requestor_1_req_bits_prv;
  assign arb_io_in_1_bits_pum = io_requestor_1_req_bits_pum;
  assign arb_io_in_1_bits_mxr = io_requestor_1_req_bits_mxr;
  assign arb_io_in_1_bits_addr = io_requestor_1_req_bits_addr;
  assign arb_io_in_1_bits_store = io_requestor_1_req_bits_store;
  assign arb_io_in_1_bits_fetch = io_requestor_1_req_bits_fetch;
  assign arb_io_out_ready = T_2204;
  assign T_2204 = state == 3'h0;
  assign T_2229_reserved_for_hardware = T_2251;
  assign T_2229_ppn = T_2250;
  assign T_2229_reserved_for_software = T_2249;
  assign T_2229_d = T_2248;
  assign T_2229_a = T_2247;
  assign T_2229_g = T_2246;
  assign T_2229_u = T_2245;
  assign T_2229_x = T_2244;
  assign T_2229_w = T_2243;
  assign T_2229_r = T_2242;
  assign T_2229_v = T_2241;
  assign T_2241 = io_mem_resp_bits_data[0];
  assign T_2242 = io_mem_resp_bits_data[1];
  assign T_2243 = io_mem_resp_bits_data[2];
  assign T_2244 = io_mem_resp_bits_data[3];
  assign T_2245 = io_mem_resp_bits_data[4];
  assign T_2246 = io_mem_resp_bits_data[5];
  assign T_2247 = io_mem_resp_bits_data[6];
  assign T_2248 = io_mem_resp_bits_data[7];
  assign T_2249 = io_mem_resp_bits_data[9:8];
  assign T_2250 = io_mem_resp_bits_data[47:10];
  assign T_2251 = io_mem_resp_bits_data[63:48];
  assign T_2276_reserved_for_hardware = T_2251;
  assign T_2276_ppn = T_2250;
  assign T_2276_reserved_for_software = T_2249;
  assign T_2276_d = T_2248;
  assign T_2276_a = T_2247;
  assign T_2276_g = T_2246;
  assign T_2276_u = T_2245;
  assign T_2276_x = T_2244;
  assign T_2276_w = T_2243;
  assign T_2276_r = T_2242;
  assign T_2276_v = T_2241;
  assign pte_reserved_for_hardware = T_2276_reserved_for_hardware;
  assign pte_ppn = {{18'd0}, T_2310};
  assign pte_reserved_for_software = T_2276_reserved_for_software;
  assign pte_d = T_2276_d;
  assign pte_a = T_2276_a;
  assign pte_g = T_2276_g;
  assign pte_u = T_2276_u;
  assign pte_x = T_2276_x;
  assign pte_w = T_2276_w;
  assign pte_r = T_2276_r;
  assign pte_v = GEN_2;
  assign T_2310 = T_2229_ppn[19:0];
  assign T_2311 = T_2229_ppn[37:20];
  assign T_2313 = T_2311 != 18'h0;
  assign GEN_2 = T_2313 ? 1'h0 : T_2276_v;
  assign T_2315 = {r_pte_ppn,vpn_idx};
  assign GEN_115 = {{3'd0}, T_2315};
  assign pte_addr = GEN_115 << 3;
  assign T_2316 = arb_io_out_ready & arb_io_out_valid;
  assign GEN_3 = T_2316 ? arb_io_out_bits_prv : r_req_prv;
  assign GEN_4 = T_2316 ? arb_io_out_bits_pum : r_req_pum;
  assign GEN_5 = T_2316 ? arb_io_out_bits_mxr : r_req_mxr;
  assign GEN_6 = T_2316 ? arb_io_out_bits_addr : r_req_addr;
  assign GEN_7 = T_2316 ? arb_io_out_bits_store : r_req_store;
  assign GEN_8 = T_2316 ? arb_io_out_bits_fetch : r_req_fetch;
  assign GEN_9 = T_2316 ? arb_io_chosen : r_req_dest;
  assign GEN_10 = T_2316 ? io_dpath_ptbr_ppn : r_pte_ppn;
  assign GEN_116 = {{18'd0}, T_2327_0};
  assign T_2337 = GEN_116 == pte_addr;
  assign GEN_117 = {{18'd0}, T_2327_1};
  assign T_2338 = GEN_117 == pte_addr;
  assign GEN_118 = {{18'd0}, T_2327_2};
  assign T_2339 = GEN_118 == pte_addr;
  assign GEN_119 = {{18'd0}, T_2327_3};
  assign T_2340 = GEN_119 == pte_addr;
  assign GEN_120 = {{18'd0}, T_2327_4};
  assign T_2341 = GEN_120 == pte_addr;
  assign GEN_121 = {{18'd0}, T_2327_5};
  assign T_2342 = GEN_121 == pte_addr;
  assign GEN_122 = {{18'd0}, T_2327_6};
  assign T_2343 = GEN_122 == pte_addr;
  assign GEN_123 = {{18'd0}, T_2327_7};
  assign T_2344 = GEN_123 == pte_addr;
  assign T_2345 = {T_2338,T_2337};
  assign T_2346 = {T_2340,T_2339};
  assign T_2347 = {T_2346,T_2345};
  assign T_2348 = {T_2342,T_2341};
  assign T_2349 = {T_2344,T_2343};
  assign T_2350 = {T_2349,T_2348};
  assign T_2351 = {T_2350,T_2347};
  assign T_2352 = T_2351 & T_2320;
  assign T_2354 = T_2352 != 8'h0;
  assign T_2356 = pte_r == 1'h0;
  assign T_2357 = pte_v & T_2356;
  assign T_2359 = pte_w == 1'h0;
  assign T_2360 = T_2357 & T_2359;
  assign T_2362 = pte_x == 1'h0;
  assign T_2363 = T_2360 & T_2362;
  assign T_2364 = io_mem_resp_valid & T_2363;
  assign T_2366 = T_2354 == 1'h0;
  assign T_2367 = T_2364 & T_2366;
  assign T_2368 = ~ T_2320;
  assign T_2370 = T_2368 == 8'h0;
  assign T_2372 = T_2318 >> 1'h1;
  assign T_2373 = T_2372[0];
  assign T_2374 = {1'h1,T_2373};
  assign T_2375 = T_2318 >> T_2374;
  assign T_2376 = T_2375[0];
  assign T_2377 = {T_2374,T_2376};
  assign T_2378 = T_2318 >> T_2377;
  assign T_2379 = T_2378[0];
  assign T_2380 = {T_2377,T_2379};
  assign T_2381 = T_2380[2:0];
  assign T_2383 = T_2368[0];
  assign T_2384 = T_2368[1];
  assign T_2385 = T_2368[2];
  assign T_2386 = T_2368[3];
  assign T_2387 = T_2368[4];
  assign T_2388 = T_2368[5];
  assign T_2389 = T_2368[6];
  assign T_2399 = T_2389 ? 3'h6 : 3'h7;
  assign T_2400 = T_2388 ? 3'h5 : T_2399;
  assign T_2401 = T_2387 ? 3'h4 : T_2400;
  assign T_2402 = T_2386 ? 3'h3 : T_2401;
  assign T_2403 = T_2385 ? 3'h2 : T_2402;
  assign T_2404 = T_2384 ? 3'h1 : T_2403;
  assign T_2405 = T_2383 ? 3'h0 : T_2404;
  assign T_2406 = T_2370 ? T_2381 : T_2405;
  assign T_2408 = 8'h1 << T_2406;
  assign T_2409 = T_2320 | T_2408;
  assign GEN_0 = pte_addr[31:0];
  assign GEN_11 = 3'h0 == T_2406 ? GEN_0 : T_2327_0;
  assign GEN_12 = 3'h1 == T_2406 ? GEN_0 : T_2327_1;
  assign GEN_13 = 3'h2 == T_2406 ? GEN_0 : T_2327_2;
  assign GEN_14 = 3'h3 == T_2406 ? GEN_0 : T_2327_3;
  assign GEN_15 = 3'h4 == T_2406 ? GEN_0 : T_2327_4;
  assign GEN_16 = 3'h5 == T_2406 ? GEN_0 : T_2327_5;
  assign GEN_17 = 3'h6 == T_2406 ? GEN_0 : T_2327_6;
  assign GEN_18 = 3'h7 == T_2406 ? GEN_0 : T_2327_7;
  assign GEN_1 = pte_ppn[19:0];
  assign GEN_19 = 3'h0 == T_2406 ? GEN_1 : T_2335_0;
  assign GEN_20 = 3'h1 == T_2406 ? GEN_1 : T_2335_1;
  assign GEN_21 = 3'h2 == T_2406 ? GEN_1 : T_2335_2;
  assign GEN_22 = 3'h3 == T_2406 ? GEN_1 : T_2335_3;
  assign GEN_23 = 3'h4 == T_2406 ? GEN_1 : T_2335_4;
  assign GEN_24 = 3'h5 == T_2406 ? GEN_1 : T_2335_5;
  assign GEN_25 = 3'h6 == T_2406 ? GEN_1 : T_2335_6;
  assign GEN_26 = 3'h7 == T_2406 ? GEN_1 : T_2335_7;
  assign GEN_27 = T_2367 ? T_2409 : T_2320;
  assign GEN_29 = T_2367 ? GEN_11 : T_2327_0;
  assign GEN_30 = T_2367 ? GEN_12 : T_2327_1;
  assign GEN_31 = T_2367 ? GEN_13 : T_2327_2;
  assign GEN_32 = T_2367 ? GEN_14 : T_2327_3;
  assign GEN_33 = T_2367 ? GEN_15 : T_2327_4;
  assign GEN_34 = T_2367 ? GEN_16 : T_2327_5;
  assign GEN_35 = T_2367 ? GEN_17 : T_2327_6;
  assign GEN_36 = T_2367 ? GEN_18 : T_2327_7;
  assign GEN_38 = T_2367 ? GEN_19 : T_2335_0;
  assign GEN_39 = T_2367 ? GEN_20 : T_2335_1;
  assign GEN_40 = T_2367 ? GEN_21 : T_2335_2;
  assign GEN_41 = T_2367 ? GEN_22 : T_2335_3;
  assign GEN_42 = T_2367 ? GEN_23 : T_2335_4;
  assign GEN_43 = T_2367 ? GEN_24 : T_2335_5;
  assign GEN_44 = T_2367 ? GEN_25 : T_2335_6;
  assign GEN_45 = T_2367 ? GEN_26 : T_2335_7;
  assign T_2410 = state == 3'h1;
  assign T_2411 = T_2354 & T_2410;
  assign T_2412 = T_2352[7:4];
  assign T_2413 = T_2352[3:0];
  assign T_2415 = T_2412 != 4'h0;
  assign T_2416 = T_2412 | T_2413;
  assign T_2417 = T_2416[3:2];
  assign T_2418 = T_2416[1:0];
  assign T_2420 = T_2417 != 2'h0;
  assign T_2421 = T_2417 | T_2418;
  assign T_2422 = T_2421[1];
  assign T_2423 = {T_2420,T_2422};
  assign T_2424 = {T_2415,T_2423};
  assign T_2426 = T_2424[2];
  assign T_2428 = T_2426 == 1'h0;
  assign T_2430 = 2'h1 << 1'h1;
  assign GEN_124 = {{6'd0}, T_2430};
  assign T_2431 = T_2318 | GEN_124;
  assign T_2432 = ~ T_2318;
  assign T_2433 = T_2432 | GEN_124;
  assign T_2434 = ~ T_2433;
  assign T_2435 = T_2428 ? T_2431 : T_2434;
  assign T_2436 = {1'h1,T_2426};
  assign T_2437 = T_2424[1];
  assign T_2439 = T_2437 == 1'h0;
  assign T_2441 = 4'h1 << T_2436;
  assign GEN_126 = {{4'd0}, T_2441};
  assign T_2442 = T_2435 | GEN_126;
  assign T_2443 = ~ T_2435;
  assign T_2444 = T_2443 | GEN_126;
  assign T_2445 = ~ T_2444;
  assign T_2446 = T_2439 ? T_2442 : T_2445;
  assign T_2447 = {T_2436,T_2437};
  assign T_2448 = T_2424[0];
  assign T_2450 = T_2448 == 1'h0;
  assign T_2452 = 8'h1 << T_2447;
  assign T_2453 = T_2446 | T_2452;
  assign T_2454 = ~ T_2446;
  assign T_2455 = T_2454 | T_2452;
  assign T_2456 = ~ T_2455;
  assign T_2457 = T_2450 ? T_2453 : T_2456;
  assign GEN_46 = T_2411 ? T_2457 : T_2318;
  assign GEN_47 = io_dpath_invalidate ? 8'h0 : GEN_27;
  assign T_2461 = count < 2'h2;
  assign pte_cache_hit = T_2354 & T_2461;
  assign T_2462 = T_2352[0];
  assign T_2463 = T_2352[1];
  assign T_2464 = T_2352[2];
  assign T_2465 = T_2352[3];
  assign T_2466 = T_2352[4];
  assign T_2467 = T_2352[5];
  assign T_2468 = T_2352[6];
  assign T_2469 = T_2352[7];
  assign T_2471 = T_2462 ? T_2335_0 : 20'h0;
  assign T_2473 = T_2463 ? T_2335_1 : 20'h0;
  assign T_2475 = T_2464 ? T_2335_2 : 20'h0;
  assign T_2477 = T_2465 ? T_2335_3 : 20'h0;
  assign T_2479 = T_2466 ? T_2335_4 : 20'h0;
  assign T_2481 = T_2467 ? T_2335_5 : 20'h0;
  assign T_2483 = T_2468 ? T_2335_6 : 20'h0;
  assign T_2485 = T_2469 ? T_2335_7 : 20'h0;
  assign T_2487 = T_2471 | T_2473;
  assign T_2488 = T_2487 | T_2475;
  assign T_2489 = T_2488 | T_2477;
  assign T_2490 = T_2489 | T_2479;
  assign T_2491 = T_2490 | T_2481;
  assign T_2492 = T_2491 | T_2483;
  assign T_2493 = T_2492 | T_2485;
  assign pte_cache_data = T_2493;
  assign T_2519_reserved_for_hardware = T_2543;
  assign T_2519_ppn = T_2542;
  assign T_2519_reserved_for_software = T_2541;
  assign T_2519_d = T_2540;
  assign T_2519_a = T_2539;
  assign T_2519_g = T_2538;
  assign T_2519_u = T_2537;
  assign T_2519_x = T_2536;
  assign T_2519_w = T_2535;
  assign T_2519_r = T_2534;
  assign T_2519_v = T_2533;
  assign T_2532 = 64'h0;
  assign T_2533 = T_2532[0];
  assign T_2534 = T_2532[1];
  assign T_2535 = T_2532[2];
  assign T_2536 = T_2532[3];
  assign T_2537 = T_2532[4];
  assign T_2538 = T_2532[5];
  assign T_2539 = T_2532[6];
  assign T_2540 = T_2532[7];
  assign T_2541 = T_2532[9:8];
  assign T_2542 = T_2532[47:10];
  assign T_2543 = T_2532[63:48];
  assign pte_wdata_reserved_for_hardware = T_2519_reserved_for_hardware;
  assign pte_wdata_ppn = T_2519_ppn;
  assign pte_wdata_reserved_for_software = T_2519_reserved_for_software;
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_a = 1'h1;
  assign pte_wdata_g = T_2519_g;
  assign pte_wdata_u = T_2519_u;
  assign pte_wdata_x = T_2519_x;
  assign pte_wdata_w = T_2519_w;
  assign pte_wdata_r = T_2519_r;
  assign pte_wdata_v = T_2519_v;
  assign T_2557 = state == 3'h4;
  assign T_2558 = T_2410 | T_2557;
  assign T_2561 = T_2557 ? 5'ha : 5'h0;
  assign T_2563 = {pte_wdata_r,pte_wdata_v};
  assign T_2564 = {pte_wdata_u,pte_wdata_x};
  assign T_2565 = {T_2564,pte_wdata_w};
  assign T_2566 = {T_2565,T_2563};
  assign T_2567 = {pte_wdata_d,pte_wdata_a};
  assign T_2568 = {T_2567,pte_wdata_g};
  assign T_2569 = {pte_wdata_reserved_for_hardware,pte_wdata_ppn};
  assign T_2570 = {T_2569,pte_wdata_reserved_for_software};
  assign T_2571 = {T_2570,T_2568};
  assign T_2572 = {T_2571,T_2566};
  assign T_2574 = pte_addr[49:30];
  assign T_2575 = r_req_addr[17:0];
  assign resp_ppns_0 = {T_2574,T_2575};
  assign T_2576 = pte_addr[49:21];
  assign resp_ppns_1 = {T_2576,vpn_idxs_2};
  assign resp_ppns_2 = pte_addr[49:12];
  assign T_2578 = state == 3'h7;
  assign T_2580 = r_req_dest == 1'h0;
  assign T_2581 = T_2578 & T_2580;
  assign T_2590 = T_2195 ? resp_ppns_1 : resp_ppns_0;
  assign T_2591 = T_2191 ? resp_ppns_2 : T_2590;
  assign T_2595 = T_2578 & r_req_dest;
  assign T_2606 = 3'h0 == state;
  assign GEN_48 = arb_io_out_valid ? 3'h1 : state;
  assign GEN_49 = T_2606 ? GEN_48 : state;
  assign GEN_50 = T_2606 ? 2'h0 : count;
  assign T_2608 = 3'h1 == state;
  assign T_2611 = count + 2'h1;
  assign T_2612 = T_2611[1:0];
  assign GEN_52 = pte_cache_hit ? 3'h1 : GEN_49;
  assign GEN_53 = pte_cache_hit ? T_2612 : GEN_50;
  assign GEN_54 = pte_cache_hit ? {{18'd0}, pte_cache_data} : GEN_10;
  assign T_2614 = pte_cache_hit == 1'h0;
  assign T_2615 = T_2614 & io_mem_req_ready;
  assign GEN_55 = T_2615 ? 3'h2 : GEN_52;
  assign GEN_56 = T_2608 ? pte_cache_hit : 1'h0;
  assign GEN_57 = T_2608 ? GEN_55 : GEN_49;
  assign GEN_58 = T_2608 ? GEN_53 : GEN_50;
  assign GEN_59 = T_2608 ? GEN_54 : GEN_10;
  assign T_2616 = 3'h2 == state;
  assign GEN_60 = io_mem_xcpt_pf_ld ? 1'h0 : r_pte_v;
  assign GEN_61 = io_mem_xcpt_pf_ld ? 3'h7 : 3'h3;
  assign GEN_62 = T_2616 ? GEN_61 : GEN_57;
  assign GEN_63 = T_2616 ? GEN_60 : r_pte_v;
  assign T_2618 = 3'h3 == state;
  assign GEN_64 = io_mem_s2_nack ? 3'h1 : GEN_62;
  assign T_2619 = pte_x & r_req_mxr;
  assign T_2620 = pte_r | T_2619;
  assign T_2621 = r_req_store ? pte_w : T_2620;
  assign T_2622 = r_req_fetch ? pte_x : T_2621;
  assign T_2624 = r_req_pum == 1'h0;
  assign T_2625 = r_req_prv[0];
  assign T_2626 = pte_u ? T_2624 : T_2625;
  assign T_2629 = pte_x & T_2359;
  assign T_2630 = pte_r | T_2629;
  assign T_2631 = pte_v & T_2630;
  assign T_2632 = T_2631 & T_2626;
  assign T_2633 = T_2632 & T_2622;
  assign T_2635 = pte_a == 1'h0;
  assign T_2637 = pte_d == 1'h0;
  assign T_2638 = r_req_store & T_2637;
  assign T_2639 = T_2635 | T_2638;
  assign T_2640 = T_2633 & T_2639;
  assign GEN_65 = T_2640 ? 3'h4 : 3'h7;
  assign T_2642 = T_2640 == 1'h0;
  assign GEN_66 = T_2642 ? pte_reserved_for_hardware : r_pte_reserved_for_hardware;
  assign GEN_67 = T_2642 ? pte_ppn : GEN_59;
  assign GEN_68 = T_2642 ? pte_reserved_for_software : r_pte_reserved_for_software;
  assign GEN_69 = T_2642 ? pte_d : r_pte_d;
  assign GEN_70 = T_2642 ? pte_a : r_pte_a;
  assign GEN_71 = T_2642 ? pte_g : r_pte_g;
  assign GEN_72 = T_2642 ? pte_u : r_pte_u;
  assign GEN_73 = T_2642 ? pte_x : r_pte_x;
  assign GEN_74 = T_2642 ? pte_w : r_pte_w;
  assign GEN_75 = T_2642 ? pte_r : r_pte_r;
  assign GEN_76 = T_2642 ? pte_v : GEN_63;
  assign T_2654 = T_2363 & T_2461;
  assign GEN_77 = T_2654 ? 3'h1 : GEN_65;
  assign GEN_78 = T_2654 ? T_2612 : GEN_58;
  assign GEN_79 = io_mem_resp_valid ? GEN_77 : GEN_64;
  assign GEN_80 = io_mem_resp_valid ? GEN_66 : r_pte_reserved_for_hardware;
  assign GEN_81 = io_mem_resp_valid ? GEN_67 : GEN_59;
  assign GEN_82 = io_mem_resp_valid ? GEN_68 : r_pte_reserved_for_software;
  assign GEN_83 = io_mem_resp_valid ? GEN_69 : r_pte_d;
  assign GEN_84 = io_mem_resp_valid ? GEN_70 : r_pte_a;
  assign GEN_85 = io_mem_resp_valid ? GEN_71 : r_pte_g;
  assign GEN_86 = io_mem_resp_valid ? GEN_72 : r_pte_u;
  assign GEN_87 = io_mem_resp_valid ? GEN_73 : r_pte_x;
  assign GEN_88 = io_mem_resp_valid ? GEN_74 : r_pte_w;
  assign GEN_89 = io_mem_resp_valid ? GEN_75 : r_pte_r;
  assign GEN_90 = io_mem_resp_valid ? GEN_76 : GEN_63;
  assign GEN_91 = io_mem_resp_valid ? GEN_78 : GEN_58;
  assign GEN_92 = T_2618 ? GEN_79 : GEN_62;
  assign GEN_93 = T_2618 ? GEN_80 : r_pte_reserved_for_hardware;
  assign GEN_94 = T_2618 ? GEN_81 : GEN_59;
  assign GEN_95 = T_2618 ? GEN_82 : r_pte_reserved_for_software;
  assign GEN_96 = T_2618 ? GEN_83 : r_pte_d;
  assign GEN_97 = T_2618 ? GEN_84 : r_pte_a;
  assign GEN_98 = T_2618 ? GEN_85 : r_pte_g;
  assign GEN_99 = T_2618 ? GEN_86 : r_pte_u;
  assign GEN_100 = T_2618 ? GEN_87 : r_pte_x;
  assign GEN_101 = T_2618 ? GEN_88 : r_pte_w;
  assign GEN_102 = T_2618 ? GEN_89 : r_pte_r;
  assign GEN_103 = T_2618 ? GEN_90 : GEN_63;
  assign GEN_104 = T_2618 ? GEN_91 : GEN_58;
  assign T_2658 = 3'h4 == state;
  assign GEN_105 = io_mem_req_ready ? 3'h5 : GEN_92;
  assign GEN_106 = T_2658 ? GEN_105 : GEN_92;
  assign T_2659 = 3'h5 == state;
  assign GEN_107 = io_mem_xcpt_pf_st ? 1'h0 : GEN_103;
  assign GEN_108 = io_mem_xcpt_pf_st ? 3'h7 : 3'h6;
  assign GEN_109 = T_2659 ? GEN_108 : GEN_106;
  assign GEN_110 = T_2659 ? GEN_107 : GEN_103;
  assign T_2661 = 3'h6 == state;
  assign GEN_111 = io_mem_s2_nack ? 3'h4 : GEN_109;
  assign GEN_112 = io_mem_resp_valid ? 3'h1 : GEN_111;
  assign GEN_113 = T_2661 ? GEN_112 : GEN_109;
  assign T_2662 = 3'h7 == state;
  assign GEN_114 = T_2662 ? 3'h0 : GEN_113;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_28 = GEN_164[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_165[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  state = GEN_51[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  count = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {1{$random}};
  s1_kill = GEN_127[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {1{$random}};
  r_req_prv = GEN_128[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {1{$random}};
  r_req_pum = GEN_129[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {1{$random}};
  r_req_mxr = GEN_130[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  r_req_addr = GEN_131[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  r_req_store = GEN_132[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  r_req_fetch = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  r_req_dest = GEN_134[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  r_pte_reserved_for_hardware = GEN_135[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {2{$random}};
  r_pte_ppn = GEN_136[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  r_pte_reserved_for_software = GEN_137[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  r_pte_d = GEN_138[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  r_pte_a = GEN_139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  r_pte_g = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  r_pte_u = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  r_pte_x = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  r_pte_w = GEN_143[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  r_pte_r = GEN_144[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  r_pte_v = GEN_145[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  T_2318 = GEN_146[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  T_2320 = GEN_147[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {1{$random}};
  T_2327_0 = GEN_148[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  T_2327_1 = GEN_149[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  T_2327_2 = GEN_150[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  T_2327_3 = GEN_151[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  T_2327_4 = GEN_152[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  T_2327_5 = GEN_153[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  T_2327_6 = GEN_154[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  T_2327_7 = GEN_155[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  T_2335_0 = GEN_156[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  T_2335_1 = GEN_157[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  T_2335_2 = GEN_158[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  T_2335_3 = GEN_159[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {1{$random}};
  T_2335_4 = GEN_160[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  T_2335_5 = GEN_161[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {1{$random}};
  T_2335_6 = GEN_162[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {1{$random}};
  T_2335_7 = GEN_163[19:0];
  `endif
  GEN_164 = {1{$random}};
  GEN_165 = {2{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_2662) begin
        state <= 3'h0;
      end else begin
        if(T_2661) begin
          if(io_mem_resp_valid) begin
            state <= 3'h1;
          end else begin
            if(io_mem_s2_nack) begin
              state <= 3'h4;
            end else begin
              if(T_2659) begin
                if(io_mem_xcpt_pf_st) begin
                  state <= 3'h7;
                end else begin
                  state <= 3'h6;
                end
              end else begin
                if(T_2658) begin
                  if(io_mem_req_ready) begin
                    state <= 3'h5;
                  end else begin
                    if(T_2618) begin
                      if(io_mem_resp_valid) begin
                        if(T_2654) begin
                          state <= 3'h1;
                        end else begin
                          if(T_2640) begin
                            state <= 3'h4;
                          end else begin
                            state <= 3'h7;
                          end
                        end
                      end else begin
                        if(io_mem_s2_nack) begin
                          state <= 3'h1;
                        end else begin
                          if(T_2616) begin
                            if(io_mem_xcpt_pf_ld) begin
                              state <= 3'h7;
                            end else begin
                              state <= 3'h3;
                            end
                          end else begin
                            if(T_2608) begin
                              if(T_2615) begin
                                state <= 3'h2;
                              end else begin
                                if(pte_cache_hit) begin
                                  state <= 3'h1;
                                end else begin
                                  if(T_2606) begin
                                    if(arb_io_out_valid) begin
                                      state <= 3'h1;
                                    end
                                  end
                                end
                              end
                            end else begin
                              if(T_2606) begin
                                if(arb_io_out_valid) begin
                                  state <= 3'h1;
                                end
                              end
                            end
                          end
                        end
                      end
                    end else begin
                      if(T_2616) begin
                        if(io_mem_xcpt_pf_ld) begin
                          state <= 3'h7;
                        end else begin
                          state <= 3'h3;
                        end
                      end else begin
                        if(T_2608) begin
                          if(T_2615) begin
                            state <= 3'h2;
                          end else begin
                            if(pte_cache_hit) begin
                              state <= 3'h1;
                            end else begin
                              if(T_2606) begin
                                if(arb_io_out_valid) begin
                                  state <= 3'h1;
                                end
                              end
                            end
                          end
                        end else begin
                          if(T_2606) begin
                            if(arb_io_out_valid) begin
                              state <= 3'h1;
                            end
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if(T_2618) begin
                    if(io_mem_resp_valid) begin
                      if(T_2654) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2640) begin
                          state <= 3'h4;
                        end else begin
                          state <= 3'h7;
                        end
                      end
                    end else begin
                      if(io_mem_s2_nack) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2616) begin
                          if(io_mem_xcpt_pf_ld) begin
                            state <= 3'h7;
                          end else begin
                            state <= 3'h3;
                          end
                        end else begin
                          if(T_2608) begin
                            if(T_2615) begin
                              state <= 3'h2;
                            end else begin
                              if(pte_cache_hit) begin
                                state <= 3'h1;
                              end else begin
                                state <= GEN_49;
                              end
                            end
                          end else begin
                            state <= GEN_49;
                          end
                        end
                      end
                    end
                  end else begin
                    if(T_2616) begin
                      if(io_mem_xcpt_pf_ld) begin
                        state <= 3'h7;
                      end else begin
                        state <= 3'h3;
                      end
                    end else begin
                      if(T_2608) begin
                        if(T_2615) begin
                          state <= 3'h2;
                        end else begin
                          if(pte_cache_hit) begin
                            state <= 3'h1;
                          end else begin
                            state <= GEN_49;
                          end
                        end
                      end else begin
                        state <= GEN_49;
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if(T_2659) begin
            if(io_mem_xcpt_pf_st) begin
              state <= 3'h7;
            end else begin
              state <= 3'h6;
            end
          end else begin
            if(T_2658) begin
              if(io_mem_req_ready) begin
                state <= 3'h5;
              end else begin
                if(T_2618) begin
                  if(io_mem_resp_valid) begin
                    if(T_2654) begin
                      state <= 3'h1;
                    end else begin
                      if(T_2640) begin
                        state <= 3'h4;
                      end else begin
                        state <= 3'h7;
                      end
                    end
                  end else begin
                    if(io_mem_s2_nack) begin
                      state <= 3'h1;
                    end else begin
                      state <= GEN_62;
                    end
                  end
                end else begin
                  state <= GEN_62;
                end
              end
            end else begin
              if(T_2618) begin
                if(io_mem_resp_valid) begin
                  if(T_2654) begin
                    state <= 3'h1;
                  end else begin
                    if(T_2640) begin
                      state <= 3'h4;
                    end else begin
                      state <= 3'h7;
                    end
                  end
                end else begin
                  if(io_mem_s2_nack) begin
                    state <= 3'h1;
                  end else begin
                    state <= GEN_62;
                  end
                end
              end else begin
                state <= GEN_62;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2654) begin
            count <= T_2612;
          end else begin
            if(T_2608) begin
              if(pte_cache_hit) begin
                count <= T_2612;
              end else begin
                if(T_2606) begin
                  count <= 2'h0;
                end
              end
            end else begin
              if(T_2606) begin
                count <= 2'h0;
              end
            end
          end
        end else begin
          if(T_2608) begin
            if(pte_cache_hit) begin
              count <= T_2612;
            end else begin
              if(T_2606) begin
                count <= 2'h0;
              end
            end
          end else begin
            if(T_2606) begin
              count <= 2'h0;
            end
          end
        end
      end else begin
        if(T_2608) begin
          if(pte_cache_hit) begin
            count <= T_2612;
          end else begin
            count <= GEN_50;
          end
        end else begin
          count <= GEN_50;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2608) begin
        s1_kill <= pte_cache_hit;
      end else begin
        s1_kill <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_prv <= arb_io_out_bits_prv;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_pum <= arb_io_out_bits_pum;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_mxr <= arb_io_out_bits_mxr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_addr <= arb_io_out_bits_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_store <= arb_io_out_bits_store;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_fetch <= arb_io_out_bits_fetch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2316) begin
        r_req_dest <= arb_io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_reserved_for_hardware <= pte_reserved_for_hardware;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_ppn <= pte_ppn;
          end else begin
            if(T_2608) begin
              if(pte_cache_hit) begin
                r_pte_ppn <= {{18'd0}, pte_cache_data};
              end else begin
                if(T_2316) begin
                  r_pte_ppn <= io_dpath_ptbr_ppn;
                end
              end
            end else begin
              if(T_2316) begin
                r_pte_ppn <= io_dpath_ptbr_ppn;
              end
            end
          end
        end else begin
          if(T_2608) begin
            if(pte_cache_hit) begin
              r_pte_ppn <= {{18'd0}, pte_cache_data};
            end else begin
              if(T_2316) begin
                r_pte_ppn <= io_dpath_ptbr_ppn;
              end
            end
          end else begin
            if(T_2316) begin
              r_pte_ppn <= io_dpath_ptbr_ppn;
            end
          end
        end
      end else begin
        if(T_2608) begin
          if(pte_cache_hit) begin
            r_pte_ppn <= {{18'd0}, pte_cache_data};
          end else begin
            r_pte_ppn <= GEN_10;
          end
        end else begin
          r_pte_ppn <= GEN_10;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_reserved_for_software <= pte_reserved_for_software;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_d <= pte_d;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_a <= pte_a;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_g <= pte_g;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_u <= pte_u;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_x <= pte_x;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_w <= pte_w;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2618) begin
        if(io_mem_resp_valid) begin
          if(T_2642) begin
            r_pte_r <= pte_r;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2659) begin
        if(io_mem_xcpt_pf_st) begin
          r_pte_v <= 1'h0;
        end else begin
          if(T_2618) begin
            if(io_mem_resp_valid) begin
              if(T_2642) begin
                r_pte_v <= pte_v;
              end else begin
                if(T_2616) begin
                  if(io_mem_xcpt_pf_ld) begin
                    r_pte_v <= 1'h0;
                  end
                end
              end
            end else begin
              if(T_2616) begin
                if(io_mem_xcpt_pf_ld) begin
                  r_pte_v <= 1'h0;
                end
              end
            end
          end else begin
            if(T_2616) begin
              if(io_mem_xcpt_pf_ld) begin
                r_pte_v <= 1'h0;
              end
            end
          end
        end
      end else begin
        if(T_2618) begin
          if(io_mem_resp_valid) begin
            if(T_2642) begin
              r_pte_v <= pte_v;
            end else begin
              if(T_2616) begin
                if(io_mem_xcpt_pf_ld) begin
                  r_pte_v <= 1'h0;
                end
              end
            end
          end else begin
            r_pte_v <= GEN_63;
          end
        end else begin
          r_pte_v <= GEN_63;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2411) begin
        if(T_2450) begin
          T_2318 <= T_2453;
        end else begin
          T_2318 <= T_2456;
        end
      end
    end
    if(reset) begin
      T_2320 <= 8'h0;
    end else begin
      if(io_dpath_invalidate) begin
        T_2320 <= 8'h0;
      end else begin
        if(T_2367) begin
          T_2320 <= T_2409;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h0 == T_2406) begin
          T_2327_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h1 == T_2406) begin
          T_2327_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h2 == T_2406) begin
          T_2327_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h3 == T_2406) begin
          T_2327_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h4 == T_2406) begin
          T_2327_4 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h5 == T_2406) begin
          T_2327_5 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h6 == T_2406) begin
          T_2327_6 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h7 == T_2406) begin
          T_2327_7 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h0 == T_2406) begin
          T_2335_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h1 == T_2406) begin
          T_2335_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h2 == T_2406) begin
          T_2335_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h3 == T_2406) begin
          T_2335_3 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h4 == T_2406) begin
          T_2335_4 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h5 == T_2406) begin
          T_2335_5 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h6 == T_2406) begin
          T_2335_6 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2367) begin
        if(3'h7 == T_2406) begin
          T_2335_7 <= GEN_1;
        end
      end
    end
  end
endmodule
module HellaCacheArbiter(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input  [6:0] io_requestor_0_req_bits_tag,
  input  [4:0] io_requestor_0_req_bits_cmd,
  input  [2:0] io_requestor_0_req_bits_typ,
  input   io_requestor_0_req_bits_phys,
  input  [63:0] io_requestor_0_req_bits_data,
  input   io_requestor_0_s1_kill,
  input  [63:0] io_requestor_0_s1_data,
  output  io_requestor_0_s2_nack,
  output  io_requestor_0_resp_valid,
  output [39:0] io_requestor_0_resp_bits_addr,
  output [6:0] io_requestor_0_resp_bits_tag,
  output [4:0] io_requestor_0_resp_bits_cmd,
  output [2:0] io_requestor_0_resp_bits_typ,
  output [63:0] io_requestor_0_resp_bits_data,
  output  io_requestor_0_resp_bits_replay,
  output  io_requestor_0_resp_bits_has_data,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output [63:0] io_requestor_0_resp_bits_store_data,
  output  io_requestor_0_replay_next,
  output  io_requestor_0_xcpt_ma_ld,
  output  io_requestor_0_xcpt_ma_st,
  output  io_requestor_0_xcpt_pf_ld,
  output  io_requestor_0_xcpt_pf_st,
  input   io_requestor_0_invalidate_lr,
  output  io_requestor_0_ordered,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [6:0] io_requestor_1_req_bits_tag,
  input  [4:0] io_requestor_1_req_bits_cmd,
  input  [2:0] io_requestor_1_req_bits_typ,
  input   io_requestor_1_req_bits_phys,
  input  [63:0] io_requestor_1_req_bits_data,
  input   io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data,
  output  io_requestor_1_s2_nack,
  output  io_requestor_1_resp_valid,
  output [39:0] io_requestor_1_resp_bits_addr,
  output [6:0] io_requestor_1_resp_bits_tag,
  output [4:0] io_requestor_1_resp_bits_cmd,
  output [2:0] io_requestor_1_resp_bits_typ,
  output [63:0] io_requestor_1_resp_bits_data,
  output  io_requestor_1_resp_bits_replay,
  output  io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output [63:0] io_requestor_1_resp_bits_store_data,
  output  io_requestor_1_replay_next,
  output  io_requestor_1_xcpt_ma_ld,
  output  io_requestor_1_xcpt_ma_st,
  output  io_requestor_1_xcpt_pf_ld,
  output  io_requestor_1_xcpt_pf_st,
  input   io_requestor_1_invalidate_lr,
  output  io_requestor_1_ordered,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [6:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered
);
  reg  T_6368;
  reg [31:0] GEN_9;
  reg  T_6369;
  reg [31:0] GEN_10;
  wire  T_6370;
  wire  T_6371;
  wire  T_6373;
  wire  T_6374;
  wire [7:0] T_6376;
  wire [7:0] T_6379;
  wire [4:0] GEN_0;
  wire [2:0] GEN_1;
  wire [39:0] GEN_2;
  wire  GEN_3;
  wire [7:0] GEN_4;
  wire  GEN_5;
  wire  T_6382;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire  T_6383;
  wire  T_6385;
  wire  T_6386;
  wire  T_6388;
  wire  T_6389;
  wire [5:0] T_6390;
  wire  T_6394;
  wire  T_6397;
  wire [63:0] GEN_8;
  reg [63:0] GEN_11;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = T_6389;
  assign io_requestor_0_resp_valid = T_6386;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_tag = {{1'd0}, T_6390};
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_replay_next = io_mem_replay_next;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_1_req_ready = T_6374;
  assign io_requestor_1_s2_nack = T_6397;
  assign io_requestor_1_resp_valid = T_6394;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_tag = {{1'd0}, T_6390};
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_replay_next = io_mem_replay_next;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_mem_req_valid = T_6371;
  assign io_mem_req_bits_addr = GEN_2;
  assign io_mem_req_bits_tag = GEN_4[6:0];
  assign io_mem_req_bits_cmd = GEN_0;
  assign io_mem_req_bits_typ = GEN_1;
  assign io_mem_req_bits_phys = GEN_3;
  assign io_mem_req_bits_data = GEN_8;
  assign io_mem_s1_kill = GEN_6;
  assign io_mem_s1_data = GEN_7;
  assign io_mem_invalidate_lr = T_6370;
  assign T_6370 = io_requestor_0_invalidate_lr | io_requestor_1_invalidate_lr;
  assign T_6371 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign T_6373 = io_requestor_0_req_valid == 1'h0;
  assign T_6374 = io_requestor_0_req_ready & T_6373;
  assign T_6376 = {io_requestor_1_req_bits_tag,1'h1};
  assign T_6379 = {io_requestor_0_req_bits_tag,1'h0};
  assign GEN_0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign GEN_1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign GEN_2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign GEN_3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign GEN_4 = io_requestor_0_req_valid ? T_6379 : T_6376;
  assign GEN_5 = io_requestor_0_req_valid ? 1'h0 : 1'h1;
  assign T_6382 = T_6368 == 1'h0;
  assign GEN_6 = T_6382 ? io_requestor_0_s1_kill : io_requestor_1_s1_kill;
  assign GEN_7 = T_6382 ? io_requestor_0_s1_data : io_requestor_1_s1_data;
  assign T_6383 = io_mem_resp_bits_tag[0];
  assign T_6385 = T_6383 == 1'h0;
  assign T_6386 = io_mem_resp_valid & T_6385;
  assign T_6388 = T_6369 == 1'h0;
  assign T_6389 = io_mem_s2_nack & T_6388;
  assign T_6390 = io_mem_resp_bits_tag[6:1];
  assign T_6394 = io_mem_resp_valid & T_6383;
  assign T_6397 = io_mem_s2_nack & T_6369;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_11[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  T_6368 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  T_6369 = GEN_10[0:0];
  `endif
  GEN_11 = {2{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_requestor_0_req_valid) begin
        T_6368 <= 1'h0;
      end else begin
        T_6368 <= 1'h1;
      end
    end
    if(1'h0) begin
    end else begin
      T_6369 <= T_6368;
    end
  end
endmodule
module RocketTile(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output [1:0] io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [10:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output [1:0] io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input  [1:0] io_cached_0_grant_bits_client_xact_id,
  input  [2:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [2:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output [1:0] io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [10:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input  [1:0] io_uncached_0_grant_bits_client_xact_id,
  input  [2:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip
);
  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [39:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire  core_io_imem_resp_bits_btb_valid;
  wire  core_io_imem_resp_bits_btb_bits_taken;
  wire [1:0] core_io_imem_resp_bits_btb_bits_mask;
  wire  core_io_imem_resp_bits_btb_bits_bridx;
  wire [38:0] core_io_imem_resp_bits_btb_bits_target;
  wire [5:0] core_io_imem_resp_bits_btb_bits_entry;
  wire [6:0] core_io_imem_resp_bits_btb_bits_bht_history;
  wire [1:0] core_io_imem_resp_bits_btb_bits_bht_value;
  wire [39:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data;
  wire [1:0] core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_btb_update_bits_pc;
  wire [38:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isValid;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [38:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [38:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [39:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [39:0] core_io_dmem_req_bits_addr;
  wire [6:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [63:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [63:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [39:0] core_io_dmem_resp_bits_addr;
  wire [6:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [63:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [63:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [6:0] core_io_ptw_ptbr_asid;
  wire [37:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [3:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [63:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [63:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] core_io_rocc_cmd_bits_rs1;
  wire [63:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_cmd_bits_status_debug;
  wire [1:0] core_io_rocc_cmd_bits_status_prv;
  wire  core_io_rocc_cmd_bits_status_sd;
  wire [30:0] core_io_rocc_cmd_bits_status_zero3;
  wire  core_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] core_io_rocc_cmd_bits_status_zero2;
  wire [4:0] core_io_rocc_cmd_bits_status_vm;
  wire [3:0] core_io_rocc_cmd_bits_status_zero1;
  wire  core_io_rocc_cmd_bits_status_mxr;
  wire  core_io_rocc_cmd_bits_status_pum;
  wire  core_io_rocc_cmd_bits_status_mprv;
  wire [1:0] core_io_rocc_cmd_bits_status_xs;
  wire [1:0] core_io_rocc_cmd_bits_status_fs;
  wire [1:0] core_io_rocc_cmd_bits_status_mpp;
  wire [1:0] core_io_rocc_cmd_bits_status_hpp;
  wire  core_io_rocc_cmd_bits_status_spp;
  wire  core_io_rocc_cmd_bits_status_mpie;
  wire  core_io_rocc_cmd_bits_status_hpie;
  wire  core_io_rocc_cmd_bits_status_spie;
  wire  core_io_rocc_cmd_bits_status_upie;
  wire  core_io_rocc_cmd_bits_status_mie;
  wire  core_io_rocc_cmd_bits_status_hie;
  wire  core_io_rocc_cmd_bits_status_sie;
  wire  core_io_rocc_cmd_bits_status_uie;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [63:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [39:0] core_io_rocc_mem_req_bits_addr;
  wire [6:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [63:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [63:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [39:0] core_io_rocc_mem_resp_bits_addr;
  wire [6:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [63:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [63:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [10:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] core_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [39:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_req_bits_speculative;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire  icache_io_cpu_resp_bits_btb_valid;
  wire  icache_io_cpu_resp_bits_btb_bits_taken;
  wire [1:0] icache_io_cpu_resp_bits_btb_bits_mask;
  wire  icache_io_cpu_resp_bits_btb_bits_bridx;
  wire [38:0] icache_io_cpu_resp_bits_btb_bits_target;
  wire [5:0] icache_io_cpu_resp_bits_btb_bits_entry;
  wire [6:0] icache_io_cpu_resp_bits_btb_bits_bht_history;
  wire [1:0] icache_io_cpu_resp_bits_btb_bits_bht_value;
  wire [39:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data;
  wire [1:0] icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_resp_bits_replay;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_btb_update_bits_pc;
  wire [38:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isValid;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [38:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [38:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [39:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_pum;
  wire  icache_io_ptw_req_bits_mxr;
  wire [26:0] icache_io_ptw_req_bits_addr;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [15:0] icache_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [1:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_a;
  wire  icache_io_ptw_resp_bits_pte_g;
  wire  icache_io_ptw_resp_bits_pte_u;
  wire  icache_io_ptw_resp_bits_pte_x;
  wire  icache_io_ptw_resp_bits_pte_w;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire [6:0] icache_io_ptw_ptbr_asid;
  wire [37:0] icache_io_ptw_ptbr_ppn;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [3:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_mxr;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [10:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  HellaCache_1_clk;
  wire  HellaCache_1_reset;
  wire  HellaCache_1_io_cpu_req_ready;
  wire  HellaCache_1_io_cpu_req_valid;
  wire [39:0] HellaCache_1_io_cpu_req_bits_addr;
  wire [6:0] HellaCache_1_io_cpu_req_bits_tag;
  wire [4:0] HellaCache_1_io_cpu_req_bits_cmd;
  wire [2:0] HellaCache_1_io_cpu_req_bits_typ;
  wire  HellaCache_1_io_cpu_req_bits_phys;
  wire [63:0] HellaCache_1_io_cpu_req_bits_data;
  wire  HellaCache_1_io_cpu_s1_kill;
  wire [63:0] HellaCache_1_io_cpu_s1_data;
  wire  HellaCache_1_io_cpu_s2_nack;
  wire  HellaCache_1_io_cpu_resp_valid;
  wire [39:0] HellaCache_1_io_cpu_resp_bits_addr;
  wire [6:0] HellaCache_1_io_cpu_resp_bits_tag;
  wire [4:0] HellaCache_1_io_cpu_resp_bits_cmd;
  wire [2:0] HellaCache_1_io_cpu_resp_bits_typ;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_data;
  wire  HellaCache_1_io_cpu_resp_bits_replay;
  wire  HellaCache_1_io_cpu_resp_bits_has_data;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_data_word_bypass;
  wire [63:0] HellaCache_1_io_cpu_resp_bits_store_data;
  wire  HellaCache_1_io_cpu_replay_next;
  wire  HellaCache_1_io_cpu_xcpt_ma_ld;
  wire  HellaCache_1_io_cpu_xcpt_ma_st;
  wire  HellaCache_1_io_cpu_xcpt_pf_ld;
  wire  HellaCache_1_io_cpu_xcpt_pf_st;
  wire  HellaCache_1_io_cpu_invalidate_lr;
  wire  HellaCache_1_io_cpu_ordered;
  wire  HellaCache_1_io_ptw_req_ready;
  wire  HellaCache_1_io_ptw_req_valid;
  wire [1:0] HellaCache_1_io_ptw_req_bits_prv;
  wire  HellaCache_1_io_ptw_req_bits_pum;
  wire  HellaCache_1_io_ptw_req_bits_mxr;
  wire [26:0] HellaCache_1_io_ptw_req_bits_addr;
  wire  HellaCache_1_io_ptw_req_bits_store;
  wire  HellaCache_1_io_ptw_req_bits_fetch;
  wire  HellaCache_1_io_ptw_resp_valid;
  wire [15:0] HellaCache_1_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] HellaCache_1_io_ptw_resp_bits_pte_ppn;
  wire [1:0] HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software;
  wire  HellaCache_1_io_ptw_resp_bits_pte_d;
  wire  HellaCache_1_io_ptw_resp_bits_pte_a;
  wire  HellaCache_1_io_ptw_resp_bits_pte_g;
  wire  HellaCache_1_io_ptw_resp_bits_pte_u;
  wire  HellaCache_1_io_ptw_resp_bits_pte_x;
  wire  HellaCache_1_io_ptw_resp_bits_pte_w;
  wire  HellaCache_1_io_ptw_resp_bits_pte_r;
  wire  HellaCache_1_io_ptw_resp_bits_pte_v;
  wire [6:0] HellaCache_1_io_ptw_ptbr_asid;
  wire [37:0] HellaCache_1_io_ptw_ptbr_ppn;
  wire  HellaCache_1_io_ptw_invalidate;
  wire  HellaCache_1_io_ptw_status_debug;
  wire [1:0] HellaCache_1_io_ptw_status_prv;
  wire  HellaCache_1_io_ptw_status_sd;
  wire [30:0] HellaCache_1_io_ptw_status_zero3;
  wire  HellaCache_1_io_ptw_status_sd_rv32;
  wire [1:0] HellaCache_1_io_ptw_status_zero2;
  wire [4:0] HellaCache_1_io_ptw_status_vm;
  wire [3:0] HellaCache_1_io_ptw_status_zero1;
  wire  HellaCache_1_io_ptw_status_mxr;
  wire  HellaCache_1_io_ptw_status_pum;
  wire  HellaCache_1_io_ptw_status_mprv;
  wire [1:0] HellaCache_1_io_ptw_status_xs;
  wire [1:0] HellaCache_1_io_ptw_status_fs;
  wire [1:0] HellaCache_1_io_ptw_status_mpp;
  wire [1:0] HellaCache_1_io_ptw_status_hpp;
  wire  HellaCache_1_io_ptw_status_spp;
  wire  HellaCache_1_io_ptw_status_mpie;
  wire  HellaCache_1_io_ptw_status_hpie;
  wire  HellaCache_1_io_ptw_status_spie;
  wire  HellaCache_1_io_ptw_status_upie;
  wire  HellaCache_1_io_ptw_status_mie;
  wire  HellaCache_1_io_ptw_status_hie;
  wire  HellaCache_1_io_ptw_status_sie;
  wire  HellaCache_1_io_ptw_status_uie;
  wire  HellaCache_1_io_mem_acquire_ready;
  wire  HellaCache_1_io_mem_acquire_valid;
  wire [25:0] HellaCache_1_io_mem_acquire_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_acquire_bits_client_xact_id;
  wire [2:0] HellaCache_1_io_mem_acquire_bits_addr_beat;
  wire  HellaCache_1_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] HellaCache_1_io_mem_acquire_bits_a_type;
  wire [10:0] HellaCache_1_io_mem_acquire_bits_union;
  wire [63:0] HellaCache_1_io_mem_acquire_bits_data;
  wire  HellaCache_1_io_mem_probe_ready;
  wire  HellaCache_1_io_mem_probe_valid;
  wire [25:0] HellaCache_1_io_mem_probe_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_probe_bits_p_type;
  wire  HellaCache_1_io_mem_release_ready;
  wire  HellaCache_1_io_mem_release_valid;
  wire [2:0] HellaCache_1_io_mem_release_bits_addr_beat;
  wire [25:0] HellaCache_1_io_mem_release_bits_addr_block;
  wire [1:0] HellaCache_1_io_mem_release_bits_client_xact_id;
  wire  HellaCache_1_io_mem_release_bits_voluntary;
  wire [2:0] HellaCache_1_io_mem_release_bits_r_type;
  wire [63:0] HellaCache_1_io_mem_release_bits_data;
  wire  HellaCache_1_io_mem_grant_ready;
  wire  HellaCache_1_io_mem_grant_valid;
  wire [2:0] HellaCache_1_io_mem_grant_bits_addr_beat;
  wire [1:0] HellaCache_1_io_mem_grant_bits_client_xact_id;
  wire [2:0] HellaCache_1_io_mem_grant_bits_manager_xact_id;
  wire  HellaCache_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] HellaCache_1_io_mem_grant_bits_g_type;
  wire [63:0] HellaCache_1_io_mem_grant_bits_data;
  wire  HellaCache_1_io_mem_grant_bits_manager_id;
  wire  HellaCache_1_io_mem_finish_ready;
  wire  HellaCache_1_io_mem_finish_valid;
  wire [2:0] HellaCache_1_io_mem_finish_bits_manager_xact_id;
  wire  HellaCache_1_io_mem_finish_bits_manager_id;
  wire  fpuOpt_clk;
  wire  fpuOpt_reset;
  wire [31:0] fpuOpt_io_inst;
  wire [63:0] fpuOpt_io_fromint_data;
  wire [2:0] fpuOpt_io_fcsr_rm;
  wire  fpuOpt_io_fcsr_flags_valid;
  wire [4:0] fpuOpt_io_fcsr_flags_bits;
  wire [63:0] fpuOpt_io_store_data;
  wire [63:0] fpuOpt_io_toint_data;
  wire  fpuOpt_io_dmem_resp_val;
  wire [2:0] fpuOpt_io_dmem_resp_type;
  wire [4:0] fpuOpt_io_dmem_resp_tag;
  wire [63:0] fpuOpt_io_dmem_resp_data;
  wire  fpuOpt_io_valid;
  wire  fpuOpt_io_fcsr_rdy;
  wire  fpuOpt_io_nack_mem;
  wire  fpuOpt_io_illegal_rm;
  wire  fpuOpt_io_killx;
  wire  fpuOpt_io_killm;
  wire [4:0] fpuOpt_io_dec_cmd;
  wire  fpuOpt_io_dec_ldst;
  wire  fpuOpt_io_dec_wen;
  wire  fpuOpt_io_dec_ren1;
  wire  fpuOpt_io_dec_ren2;
  wire  fpuOpt_io_dec_ren3;
  wire  fpuOpt_io_dec_swap12;
  wire  fpuOpt_io_dec_swap23;
  wire  fpuOpt_io_dec_single;
  wire  fpuOpt_io_dec_fromint;
  wire  fpuOpt_io_dec_toint;
  wire  fpuOpt_io_dec_fastpipe;
  wire  fpuOpt_io_dec_fma;
  wire  fpuOpt_io_dec_div;
  wire  fpuOpt_io_dec_sqrt;
  wire  fpuOpt_io_dec_round;
  wire  fpuOpt_io_dec_wflags;
  wire  fpuOpt_io_sboard_set;
  wire  fpuOpt_io_sboard_clr;
  wire [4:0] fpuOpt_io_sboard_clra;
  wire  fpuOpt_io_cp_req_ready;
  wire  fpuOpt_io_cp_req_valid;
  wire [4:0] fpuOpt_io_cp_req_bits_cmd;
  wire  fpuOpt_io_cp_req_bits_ldst;
  wire  fpuOpt_io_cp_req_bits_wen;
  wire  fpuOpt_io_cp_req_bits_ren1;
  wire  fpuOpt_io_cp_req_bits_ren2;
  wire  fpuOpt_io_cp_req_bits_ren3;
  wire  fpuOpt_io_cp_req_bits_swap12;
  wire  fpuOpt_io_cp_req_bits_swap23;
  wire  fpuOpt_io_cp_req_bits_single;
  wire  fpuOpt_io_cp_req_bits_fromint;
  wire  fpuOpt_io_cp_req_bits_toint;
  wire  fpuOpt_io_cp_req_bits_fastpipe;
  wire  fpuOpt_io_cp_req_bits_fma;
  wire  fpuOpt_io_cp_req_bits_div;
  wire  fpuOpt_io_cp_req_bits_sqrt;
  wire  fpuOpt_io_cp_req_bits_round;
  wire  fpuOpt_io_cp_req_bits_wflags;
  wire [2:0] fpuOpt_io_cp_req_bits_rm;
  wire [1:0] fpuOpt_io_cp_req_bits_typ;
  wire [64:0] fpuOpt_io_cp_req_bits_in1;
  wire [64:0] fpuOpt_io_cp_req_bits_in2;
  wire [64:0] fpuOpt_io_cp_req_bits_in3;
  wire  fpuOpt_io_cp_resp_ready;
  wire  fpuOpt_io_cp_resp_valid;
  wire [64:0] fpuOpt_io_cp_resp_bits_data;
  wire [4:0] fpuOpt_io_cp_resp_bits_exc;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [10:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [10:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_out_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  PTW_1_clk;
  wire  PTW_1_reset;
  wire  PTW_1_io_requestor_0_req_ready;
  wire  PTW_1_io_requestor_0_req_valid;
  wire [1:0] PTW_1_io_requestor_0_req_bits_prv;
  wire  PTW_1_io_requestor_0_req_bits_pum;
  wire  PTW_1_io_requestor_0_req_bits_mxr;
  wire [26:0] PTW_1_io_requestor_0_req_bits_addr;
  wire  PTW_1_io_requestor_0_req_bits_store;
  wire  PTW_1_io_requestor_0_req_bits_fetch;
  wire  PTW_1_io_requestor_0_resp_valid;
  wire [15:0] PTW_1_io_requestor_0_resp_bits_pte_reserved_for_hardware;
  wire [37:0] PTW_1_io_requestor_0_resp_bits_pte_ppn;
  wire [1:0] PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire  PTW_1_io_requestor_0_resp_bits_pte_d;
  wire  PTW_1_io_requestor_0_resp_bits_pte_a;
  wire  PTW_1_io_requestor_0_resp_bits_pte_g;
  wire  PTW_1_io_requestor_0_resp_bits_pte_u;
  wire  PTW_1_io_requestor_0_resp_bits_pte_x;
  wire  PTW_1_io_requestor_0_resp_bits_pte_w;
  wire  PTW_1_io_requestor_0_resp_bits_pte_r;
  wire  PTW_1_io_requestor_0_resp_bits_pte_v;
  wire [6:0] PTW_1_io_requestor_0_ptbr_asid;
  wire [37:0] PTW_1_io_requestor_0_ptbr_ppn;
  wire  PTW_1_io_requestor_0_invalidate;
  wire  PTW_1_io_requestor_0_status_debug;
  wire [1:0] PTW_1_io_requestor_0_status_prv;
  wire  PTW_1_io_requestor_0_status_sd;
  wire [30:0] PTW_1_io_requestor_0_status_zero3;
  wire  PTW_1_io_requestor_0_status_sd_rv32;
  wire [1:0] PTW_1_io_requestor_0_status_zero2;
  wire [4:0] PTW_1_io_requestor_0_status_vm;
  wire [3:0] PTW_1_io_requestor_0_status_zero1;
  wire  PTW_1_io_requestor_0_status_mxr;
  wire  PTW_1_io_requestor_0_status_pum;
  wire  PTW_1_io_requestor_0_status_mprv;
  wire [1:0] PTW_1_io_requestor_0_status_xs;
  wire [1:0] PTW_1_io_requestor_0_status_fs;
  wire [1:0] PTW_1_io_requestor_0_status_mpp;
  wire [1:0] PTW_1_io_requestor_0_status_hpp;
  wire  PTW_1_io_requestor_0_status_spp;
  wire  PTW_1_io_requestor_0_status_mpie;
  wire  PTW_1_io_requestor_0_status_hpie;
  wire  PTW_1_io_requestor_0_status_spie;
  wire  PTW_1_io_requestor_0_status_upie;
  wire  PTW_1_io_requestor_0_status_mie;
  wire  PTW_1_io_requestor_0_status_hie;
  wire  PTW_1_io_requestor_0_status_sie;
  wire  PTW_1_io_requestor_0_status_uie;
  wire  PTW_1_io_requestor_1_req_ready;
  wire  PTW_1_io_requestor_1_req_valid;
  wire [1:0] PTW_1_io_requestor_1_req_bits_prv;
  wire  PTW_1_io_requestor_1_req_bits_pum;
  wire  PTW_1_io_requestor_1_req_bits_mxr;
  wire [26:0] PTW_1_io_requestor_1_req_bits_addr;
  wire  PTW_1_io_requestor_1_req_bits_store;
  wire  PTW_1_io_requestor_1_req_bits_fetch;
  wire  PTW_1_io_requestor_1_resp_valid;
  wire [15:0] PTW_1_io_requestor_1_resp_bits_pte_reserved_for_hardware;
  wire [37:0] PTW_1_io_requestor_1_resp_bits_pte_ppn;
  wire [1:0] PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire  PTW_1_io_requestor_1_resp_bits_pte_d;
  wire  PTW_1_io_requestor_1_resp_bits_pte_a;
  wire  PTW_1_io_requestor_1_resp_bits_pte_g;
  wire  PTW_1_io_requestor_1_resp_bits_pte_u;
  wire  PTW_1_io_requestor_1_resp_bits_pte_x;
  wire  PTW_1_io_requestor_1_resp_bits_pte_w;
  wire  PTW_1_io_requestor_1_resp_bits_pte_r;
  wire  PTW_1_io_requestor_1_resp_bits_pte_v;
  wire [6:0] PTW_1_io_requestor_1_ptbr_asid;
  wire [37:0] PTW_1_io_requestor_1_ptbr_ppn;
  wire  PTW_1_io_requestor_1_invalidate;
  wire  PTW_1_io_requestor_1_status_debug;
  wire [1:0] PTW_1_io_requestor_1_status_prv;
  wire  PTW_1_io_requestor_1_status_sd;
  wire [30:0] PTW_1_io_requestor_1_status_zero3;
  wire  PTW_1_io_requestor_1_status_sd_rv32;
  wire [1:0] PTW_1_io_requestor_1_status_zero2;
  wire [4:0] PTW_1_io_requestor_1_status_vm;
  wire [3:0] PTW_1_io_requestor_1_status_zero1;
  wire  PTW_1_io_requestor_1_status_mxr;
  wire  PTW_1_io_requestor_1_status_pum;
  wire  PTW_1_io_requestor_1_status_mprv;
  wire [1:0] PTW_1_io_requestor_1_status_xs;
  wire [1:0] PTW_1_io_requestor_1_status_fs;
  wire [1:0] PTW_1_io_requestor_1_status_mpp;
  wire [1:0] PTW_1_io_requestor_1_status_hpp;
  wire  PTW_1_io_requestor_1_status_spp;
  wire  PTW_1_io_requestor_1_status_mpie;
  wire  PTW_1_io_requestor_1_status_hpie;
  wire  PTW_1_io_requestor_1_status_spie;
  wire  PTW_1_io_requestor_1_status_upie;
  wire  PTW_1_io_requestor_1_status_mie;
  wire  PTW_1_io_requestor_1_status_hie;
  wire  PTW_1_io_requestor_1_status_sie;
  wire  PTW_1_io_requestor_1_status_uie;
  wire  PTW_1_io_mem_req_ready;
  wire  PTW_1_io_mem_req_valid;
  wire [39:0] PTW_1_io_mem_req_bits_addr;
  wire [6:0] PTW_1_io_mem_req_bits_tag;
  wire [4:0] PTW_1_io_mem_req_bits_cmd;
  wire [2:0] PTW_1_io_mem_req_bits_typ;
  wire  PTW_1_io_mem_req_bits_phys;
  wire [63:0] PTW_1_io_mem_req_bits_data;
  wire  PTW_1_io_mem_s1_kill;
  wire [63:0] PTW_1_io_mem_s1_data;
  wire  PTW_1_io_mem_s2_nack;
  wire  PTW_1_io_mem_resp_valid;
  wire [39:0] PTW_1_io_mem_resp_bits_addr;
  wire [6:0] PTW_1_io_mem_resp_bits_tag;
  wire [4:0] PTW_1_io_mem_resp_bits_cmd;
  wire [2:0] PTW_1_io_mem_resp_bits_typ;
  wire [63:0] PTW_1_io_mem_resp_bits_data;
  wire  PTW_1_io_mem_resp_bits_replay;
  wire  PTW_1_io_mem_resp_bits_has_data;
  wire [63:0] PTW_1_io_mem_resp_bits_data_word_bypass;
  wire [63:0] PTW_1_io_mem_resp_bits_store_data;
  wire  PTW_1_io_mem_replay_next;
  wire  PTW_1_io_mem_xcpt_ma_ld;
  wire  PTW_1_io_mem_xcpt_ma_st;
  wire  PTW_1_io_mem_xcpt_pf_ld;
  wire  PTW_1_io_mem_xcpt_pf_st;
  wire  PTW_1_io_mem_invalidate_lr;
  wire  PTW_1_io_mem_ordered;
  wire [6:0] PTW_1_io_dpath_ptbr_asid;
  wire [37:0] PTW_1_io_dpath_ptbr_ppn;
  wire  PTW_1_io_dpath_invalidate;
  wire  PTW_1_io_dpath_status_debug;
  wire [1:0] PTW_1_io_dpath_status_prv;
  wire  PTW_1_io_dpath_status_sd;
  wire [30:0] PTW_1_io_dpath_status_zero3;
  wire  PTW_1_io_dpath_status_sd_rv32;
  wire [1:0] PTW_1_io_dpath_status_zero2;
  wire [4:0] PTW_1_io_dpath_status_vm;
  wire [3:0] PTW_1_io_dpath_status_zero1;
  wire  PTW_1_io_dpath_status_mxr;
  wire  PTW_1_io_dpath_status_pum;
  wire  PTW_1_io_dpath_status_mprv;
  wire [1:0] PTW_1_io_dpath_status_xs;
  wire [1:0] PTW_1_io_dpath_status_fs;
  wire [1:0] PTW_1_io_dpath_status_mpp;
  wire [1:0] PTW_1_io_dpath_status_hpp;
  wire  PTW_1_io_dpath_status_spp;
  wire  PTW_1_io_dpath_status_mpie;
  wire  PTW_1_io_dpath_status_hpie;
  wire  PTW_1_io_dpath_status_spie;
  wire  PTW_1_io_dpath_status_upie;
  wire  PTW_1_io_dpath_status_mie;
  wire  PTW_1_io_dpath_status_hie;
  wire  PTW_1_io_dpath_status_sie;
  wire  PTW_1_io_dpath_status_uie;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [39:0] dcArb_io_requestor_0_req_bits_addr;
  wire [6:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [63:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [63:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [6:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_requestor_1_req_ready;
  wire  dcArb_io_requestor_1_req_valid;
  wire [39:0] dcArb_io_requestor_1_req_bits_addr;
  wire [6:0] dcArb_io_requestor_1_req_bits_tag;
  wire [4:0] dcArb_io_requestor_1_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_req_bits_typ;
  wire  dcArb_io_requestor_1_req_bits_phys;
  wire [63:0] dcArb_io_requestor_1_req_bits_data;
  wire  dcArb_io_requestor_1_s1_kill;
  wire [63:0] dcArb_io_requestor_1_s1_data;
  wire  dcArb_io_requestor_1_s2_nack;
  wire  dcArb_io_requestor_1_resp_valid;
  wire [39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire [6:0] dcArb_io_requestor_1_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data;
  wire  dcArb_io_requestor_1_resp_bits_replay;
  wire  dcArb_io_requestor_1_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire  dcArb_io_requestor_1_replay_next;
  wire  dcArb_io_requestor_1_xcpt_ma_ld;
  wire  dcArb_io_requestor_1_xcpt_ma_st;
  wire  dcArb_io_requestor_1_xcpt_pf_ld;
  wire  dcArb_io_requestor_1_xcpt_pf_st;
  wire  dcArb_io_requestor_1_invalidate_lr;
  wire  dcArb_io_requestor_1_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [39:0] dcArb_io_mem_req_bits_addr;
  wire [6:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [63:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [63:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [39:0] dcArb_io_mem_resp_bits_addr;
  wire [6:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [63:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [63:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  wire  GEN_0;
  reg [31:0] GEN_49;
  wire  GEN_1;
  reg [31:0] GEN_50;
  wire [4:0] GEN_2;
  reg [31:0] GEN_51;
  wire [63:0] GEN_3;
  reg [63:0] GEN_52;
  wire  GEN_4;
  reg [31:0] GEN_53;
  wire [39:0] GEN_5;
  reg [63:0] GEN_54;
  wire [6:0] GEN_6;
  reg [31:0] GEN_55;
  wire [4:0] GEN_7;
  reg [31:0] GEN_56;
  wire [2:0] GEN_8;
  reg [31:0] GEN_57;
  wire  GEN_9;
  reg [31:0] GEN_58;
  wire [63:0] GEN_10;
  reg [63:0] GEN_59;
  wire  GEN_11;
  reg [31:0] GEN_60;
  wire [63:0] GEN_12;
  reg [63:0] GEN_61;
  wire  GEN_13;
  reg [31:0] GEN_62;
  wire  GEN_14;
  reg [31:0] GEN_63;
  wire  GEN_15;
  reg [31:0] GEN_64;
  wire  GEN_16;
  reg [31:0] GEN_65;
  wire [25:0] GEN_17;
  reg [31:0] GEN_66;
  wire [1:0] GEN_18;
  reg [31:0] GEN_67;
  wire [2:0] GEN_19;
  reg [31:0] GEN_68;
  wire  GEN_20;
  reg [31:0] GEN_69;
  wire [2:0] GEN_21;
  reg [31:0] GEN_70;
  wire [10:0] GEN_22;
  reg [31:0] GEN_71;
  wire [63:0] GEN_23;
  reg [63:0] GEN_72;
  wire  GEN_24;
  reg [31:0] GEN_73;
  wire  GEN_25;
  reg [31:0] GEN_74;
  wire [4:0] GEN_26;
  reg [31:0] GEN_75;
  wire  GEN_27;
  reg [31:0] GEN_76;
  wire  GEN_28;
  reg [31:0] GEN_77;
  wire  GEN_29;
  reg [31:0] GEN_78;
  wire  GEN_30;
  reg [31:0] GEN_79;
  wire  GEN_31;
  reg [31:0] GEN_80;
  wire  GEN_32;
  reg [31:0] GEN_81;
  wire  GEN_33;
  reg [31:0] GEN_82;
  wire  GEN_34;
  reg [31:0] GEN_83;
  wire  GEN_35;
  reg [31:0] GEN_84;
  wire  GEN_36;
  reg [31:0] GEN_85;
  wire  GEN_37;
  reg [31:0] GEN_86;
  wire  GEN_38;
  reg [31:0] GEN_87;
  wire  GEN_39;
  reg [31:0] GEN_88;
  wire  GEN_40;
  reg [31:0] GEN_89;
  wire  GEN_41;
  reg [31:0] GEN_90;
  wire  GEN_42;
  reg [31:0] GEN_91;
  wire [2:0] GEN_43;
  reg [31:0] GEN_92;
  wire [1:0] GEN_44;
  reg [31:0] GEN_93;
  wire [64:0] GEN_45;
  reg [95:0] GEN_94;
  wire [64:0] GEN_46;
  reg [95:0] GEN_95;
  wire [64:0] GEN_47;
  reg [95:0] GEN_96;
  wire  GEN_48;
  reg [31:0] GEN_97;
  Rocket core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_valid(core_io_imem_resp_bits_btb_valid),
    .io_imem_resp_bits_btb_bits_taken(core_io_imem_resp_bits_btb_bits_taken),
    .io_imem_resp_bits_btb_bits_mask(core_io_imem_resp_bits_btb_bits_mask),
    .io_imem_resp_bits_btb_bits_bridx(core_io_imem_resp_bits_btb_bits_bridx),
    .io_imem_resp_bits_btb_bits_target(core_io_imem_resp_bits_btb_bits_target),
    .io_imem_resp_bits_btb_bits_entry(core_io_imem_resp_bits_btb_bits_entry),
    .io_imem_resp_bits_btb_bits_bht_history(core_io_imem_resp_bits_btb_bits_bht_history),
    .io_imem_resp_bits_btb_bits_bht_value(core_io_imem_resp_bits_btb_bits_bht_value),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isValid(core_io_imem_btb_update_bits_isValid),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(core_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(core_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(core_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(core_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(core_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(core_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(core_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(core_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(core_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(core_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(core_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(core_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(core_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(core_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(core_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(core_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(core_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(core_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(core_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(core_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(core_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(core_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(core_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(core_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception)
  );
  Frontend icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(icache_io_cpu_req_bits_speculative),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_valid(icache_io_cpu_resp_bits_btb_valid),
    .io_cpu_resp_bits_btb_bits_taken(icache_io_cpu_resp_bits_btb_bits_taken),
    .io_cpu_resp_bits_btb_bits_mask(icache_io_cpu_resp_bits_btb_bits_mask),
    .io_cpu_resp_bits_btb_bits_bridx(icache_io_cpu_resp_bits_btb_bits_bridx),
    .io_cpu_resp_bits_btb_bits_target(icache_io_cpu_resp_bits_btb_bits_target),
    .io_cpu_resp_bits_btb_bits_entry(icache_io_cpu_resp_bits_btb_bits_entry),
    .io_cpu_resp_bits_btb_bits_bht_history(icache_io_cpu_resp_bits_btb_bits_bht_history),
    .io_cpu_resp_bits_btb_bits_bht_value(icache_io_cpu_resp_bits_btb_bits_bht_value),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(icache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_resp_bits_replay(icache_io_cpu_resp_bits_replay),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isValid(icache_io_cpu_btb_update_bits_isValid),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(icache_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(icache_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(icache_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(icache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(icache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(icache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(icache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(icache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(icache_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(icache_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_mxr(icache_io_ptw_status_mxr),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  HellaCache HellaCache_1 (
    .clk(HellaCache_1_clk),
    .reset(HellaCache_1_reset),
    .io_cpu_req_ready(HellaCache_1_io_cpu_req_ready),
    .io_cpu_req_valid(HellaCache_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(HellaCache_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(HellaCache_1_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(HellaCache_1_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(HellaCache_1_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(HellaCache_1_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(HellaCache_1_io_cpu_req_bits_data),
    .io_cpu_s1_kill(HellaCache_1_io_cpu_s1_kill),
    .io_cpu_s1_data(HellaCache_1_io_cpu_s1_data),
    .io_cpu_s2_nack(HellaCache_1_io_cpu_s2_nack),
    .io_cpu_resp_valid(HellaCache_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(HellaCache_1_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(HellaCache_1_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(HellaCache_1_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(HellaCache_1_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(HellaCache_1_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(HellaCache_1_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(HellaCache_1_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(HellaCache_1_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(HellaCache_1_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(HellaCache_1_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(HellaCache_1_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(HellaCache_1_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(HellaCache_1_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(HellaCache_1_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(HellaCache_1_io_cpu_invalidate_lr),
    .io_cpu_ordered(HellaCache_1_io_cpu_ordered),
    .io_ptw_req_ready(HellaCache_1_io_ptw_req_ready),
    .io_ptw_req_valid(HellaCache_1_io_ptw_req_valid),
    .io_ptw_req_bits_prv(HellaCache_1_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(HellaCache_1_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(HellaCache_1_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(HellaCache_1_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(HellaCache_1_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(HellaCache_1_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(HellaCache_1_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(HellaCache_1_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(HellaCache_1_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(HellaCache_1_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(HellaCache_1_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(HellaCache_1_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(HellaCache_1_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(HellaCache_1_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(HellaCache_1_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(HellaCache_1_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(HellaCache_1_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(HellaCache_1_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(HellaCache_1_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(HellaCache_1_io_ptw_invalidate),
    .io_ptw_status_debug(HellaCache_1_io_ptw_status_debug),
    .io_ptw_status_prv(HellaCache_1_io_ptw_status_prv),
    .io_ptw_status_sd(HellaCache_1_io_ptw_status_sd),
    .io_ptw_status_zero3(HellaCache_1_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(HellaCache_1_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(HellaCache_1_io_ptw_status_zero2),
    .io_ptw_status_vm(HellaCache_1_io_ptw_status_vm),
    .io_ptw_status_zero1(HellaCache_1_io_ptw_status_zero1),
    .io_ptw_status_mxr(HellaCache_1_io_ptw_status_mxr),
    .io_ptw_status_pum(HellaCache_1_io_ptw_status_pum),
    .io_ptw_status_mprv(HellaCache_1_io_ptw_status_mprv),
    .io_ptw_status_xs(HellaCache_1_io_ptw_status_xs),
    .io_ptw_status_fs(HellaCache_1_io_ptw_status_fs),
    .io_ptw_status_mpp(HellaCache_1_io_ptw_status_mpp),
    .io_ptw_status_hpp(HellaCache_1_io_ptw_status_hpp),
    .io_ptw_status_spp(HellaCache_1_io_ptw_status_spp),
    .io_ptw_status_mpie(HellaCache_1_io_ptw_status_mpie),
    .io_ptw_status_hpie(HellaCache_1_io_ptw_status_hpie),
    .io_ptw_status_spie(HellaCache_1_io_ptw_status_spie),
    .io_ptw_status_upie(HellaCache_1_io_ptw_status_upie),
    .io_ptw_status_mie(HellaCache_1_io_ptw_status_mie),
    .io_ptw_status_hie(HellaCache_1_io_ptw_status_hie),
    .io_ptw_status_sie(HellaCache_1_io_ptw_status_sie),
    .io_ptw_status_uie(HellaCache_1_io_ptw_status_uie),
    .io_mem_acquire_ready(HellaCache_1_io_mem_acquire_ready),
    .io_mem_acquire_valid(HellaCache_1_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(HellaCache_1_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(HellaCache_1_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(HellaCache_1_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(HellaCache_1_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(HellaCache_1_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(HellaCache_1_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(HellaCache_1_io_mem_acquire_bits_data),
    .io_mem_probe_ready(HellaCache_1_io_mem_probe_ready),
    .io_mem_probe_valid(HellaCache_1_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(HellaCache_1_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(HellaCache_1_io_mem_probe_bits_p_type),
    .io_mem_release_ready(HellaCache_1_io_mem_release_ready),
    .io_mem_release_valid(HellaCache_1_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(HellaCache_1_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(HellaCache_1_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(HellaCache_1_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(HellaCache_1_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(HellaCache_1_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(HellaCache_1_io_mem_release_bits_data),
    .io_mem_grant_ready(HellaCache_1_io_mem_grant_ready),
    .io_mem_grant_valid(HellaCache_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(HellaCache_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(HellaCache_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(HellaCache_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(HellaCache_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(HellaCache_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(HellaCache_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(HellaCache_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(HellaCache_1_io_mem_finish_ready),
    .io_mem_finish_valid(HellaCache_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(HellaCache_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(HellaCache_1_io_mem_finish_bits_manager_id)
  );
  FPU fpuOpt (
    .clk(fpuOpt_clk),
    .reset(fpuOpt_reset),
    .io_inst(fpuOpt_io_inst),
    .io_fromint_data(fpuOpt_io_fromint_data),
    .io_fcsr_rm(fpuOpt_io_fcsr_rm),
    .io_fcsr_flags_valid(fpuOpt_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(fpuOpt_io_fcsr_flags_bits),
    .io_store_data(fpuOpt_io_store_data),
    .io_toint_data(fpuOpt_io_toint_data),
    .io_dmem_resp_val(fpuOpt_io_dmem_resp_val),
    .io_dmem_resp_type(fpuOpt_io_dmem_resp_type),
    .io_dmem_resp_tag(fpuOpt_io_dmem_resp_tag),
    .io_dmem_resp_data(fpuOpt_io_dmem_resp_data),
    .io_valid(fpuOpt_io_valid),
    .io_fcsr_rdy(fpuOpt_io_fcsr_rdy),
    .io_nack_mem(fpuOpt_io_nack_mem),
    .io_illegal_rm(fpuOpt_io_illegal_rm),
    .io_killx(fpuOpt_io_killx),
    .io_killm(fpuOpt_io_killm),
    .io_dec_cmd(fpuOpt_io_dec_cmd),
    .io_dec_ldst(fpuOpt_io_dec_ldst),
    .io_dec_wen(fpuOpt_io_dec_wen),
    .io_dec_ren1(fpuOpt_io_dec_ren1),
    .io_dec_ren2(fpuOpt_io_dec_ren2),
    .io_dec_ren3(fpuOpt_io_dec_ren3),
    .io_dec_swap12(fpuOpt_io_dec_swap12),
    .io_dec_swap23(fpuOpt_io_dec_swap23),
    .io_dec_single(fpuOpt_io_dec_single),
    .io_dec_fromint(fpuOpt_io_dec_fromint),
    .io_dec_toint(fpuOpt_io_dec_toint),
    .io_dec_fastpipe(fpuOpt_io_dec_fastpipe),
    .io_dec_fma(fpuOpt_io_dec_fma),
    .io_dec_div(fpuOpt_io_dec_div),
    .io_dec_sqrt(fpuOpt_io_dec_sqrt),
    .io_dec_round(fpuOpt_io_dec_round),
    .io_dec_wflags(fpuOpt_io_dec_wflags),
    .io_sboard_set(fpuOpt_io_sboard_set),
    .io_sboard_clr(fpuOpt_io_sboard_clr),
    .io_sboard_clra(fpuOpt_io_sboard_clra),
    .io_cp_req_ready(fpuOpt_io_cp_req_ready),
    .io_cp_req_valid(fpuOpt_io_cp_req_valid),
    .io_cp_req_bits_cmd(fpuOpt_io_cp_req_bits_cmd),
    .io_cp_req_bits_ldst(fpuOpt_io_cp_req_bits_ldst),
    .io_cp_req_bits_wen(fpuOpt_io_cp_req_bits_wen),
    .io_cp_req_bits_ren1(fpuOpt_io_cp_req_bits_ren1),
    .io_cp_req_bits_ren2(fpuOpt_io_cp_req_bits_ren2),
    .io_cp_req_bits_ren3(fpuOpt_io_cp_req_bits_ren3),
    .io_cp_req_bits_swap12(fpuOpt_io_cp_req_bits_swap12),
    .io_cp_req_bits_swap23(fpuOpt_io_cp_req_bits_swap23),
    .io_cp_req_bits_single(fpuOpt_io_cp_req_bits_single),
    .io_cp_req_bits_fromint(fpuOpt_io_cp_req_bits_fromint),
    .io_cp_req_bits_toint(fpuOpt_io_cp_req_bits_toint),
    .io_cp_req_bits_fastpipe(fpuOpt_io_cp_req_bits_fastpipe),
    .io_cp_req_bits_fma(fpuOpt_io_cp_req_bits_fma),
    .io_cp_req_bits_div(fpuOpt_io_cp_req_bits_div),
    .io_cp_req_bits_sqrt(fpuOpt_io_cp_req_bits_sqrt),
    .io_cp_req_bits_round(fpuOpt_io_cp_req_bits_round),
    .io_cp_req_bits_wflags(fpuOpt_io_cp_req_bits_wflags),
    .io_cp_req_bits_rm(fpuOpt_io_cp_req_bits_rm),
    .io_cp_req_bits_typ(fpuOpt_io_cp_req_bits_typ),
    .io_cp_req_bits_in1(fpuOpt_io_cp_req_bits_in1),
    .io_cp_req_bits_in2(fpuOpt_io_cp_req_bits_in2),
    .io_cp_req_bits_in3(fpuOpt_io_cp_req_bits_in3),
    .io_cp_resp_ready(fpuOpt_io_cp_resp_ready),
    .io_cp_resp_valid(fpuOpt_io_cp_resp_valid),
    .io_cp_resp_bits_data(fpuOpt_io_cp_resp_bits_data),
    .io_cp_resp_bits_exc(fpuOpt_io_cp_resp_bits_exc)
  );
  ClientUncachedTileLinkIOArbiter uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  PTW PTW_1 (
    .clk(PTW_1_clk),
    .reset(PTW_1_reset),
    .io_requestor_0_req_ready(PTW_1_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(PTW_1_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_prv(PTW_1_io_requestor_0_req_bits_prv),
    .io_requestor_0_req_bits_pum(PTW_1_io_requestor_0_req_bits_pum),
    .io_requestor_0_req_bits_mxr(PTW_1_io_requestor_0_req_bits_mxr),
    .io_requestor_0_req_bits_addr(PTW_1_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_store(PTW_1_io_requestor_0_req_bits_store),
    .io_requestor_0_req_bits_fetch(PTW_1_io_requestor_0_req_bits_fetch),
    .io_requestor_0_resp_valid(PTW_1_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_pte_reserved_for_hardware(PTW_1_io_requestor_0_resp_bits_pte_reserved_for_hardware),
    .io_requestor_0_resp_bits_pte_ppn(PTW_1_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_reserved_for_software(PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software),
    .io_requestor_0_resp_bits_pte_d(PTW_1_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_a(PTW_1_io_requestor_0_resp_bits_pte_a),
    .io_requestor_0_resp_bits_pte_g(PTW_1_io_requestor_0_resp_bits_pte_g),
    .io_requestor_0_resp_bits_pte_u(PTW_1_io_requestor_0_resp_bits_pte_u),
    .io_requestor_0_resp_bits_pte_x(PTW_1_io_requestor_0_resp_bits_pte_x),
    .io_requestor_0_resp_bits_pte_w(PTW_1_io_requestor_0_resp_bits_pte_w),
    .io_requestor_0_resp_bits_pte_r(PTW_1_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_v(PTW_1_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_ptbr_asid(PTW_1_io_requestor_0_ptbr_asid),
    .io_requestor_0_ptbr_ppn(PTW_1_io_requestor_0_ptbr_ppn),
    .io_requestor_0_invalidate(PTW_1_io_requestor_0_invalidate),
    .io_requestor_0_status_debug(PTW_1_io_requestor_0_status_debug),
    .io_requestor_0_status_prv(PTW_1_io_requestor_0_status_prv),
    .io_requestor_0_status_sd(PTW_1_io_requestor_0_status_sd),
    .io_requestor_0_status_zero3(PTW_1_io_requestor_0_status_zero3),
    .io_requestor_0_status_sd_rv32(PTW_1_io_requestor_0_status_sd_rv32),
    .io_requestor_0_status_zero2(PTW_1_io_requestor_0_status_zero2),
    .io_requestor_0_status_vm(PTW_1_io_requestor_0_status_vm),
    .io_requestor_0_status_zero1(PTW_1_io_requestor_0_status_zero1),
    .io_requestor_0_status_mxr(PTW_1_io_requestor_0_status_mxr),
    .io_requestor_0_status_pum(PTW_1_io_requestor_0_status_pum),
    .io_requestor_0_status_mprv(PTW_1_io_requestor_0_status_mprv),
    .io_requestor_0_status_xs(PTW_1_io_requestor_0_status_xs),
    .io_requestor_0_status_fs(PTW_1_io_requestor_0_status_fs),
    .io_requestor_0_status_mpp(PTW_1_io_requestor_0_status_mpp),
    .io_requestor_0_status_hpp(PTW_1_io_requestor_0_status_hpp),
    .io_requestor_0_status_spp(PTW_1_io_requestor_0_status_spp),
    .io_requestor_0_status_mpie(PTW_1_io_requestor_0_status_mpie),
    .io_requestor_0_status_hpie(PTW_1_io_requestor_0_status_hpie),
    .io_requestor_0_status_spie(PTW_1_io_requestor_0_status_spie),
    .io_requestor_0_status_upie(PTW_1_io_requestor_0_status_upie),
    .io_requestor_0_status_mie(PTW_1_io_requestor_0_status_mie),
    .io_requestor_0_status_hie(PTW_1_io_requestor_0_status_hie),
    .io_requestor_0_status_sie(PTW_1_io_requestor_0_status_sie),
    .io_requestor_0_status_uie(PTW_1_io_requestor_0_status_uie),
    .io_requestor_1_req_ready(PTW_1_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(PTW_1_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_prv(PTW_1_io_requestor_1_req_bits_prv),
    .io_requestor_1_req_bits_pum(PTW_1_io_requestor_1_req_bits_pum),
    .io_requestor_1_req_bits_mxr(PTW_1_io_requestor_1_req_bits_mxr),
    .io_requestor_1_req_bits_addr(PTW_1_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_store(PTW_1_io_requestor_1_req_bits_store),
    .io_requestor_1_req_bits_fetch(PTW_1_io_requestor_1_req_bits_fetch),
    .io_requestor_1_resp_valid(PTW_1_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_pte_reserved_for_hardware(PTW_1_io_requestor_1_resp_bits_pte_reserved_for_hardware),
    .io_requestor_1_resp_bits_pte_ppn(PTW_1_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_reserved_for_software(PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software),
    .io_requestor_1_resp_bits_pte_d(PTW_1_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_a(PTW_1_io_requestor_1_resp_bits_pte_a),
    .io_requestor_1_resp_bits_pte_g(PTW_1_io_requestor_1_resp_bits_pte_g),
    .io_requestor_1_resp_bits_pte_u(PTW_1_io_requestor_1_resp_bits_pte_u),
    .io_requestor_1_resp_bits_pte_x(PTW_1_io_requestor_1_resp_bits_pte_x),
    .io_requestor_1_resp_bits_pte_w(PTW_1_io_requestor_1_resp_bits_pte_w),
    .io_requestor_1_resp_bits_pte_r(PTW_1_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_v(PTW_1_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_ptbr_asid(PTW_1_io_requestor_1_ptbr_asid),
    .io_requestor_1_ptbr_ppn(PTW_1_io_requestor_1_ptbr_ppn),
    .io_requestor_1_invalidate(PTW_1_io_requestor_1_invalidate),
    .io_requestor_1_status_debug(PTW_1_io_requestor_1_status_debug),
    .io_requestor_1_status_prv(PTW_1_io_requestor_1_status_prv),
    .io_requestor_1_status_sd(PTW_1_io_requestor_1_status_sd),
    .io_requestor_1_status_zero3(PTW_1_io_requestor_1_status_zero3),
    .io_requestor_1_status_sd_rv32(PTW_1_io_requestor_1_status_sd_rv32),
    .io_requestor_1_status_zero2(PTW_1_io_requestor_1_status_zero2),
    .io_requestor_1_status_vm(PTW_1_io_requestor_1_status_vm),
    .io_requestor_1_status_zero1(PTW_1_io_requestor_1_status_zero1),
    .io_requestor_1_status_mxr(PTW_1_io_requestor_1_status_mxr),
    .io_requestor_1_status_pum(PTW_1_io_requestor_1_status_pum),
    .io_requestor_1_status_mprv(PTW_1_io_requestor_1_status_mprv),
    .io_requestor_1_status_xs(PTW_1_io_requestor_1_status_xs),
    .io_requestor_1_status_fs(PTW_1_io_requestor_1_status_fs),
    .io_requestor_1_status_mpp(PTW_1_io_requestor_1_status_mpp),
    .io_requestor_1_status_hpp(PTW_1_io_requestor_1_status_hpp),
    .io_requestor_1_status_spp(PTW_1_io_requestor_1_status_spp),
    .io_requestor_1_status_mpie(PTW_1_io_requestor_1_status_mpie),
    .io_requestor_1_status_hpie(PTW_1_io_requestor_1_status_hpie),
    .io_requestor_1_status_spie(PTW_1_io_requestor_1_status_spie),
    .io_requestor_1_status_upie(PTW_1_io_requestor_1_status_upie),
    .io_requestor_1_status_mie(PTW_1_io_requestor_1_status_mie),
    .io_requestor_1_status_hie(PTW_1_io_requestor_1_status_hie),
    .io_requestor_1_status_sie(PTW_1_io_requestor_1_status_sie),
    .io_requestor_1_status_uie(PTW_1_io_requestor_1_status_uie),
    .io_mem_req_ready(PTW_1_io_mem_req_ready),
    .io_mem_req_valid(PTW_1_io_mem_req_valid),
    .io_mem_req_bits_addr(PTW_1_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(PTW_1_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(PTW_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(PTW_1_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(PTW_1_io_mem_req_bits_phys),
    .io_mem_req_bits_data(PTW_1_io_mem_req_bits_data),
    .io_mem_s1_kill(PTW_1_io_mem_s1_kill),
    .io_mem_s1_data(PTW_1_io_mem_s1_data),
    .io_mem_s2_nack(PTW_1_io_mem_s2_nack),
    .io_mem_resp_valid(PTW_1_io_mem_resp_valid),
    .io_mem_resp_bits_addr(PTW_1_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(PTW_1_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(PTW_1_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(PTW_1_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(PTW_1_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(PTW_1_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(PTW_1_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(PTW_1_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(PTW_1_io_mem_resp_bits_store_data),
    .io_mem_replay_next(PTW_1_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(PTW_1_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(PTW_1_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(PTW_1_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(PTW_1_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(PTW_1_io_mem_invalidate_lr),
    .io_mem_ordered(PTW_1_io_mem_ordered),
    .io_dpath_ptbr_asid(PTW_1_io_dpath_ptbr_asid),
    .io_dpath_ptbr_ppn(PTW_1_io_dpath_ptbr_ppn),
    .io_dpath_invalidate(PTW_1_io_dpath_invalidate),
    .io_dpath_status_debug(PTW_1_io_dpath_status_debug),
    .io_dpath_status_prv(PTW_1_io_dpath_status_prv),
    .io_dpath_status_sd(PTW_1_io_dpath_status_sd),
    .io_dpath_status_zero3(PTW_1_io_dpath_status_zero3),
    .io_dpath_status_sd_rv32(PTW_1_io_dpath_status_sd_rv32),
    .io_dpath_status_zero2(PTW_1_io_dpath_status_zero2),
    .io_dpath_status_vm(PTW_1_io_dpath_status_vm),
    .io_dpath_status_zero1(PTW_1_io_dpath_status_zero1),
    .io_dpath_status_mxr(PTW_1_io_dpath_status_mxr),
    .io_dpath_status_pum(PTW_1_io_dpath_status_pum),
    .io_dpath_status_mprv(PTW_1_io_dpath_status_mprv),
    .io_dpath_status_xs(PTW_1_io_dpath_status_xs),
    .io_dpath_status_fs(PTW_1_io_dpath_status_fs),
    .io_dpath_status_mpp(PTW_1_io_dpath_status_mpp),
    .io_dpath_status_hpp(PTW_1_io_dpath_status_hpp),
    .io_dpath_status_spp(PTW_1_io_dpath_status_spp),
    .io_dpath_status_mpie(PTW_1_io_dpath_status_mpie),
    .io_dpath_status_hpie(PTW_1_io_dpath_status_hpie),
    .io_dpath_status_spie(PTW_1_io_dpath_status_spie),
    .io_dpath_status_upie(PTW_1_io_dpath_status_upie),
    .io_dpath_status_mie(PTW_1_io_dpath_status_mie),
    .io_dpath_status_hie(PTW_1_io_dpath_status_hie),
    .io_dpath_status_sie(PTW_1_io_dpath_status_sie),
    .io_dpath_status_uie(PTW_1_io_dpath_status_uie)
  );
  HellaCacheArbiter dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_requestor_1_req_ready(dcArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_req_bits_phys(dcArb_io_requestor_1_req_bits_phys),
    .io_requestor_1_req_bits_data(dcArb_io_requestor_1_req_bits_data),
    .io_requestor_1_s1_kill(dcArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data(dcArb_io_requestor_1_s1_data),
    .io_requestor_1_s2_nack(dcArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_addr(dcArb_io_requestor_1_resp_bits_addr),
    .io_requestor_1_resp_bits_tag(dcArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_cmd(dcArb_io_requestor_1_resp_bits_cmd),
    .io_requestor_1_resp_bits_typ(dcArb_io_requestor_1_resp_bits_typ),
    .io_requestor_1_resp_bits_data(dcArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_resp_bits_store_data(dcArb_io_requestor_1_resp_bits_store_data),
    .io_requestor_1_replay_next(dcArb_io_requestor_1_replay_next),
    .io_requestor_1_xcpt_ma_ld(dcArb_io_requestor_1_xcpt_ma_ld),
    .io_requestor_1_xcpt_ma_st(dcArb_io_requestor_1_xcpt_ma_st),
    .io_requestor_1_xcpt_pf_ld(dcArb_io_requestor_1_xcpt_pf_ld),
    .io_requestor_1_xcpt_pf_st(dcArb_io_requestor_1_xcpt_pf_st),
    .io_requestor_1_invalidate_lr(dcArb_io_requestor_1_invalidate_lr),
    .io_requestor_1_ordered(dcArb_io_requestor_1_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = HellaCache_1_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = HellaCache_1_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = HellaCache_1_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = HellaCache_1_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = HellaCache_1_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = HellaCache_1_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = HellaCache_1_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = HellaCache_1_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = HellaCache_1_io_mem_probe_ready;
  assign io_cached_0_release_valid = HellaCache_1_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = HellaCache_1_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = HellaCache_1_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = HellaCache_1_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = HellaCache_1_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = HellaCache_1_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = HellaCache_1_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = HellaCache_1_io_mem_grant_ready;
  assign io_cached_0_finish_valid = HellaCache_1_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = HellaCache_1_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = HellaCache_1_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_btb_valid = icache_io_cpu_resp_bits_btb_valid;
  assign core_io_imem_resp_bits_btb_bits_taken = icache_io_cpu_resp_bits_btb_bits_taken;
  assign core_io_imem_resp_bits_btb_bits_mask = icache_io_cpu_resp_bits_btb_bits_mask;
  assign core_io_imem_resp_bits_btb_bits_bridx = icache_io_cpu_resp_bits_btb_bits_bridx;
  assign core_io_imem_resp_bits_btb_bits_target = icache_io_cpu_resp_bits_btb_bits_target;
  assign core_io_imem_resp_bits_btb_bits_entry = icache_io_cpu_resp_bits_btb_bits_entry;
  assign core_io_imem_resp_bits_btb_bits_bht_history = icache_io_cpu_resp_bits_btb_bits_bht_history;
  assign core_io_imem_resp_bits_btb_bits_bht_value = icache_io_cpu_resp_bits_btb_bits_bht_value;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data = icache_io_cpu_resp_bits_data;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_resp_bits_replay = icache_io_cpu_resp_bits_replay;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_1_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_1_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_1_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_1_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_1_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_1_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_1_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_1_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_1_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_1_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_1_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_1_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_1_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_1_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_1_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_1_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_1_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_1_ordered;
  assign core_io_fpu_fcsr_flags_valid = fpuOpt_io_fcsr_flags_valid;
  assign core_io_fpu_fcsr_flags_bits = fpuOpt_io_fcsr_flags_bits;
  assign core_io_fpu_store_data = fpuOpt_io_store_data;
  assign core_io_fpu_toint_data = fpuOpt_io_toint_data;
  assign core_io_fpu_fcsr_rdy = fpuOpt_io_fcsr_rdy;
  assign core_io_fpu_nack_mem = fpuOpt_io_nack_mem;
  assign core_io_fpu_illegal_rm = fpuOpt_io_illegal_rm;
  assign core_io_fpu_dec_cmd = fpuOpt_io_dec_cmd;
  assign core_io_fpu_dec_ldst = fpuOpt_io_dec_ldst;
  assign core_io_fpu_dec_wen = fpuOpt_io_dec_wen;
  assign core_io_fpu_dec_ren1 = fpuOpt_io_dec_ren1;
  assign core_io_fpu_dec_ren2 = fpuOpt_io_dec_ren2;
  assign core_io_fpu_dec_ren3 = fpuOpt_io_dec_ren3;
  assign core_io_fpu_dec_swap12 = fpuOpt_io_dec_swap12;
  assign core_io_fpu_dec_swap23 = fpuOpt_io_dec_swap23;
  assign core_io_fpu_dec_single = fpuOpt_io_dec_single;
  assign core_io_fpu_dec_fromint = fpuOpt_io_dec_fromint;
  assign core_io_fpu_dec_toint = fpuOpt_io_dec_toint;
  assign core_io_fpu_dec_fastpipe = fpuOpt_io_dec_fastpipe;
  assign core_io_fpu_dec_fma = fpuOpt_io_dec_fma;
  assign core_io_fpu_dec_div = fpuOpt_io_dec_div;
  assign core_io_fpu_dec_sqrt = fpuOpt_io_dec_sqrt;
  assign core_io_fpu_dec_round = fpuOpt_io_dec_round;
  assign core_io_fpu_dec_wflags = fpuOpt_io_dec_wflags;
  assign core_io_fpu_sboard_set = fpuOpt_io_sboard_set;
  assign core_io_fpu_sboard_clr = fpuOpt_io_sboard_clr;
  assign core_io_fpu_sboard_clra = fpuOpt_io_sboard_clra;
  assign core_io_fpu_cp_req_ready = fpuOpt_io_cp_req_ready;
  assign core_io_fpu_cp_resp_valid = fpuOpt_io_cp_resp_valid;
  assign core_io_fpu_cp_resp_bits_data = fpuOpt_io_cp_resp_bits_data;
  assign core_io_fpu_cp_resp_bits_exc = fpuOpt_io_cp_resp_bits_exc;
  assign core_io_rocc_cmd_ready = GEN_0;
  assign core_io_rocc_resp_valid = GEN_1;
  assign core_io_rocc_resp_bits_rd = GEN_2;
  assign core_io_rocc_resp_bits_data = GEN_3;
  assign core_io_rocc_mem_req_valid = GEN_4;
  assign core_io_rocc_mem_req_bits_addr = GEN_5;
  assign core_io_rocc_mem_req_bits_tag = GEN_6;
  assign core_io_rocc_mem_req_bits_cmd = GEN_7;
  assign core_io_rocc_mem_req_bits_typ = GEN_8;
  assign core_io_rocc_mem_req_bits_phys = GEN_9;
  assign core_io_rocc_mem_req_bits_data = GEN_10;
  assign core_io_rocc_mem_s1_kill = GEN_11;
  assign core_io_rocc_mem_s1_data = GEN_12;
  assign core_io_rocc_mem_invalidate_lr = GEN_13;
  assign core_io_rocc_busy = GEN_14;
  assign core_io_rocc_interrupt = GEN_15;
  assign core_io_rocc_autl_acquire_valid = GEN_16;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_17;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_18;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_19;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_20;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_21;
  assign core_io_rocc_autl_acquire_bits_union = GEN_22;
  assign core_io_rocc_autl_acquire_bits_data = GEN_23;
  assign core_io_rocc_autl_grant_ready = GEN_24;
  assign core_io_rocc_fpu_req_valid = GEN_25;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_26;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_27;
  assign core_io_rocc_fpu_req_bits_wen = GEN_28;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_29;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_30;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_31;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_32;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_33;
  assign core_io_rocc_fpu_req_bits_single = GEN_34;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_35;
  assign core_io_rocc_fpu_req_bits_toint = GEN_36;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_37;
  assign core_io_rocc_fpu_req_bits_fma = GEN_38;
  assign core_io_rocc_fpu_req_bits_div = GEN_39;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_40;
  assign core_io_rocc_fpu_req_bits_round = GEN_41;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_42;
  assign core_io_rocc_fpu_req_bits_rm = GEN_43;
  assign core_io_rocc_fpu_req_bits_typ = GEN_44;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_45;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_46;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_47;
  assign core_io_rocc_fpu_resp_ready = GEN_48;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = PTW_1_io_requestor_0_req_ready;
  assign icache_io_ptw_resp_valid = PTW_1_io_requestor_0_resp_valid;
  assign icache_io_ptw_resp_bits_pte_reserved_for_hardware = PTW_1_io_requestor_0_resp_bits_pte_reserved_for_hardware;
  assign icache_io_ptw_resp_bits_pte_ppn = PTW_1_io_requestor_0_resp_bits_pte_ppn;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = PTW_1_io_requestor_0_resp_bits_pte_reserved_for_software;
  assign icache_io_ptw_resp_bits_pte_d = PTW_1_io_requestor_0_resp_bits_pte_d;
  assign icache_io_ptw_resp_bits_pte_a = PTW_1_io_requestor_0_resp_bits_pte_a;
  assign icache_io_ptw_resp_bits_pte_g = PTW_1_io_requestor_0_resp_bits_pte_g;
  assign icache_io_ptw_resp_bits_pte_u = PTW_1_io_requestor_0_resp_bits_pte_u;
  assign icache_io_ptw_resp_bits_pte_x = PTW_1_io_requestor_0_resp_bits_pte_x;
  assign icache_io_ptw_resp_bits_pte_w = PTW_1_io_requestor_0_resp_bits_pte_w;
  assign icache_io_ptw_resp_bits_pte_r = PTW_1_io_requestor_0_resp_bits_pte_r;
  assign icache_io_ptw_resp_bits_pte_v = PTW_1_io_requestor_0_resp_bits_pte_v;
  assign icache_io_ptw_ptbr_asid = PTW_1_io_requestor_0_ptbr_asid;
  assign icache_io_ptw_ptbr_ppn = PTW_1_io_requestor_0_ptbr_ppn;
  assign icache_io_ptw_invalidate = PTW_1_io_requestor_0_invalidate;
  assign icache_io_ptw_status_debug = PTW_1_io_requestor_0_status_debug;
  assign icache_io_ptw_status_prv = PTW_1_io_requestor_0_status_prv;
  assign icache_io_ptw_status_sd = PTW_1_io_requestor_0_status_sd;
  assign icache_io_ptw_status_zero3 = PTW_1_io_requestor_0_status_zero3;
  assign icache_io_ptw_status_sd_rv32 = PTW_1_io_requestor_0_status_sd_rv32;
  assign icache_io_ptw_status_zero2 = PTW_1_io_requestor_0_status_zero2;
  assign icache_io_ptw_status_vm = PTW_1_io_requestor_0_status_vm;
  assign icache_io_ptw_status_zero1 = PTW_1_io_requestor_0_status_zero1;
  assign icache_io_ptw_status_mxr = PTW_1_io_requestor_0_status_mxr;
  assign icache_io_ptw_status_pum = PTW_1_io_requestor_0_status_pum;
  assign icache_io_ptw_status_mprv = PTW_1_io_requestor_0_status_mprv;
  assign icache_io_ptw_status_xs = PTW_1_io_requestor_0_status_xs;
  assign icache_io_ptw_status_fs = PTW_1_io_requestor_0_status_fs;
  assign icache_io_ptw_status_mpp = PTW_1_io_requestor_0_status_mpp;
  assign icache_io_ptw_status_hpp = PTW_1_io_requestor_0_status_hpp;
  assign icache_io_ptw_status_spp = PTW_1_io_requestor_0_status_spp;
  assign icache_io_ptw_status_mpie = PTW_1_io_requestor_0_status_mpie;
  assign icache_io_ptw_status_hpie = PTW_1_io_requestor_0_status_hpie;
  assign icache_io_ptw_status_spie = PTW_1_io_requestor_0_status_spie;
  assign icache_io_ptw_status_upie = PTW_1_io_requestor_0_status_upie;
  assign icache_io_ptw_status_mie = PTW_1_io_requestor_0_status_mie;
  assign icache_io_ptw_status_hie = PTW_1_io_requestor_0_status_hie;
  assign icache_io_ptw_status_sie = PTW_1_io_requestor_0_status_sie;
  assign icache_io_ptw_status_uie = PTW_1_io_requestor_0_status_uie;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign HellaCache_1_clk = clk;
  assign HellaCache_1_reset = reset;
  assign HellaCache_1_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign HellaCache_1_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign HellaCache_1_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign HellaCache_1_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign HellaCache_1_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign HellaCache_1_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign HellaCache_1_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign HellaCache_1_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign HellaCache_1_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign HellaCache_1_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign HellaCache_1_io_ptw_req_ready = PTW_1_io_requestor_1_req_ready;
  assign HellaCache_1_io_ptw_resp_valid = PTW_1_io_requestor_1_resp_valid;
  assign HellaCache_1_io_ptw_resp_bits_pte_reserved_for_hardware = PTW_1_io_requestor_1_resp_bits_pte_reserved_for_hardware;
  assign HellaCache_1_io_ptw_resp_bits_pte_ppn = PTW_1_io_requestor_1_resp_bits_pte_ppn;
  assign HellaCache_1_io_ptw_resp_bits_pte_reserved_for_software = PTW_1_io_requestor_1_resp_bits_pte_reserved_for_software;
  assign HellaCache_1_io_ptw_resp_bits_pte_d = PTW_1_io_requestor_1_resp_bits_pte_d;
  assign HellaCache_1_io_ptw_resp_bits_pte_a = PTW_1_io_requestor_1_resp_bits_pte_a;
  assign HellaCache_1_io_ptw_resp_bits_pte_g = PTW_1_io_requestor_1_resp_bits_pte_g;
  assign HellaCache_1_io_ptw_resp_bits_pte_u = PTW_1_io_requestor_1_resp_bits_pte_u;
  assign HellaCache_1_io_ptw_resp_bits_pte_x = PTW_1_io_requestor_1_resp_bits_pte_x;
  assign HellaCache_1_io_ptw_resp_bits_pte_w = PTW_1_io_requestor_1_resp_bits_pte_w;
  assign HellaCache_1_io_ptw_resp_bits_pte_r = PTW_1_io_requestor_1_resp_bits_pte_r;
  assign HellaCache_1_io_ptw_resp_bits_pte_v = PTW_1_io_requestor_1_resp_bits_pte_v;
  assign HellaCache_1_io_ptw_ptbr_asid = PTW_1_io_requestor_1_ptbr_asid;
  assign HellaCache_1_io_ptw_ptbr_ppn = PTW_1_io_requestor_1_ptbr_ppn;
  assign HellaCache_1_io_ptw_invalidate = PTW_1_io_requestor_1_invalidate;
  assign HellaCache_1_io_ptw_status_debug = PTW_1_io_requestor_1_status_debug;
  assign HellaCache_1_io_ptw_status_prv = PTW_1_io_requestor_1_status_prv;
  assign HellaCache_1_io_ptw_status_sd = PTW_1_io_requestor_1_status_sd;
  assign HellaCache_1_io_ptw_status_zero3 = PTW_1_io_requestor_1_status_zero3;
  assign HellaCache_1_io_ptw_status_sd_rv32 = PTW_1_io_requestor_1_status_sd_rv32;
  assign HellaCache_1_io_ptw_status_zero2 = PTW_1_io_requestor_1_status_zero2;
  assign HellaCache_1_io_ptw_status_vm = PTW_1_io_requestor_1_status_vm;
  assign HellaCache_1_io_ptw_status_zero1 = PTW_1_io_requestor_1_status_zero1;
  assign HellaCache_1_io_ptw_status_mxr = PTW_1_io_requestor_1_status_mxr;
  assign HellaCache_1_io_ptw_status_pum = PTW_1_io_requestor_1_status_pum;
  assign HellaCache_1_io_ptw_status_mprv = PTW_1_io_requestor_1_status_mprv;
  assign HellaCache_1_io_ptw_status_xs = PTW_1_io_requestor_1_status_xs;
  assign HellaCache_1_io_ptw_status_fs = PTW_1_io_requestor_1_status_fs;
  assign HellaCache_1_io_ptw_status_mpp = PTW_1_io_requestor_1_status_mpp;
  assign HellaCache_1_io_ptw_status_hpp = PTW_1_io_requestor_1_status_hpp;
  assign HellaCache_1_io_ptw_status_spp = PTW_1_io_requestor_1_status_spp;
  assign HellaCache_1_io_ptw_status_mpie = PTW_1_io_requestor_1_status_mpie;
  assign HellaCache_1_io_ptw_status_hpie = PTW_1_io_requestor_1_status_hpie;
  assign HellaCache_1_io_ptw_status_spie = PTW_1_io_requestor_1_status_spie;
  assign HellaCache_1_io_ptw_status_upie = PTW_1_io_requestor_1_status_upie;
  assign HellaCache_1_io_ptw_status_mie = PTW_1_io_requestor_1_status_mie;
  assign HellaCache_1_io_ptw_status_hie = PTW_1_io_requestor_1_status_hie;
  assign HellaCache_1_io_ptw_status_sie = PTW_1_io_requestor_1_status_sie;
  assign HellaCache_1_io_ptw_status_uie = PTW_1_io_requestor_1_status_uie;
  assign HellaCache_1_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign HellaCache_1_io_mem_probe_valid = io_cached_0_probe_valid;
  assign HellaCache_1_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign HellaCache_1_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign HellaCache_1_io_mem_release_ready = io_cached_0_release_ready;
  assign HellaCache_1_io_mem_grant_valid = io_cached_0_grant_valid;
  assign HellaCache_1_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign HellaCache_1_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign HellaCache_1_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign HellaCache_1_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign HellaCache_1_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign HellaCache_1_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign HellaCache_1_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign HellaCache_1_io_mem_finish_ready = io_cached_0_finish_ready;
  assign fpuOpt_clk = clk;
  assign fpuOpt_reset = reset;
  assign fpuOpt_io_inst = core_io_fpu_inst;
  assign fpuOpt_io_fromint_data = core_io_fpu_fromint_data;
  assign fpuOpt_io_fcsr_rm = core_io_fpu_fcsr_rm;
  assign fpuOpt_io_dmem_resp_val = core_io_fpu_dmem_resp_val;
  assign fpuOpt_io_dmem_resp_type = core_io_fpu_dmem_resp_type;
  assign fpuOpt_io_dmem_resp_tag = core_io_fpu_dmem_resp_tag;
  assign fpuOpt_io_dmem_resp_data = core_io_fpu_dmem_resp_data;
  assign fpuOpt_io_valid = core_io_fpu_valid;
  assign fpuOpt_io_killx = core_io_fpu_killx;
  assign fpuOpt_io_killm = core_io_fpu_killm;
  assign fpuOpt_io_cp_req_valid = 1'h0;
  assign fpuOpt_io_cp_req_bits_cmd = core_io_fpu_cp_req_bits_cmd;
  assign fpuOpt_io_cp_req_bits_ldst = core_io_fpu_cp_req_bits_ldst;
  assign fpuOpt_io_cp_req_bits_wen = core_io_fpu_cp_req_bits_wen;
  assign fpuOpt_io_cp_req_bits_ren1 = core_io_fpu_cp_req_bits_ren1;
  assign fpuOpt_io_cp_req_bits_ren2 = core_io_fpu_cp_req_bits_ren2;
  assign fpuOpt_io_cp_req_bits_ren3 = core_io_fpu_cp_req_bits_ren3;
  assign fpuOpt_io_cp_req_bits_swap12 = core_io_fpu_cp_req_bits_swap12;
  assign fpuOpt_io_cp_req_bits_swap23 = core_io_fpu_cp_req_bits_swap23;
  assign fpuOpt_io_cp_req_bits_single = core_io_fpu_cp_req_bits_single;
  assign fpuOpt_io_cp_req_bits_fromint = core_io_fpu_cp_req_bits_fromint;
  assign fpuOpt_io_cp_req_bits_toint = core_io_fpu_cp_req_bits_toint;
  assign fpuOpt_io_cp_req_bits_fastpipe = core_io_fpu_cp_req_bits_fastpipe;
  assign fpuOpt_io_cp_req_bits_fma = core_io_fpu_cp_req_bits_fma;
  assign fpuOpt_io_cp_req_bits_div = core_io_fpu_cp_req_bits_div;
  assign fpuOpt_io_cp_req_bits_sqrt = core_io_fpu_cp_req_bits_sqrt;
  assign fpuOpt_io_cp_req_bits_round = core_io_fpu_cp_req_bits_round;
  assign fpuOpt_io_cp_req_bits_wflags = core_io_fpu_cp_req_bits_wflags;
  assign fpuOpt_io_cp_req_bits_rm = core_io_fpu_cp_req_bits_rm;
  assign fpuOpt_io_cp_req_bits_typ = core_io_fpu_cp_req_bits_typ;
  assign fpuOpt_io_cp_req_bits_in1 = core_io_fpu_cp_req_bits_in1;
  assign fpuOpt_io_cp_req_bits_in2 = core_io_fpu_cp_req_bits_in2;
  assign fpuOpt_io_cp_req_bits_in3 = core_io_fpu_cp_req_bits_in3;
  assign fpuOpt_io_cp_resp_ready = 1'h0;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign PTW_1_clk = clk;
  assign PTW_1_reset = reset;
  assign PTW_1_io_requestor_0_req_valid = icache_io_ptw_req_valid;
  assign PTW_1_io_requestor_0_req_bits_prv = icache_io_ptw_req_bits_prv;
  assign PTW_1_io_requestor_0_req_bits_pum = icache_io_ptw_req_bits_pum;
  assign PTW_1_io_requestor_0_req_bits_mxr = icache_io_ptw_req_bits_mxr;
  assign PTW_1_io_requestor_0_req_bits_addr = icache_io_ptw_req_bits_addr;
  assign PTW_1_io_requestor_0_req_bits_store = icache_io_ptw_req_bits_store;
  assign PTW_1_io_requestor_0_req_bits_fetch = icache_io_ptw_req_bits_fetch;
  assign PTW_1_io_requestor_1_req_valid = HellaCache_1_io_ptw_req_valid;
  assign PTW_1_io_requestor_1_req_bits_prv = HellaCache_1_io_ptw_req_bits_prv;
  assign PTW_1_io_requestor_1_req_bits_pum = HellaCache_1_io_ptw_req_bits_pum;
  assign PTW_1_io_requestor_1_req_bits_mxr = HellaCache_1_io_ptw_req_bits_mxr;
  assign PTW_1_io_requestor_1_req_bits_addr = HellaCache_1_io_ptw_req_bits_addr;
  assign PTW_1_io_requestor_1_req_bits_store = HellaCache_1_io_ptw_req_bits_store;
  assign PTW_1_io_requestor_1_req_bits_fetch = HellaCache_1_io_ptw_req_bits_fetch;
  assign PTW_1_io_mem_req_ready = dcArb_io_requestor_0_req_ready;
  assign PTW_1_io_mem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign PTW_1_io_mem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign PTW_1_io_mem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign PTW_1_io_mem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign PTW_1_io_mem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign PTW_1_io_mem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign PTW_1_io_mem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign PTW_1_io_mem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign PTW_1_io_mem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign PTW_1_io_mem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign PTW_1_io_mem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign PTW_1_io_mem_replay_next = dcArb_io_requestor_0_replay_next;
  assign PTW_1_io_mem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign PTW_1_io_mem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign PTW_1_io_mem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign PTW_1_io_mem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign PTW_1_io_mem_ordered = dcArb_io_requestor_0_ordered;
  assign PTW_1_io_dpath_ptbr_asid = core_io_ptw_ptbr_asid;
  assign PTW_1_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn;
  assign PTW_1_io_dpath_invalidate = core_io_ptw_invalidate;
  assign PTW_1_io_dpath_status_debug = core_io_ptw_status_debug;
  assign PTW_1_io_dpath_status_prv = core_io_ptw_status_prv;
  assign PTW_1_io_dpath_status_sd = core_io_ptw_status_sd;
  assign PTW_1_io_dpath_status_zero3 = core_io_ptw_status_zero3;
  assign PTW_1_io_dpath_status_sd_rv32 = core_io_ptw_status_sd_rv32;
  assign PTW_1_io_dpath_status_zero2 = core_io_ptw_status_zero2;
  assign PTW_1_io_dpath_status_vm = core_io_ptw_status_vm;
  assign PTW_1_io_dpath_status_zero1 = core_io_ptw_status_zero1;
  assign PTW_1_io_dpath_status_mxr = core_io_ptw_status_mxr;
  assign PTW_1_io_dpath_status_pum = core_io_ptw_status_pum;
  assign PTW_1_io_dpath_status_mprv = core_io_ptw_status_mprv;
  assign PTW_1_io_dpath_status_xs = core_io_ptw_status_xs;
  assign PTW_1_io_dpath_status_fs = core_io_ptw_status_fs;
  assign PTW_1_io_dpath_status_mpp = core_io_ptw_status_mpp;
  assign PTW_1_io_dpath_status_hpp = core_io_ptw_status_hpp;
  assign PTW_1_io_dpath_status_spp = core_io_ptw_status_spp;
  assign PTW_1_io_dpath_status_mpie = core_io_ptw_status_mpie;
  assign PTW_1_io_dpath_status_hpie = core_io_ptw_status_hpie;
  assign PTW_1_io_dpath_status_spie = core_io_ptw_status_spie;
  assign PTW_1_io_dpath_status_upie = core_io_ptw_status_upie;
  assign PTW_1_io_dpath_status_mie = core_io_ptw_status_mie;
  assign PTW_1_io_dpath_status_hie = core_io_ptw_status_hie;
  assign PTW_1_io_dpath_status_sie = core_io_ptw_status_sie;
  assign PTW_1_io_dpath_status_uie = core_io_ptw_status_uie;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = PTW_1_io_mem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = PTW_1_io_mem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = PTW_1_io_mem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = PTW_1_io_mem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = PTW_1_io_mem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = PTW_1_io_mem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = PTW_1_io_mem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = PTW_1_io_mem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = PTW_1_io_mem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = PTW_1_io_mem_invalidate_lr;
  assign dcArb_io_requestor_1_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_1_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_1_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_1_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_1_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = HellaCache_1_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = HellaCache_1_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = HellaCache_1_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = HellaCache_1_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = HellaCache_1_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = HellaCache_1_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = HellaCache_1_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = HellaCache_1_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = HellaCache_1_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = HellaCache_1_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = HellaCache_1_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = HellaCache_1_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = HellaCache_1_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = HellaCache_1_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = HellaCache_1_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = HellaCache_1_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = HellaCache_1_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = HellaCache_1_io_cpu_ordered;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_51[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_52[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_53[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_54[39:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_55[6:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_56[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_57[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_58[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_59[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_60[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_12 = GEN_61[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_62[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_63[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_64[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_65[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_66[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_18 = GEN_67[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_19 = GEN_68[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_20 = GEN_69[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_21 = GEN_70[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_22 = GEN_71[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_23 = GEN_72[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_24 = GEN_73[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_25 = GEN_74[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_26 = GEN_75[4:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_27 = GEN_76[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_28 = GEN_77[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_78[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_79[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_32 = GEN_81[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_33 = GEN_82[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_83[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_84[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_87[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_39 = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_89[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_41 = GEN_90[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_42 = GEN_91[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_43 = GEN_92[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_44 = GEN_93[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_45 = GEN_94[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_46 = GEN_95[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_47 = GEN_96[64:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_48 = GEN_97[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_49 = {1{$random}};
  GEN_50 = {1{$random}};
  GEN_51 = {1{$random}};
  GEN_52 = {2{$random}};
  GEN_53 = {1{$random}};
  GEN_54 = {2{$random}};
  GEN_55 = {1{$random}};
  GEN_56 = {1{$random}};
  GEN_57 = {1{$random}};
  GEN_58 = {1{$random}};
  GEN_59 = {2{$random}};
  GEN_60 = {1{$random}};
  GEN_61 = {2{$random}};
  GEN_62 = {1{$random}};
  GEN_63 = {1{$random}};
  GEN_64 = {1{$random}};
  GEN_65 = {1{$random}};
  GEN_66 = {1{$random}};
  GEN_67 = {1{$random}};
  GEN_68 = {1{$random}};
  GEN_69 = {1{$random}};
  GEN_70 = {1{$random}};
  GEN_71 = {1{$random}};
  GEN_72 = {2{$random}};
  GEN_73 = {1{$random}};
  GEN_74 = {1{$random}};
  GEN_75 = {1{$random}};
  GEN_76 = {1{$random}};
  GEN_77 = {1{$random}};
  GEN_78 = {1{$random}};
  GEN_79 = {1{$random}};
  GEN_80 = {1{$random}};
  GEN_81 = {1{$random}};
  GEN_82 = {1{$random}};
  GEN_83 = {1{$random}};
  GEN_84 = {1{$random}};
  GEN_85 = {1{$random}};
  GEN_86 = {1{$random}};
  GEN_87 = {1{$random}};
  GEN_88 = {1{$random}};
  GEN_89 = {1{$random}};
  GEN_90 = {1{$random}};
  GEN_91 = {1{$random}};
  GEN_92 = {1{$random}};
  GEN_93 = {1{$random}};
  GEN_94 = {3{$random}};
  GEN_95 = {3{$random}};
  GEN_96 = {3{$random}};
  GEN_97 = {1{$random}};
  end
`endif
endmodule
module Queue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_is_builtin_type,
  input  [2:0] io_enq_bits_payload_a_type,
  input  [10:0] io_enq_bits_payload_union,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_is_builtin_type,
  output [2:0] io_deq_bits_payload_a_type,
  output [10:0] io_deq_bits_payload_union,
  output [63:0] io_deq_bits_payload_data,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1025_data;
  wire  ram_header_src_T_1025_addr;
  wire  ram_header_src_T_1025_mask;
  wire  ram_header_src_T_1025_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1025_data;
  wire  ram_header_dst_T_1025_addr;
  wire  ram_header_dst_T_1025_mask;
  wire  ram_header_dst_T_1025_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1025_data;
  wire  ram_payload_addr_block_T_1025_addr;
  wire  ram_payload_addr_block_T_1025_mask;
  wire  ram_payload_addr_block_T_1025_en;
  reg [1:0] ram_payload_client_xact_id [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire [1:0] ram_payload_client_xact_id_T_1025_data;
  wire  ram_payload_client_xact_id_T_1025_addr;
  wire  ram_payload_client_xact_id_T_1025_mask;
  wire  ram_payload_client_xact_id_T_1025_en;
  reg [2:0] ram_payload_addr_beat [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1025_data;
  wire  ram_payload_addr_beat_T_1025_addr;
  wire  ram_payload_addr_beat_T_1025_mask;
  wire  ram_payload_addr_beat_T_1025_en;
  reg  ram_payload_is_builtin_type [0:0];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1025_data;
  wire  ram_payload_is_builtin_type_T_1025_addr;
  wire  ram_payload_is_builtin_type_T_1025_mask;
  wire  ram_payload_is_builtin_type_T_1025_en;
  reg [2:0] ram_payload_a_type [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_a_type_T_1144_data;
  wire  ram_payload_a_type_T_1144_addr;
  wire  ram_payload_a_type_T_1144_en;
  wire [2:0] ram_payload_a_type_T_1025_data;
  wire  ram_payload_a_type_T_1025_addr;
  wire  ram_payload_a_type_T_1025_mask;
  wire  ram_payload_a_type_T_1025_en;
  reg [10:0] ram_payload_union [0:0];
  reg [31:0] GEN_7;
  wire [10:0] ram_payload_union_T_1144_data;
  wire  ram_payload_union_T_1144_addr;
  wire  ram_payload_union_T_1144_en;
  wire [10:0] ram_payload_union_T_1025_data;
  wire  ram_payload_union_T_1025_addr;
  wire  ram_payload_union_T_1025_mask;
  wire  ram_payload_union_T_1025_en;
  reg [63:0] ram_payload_data [0:0];
  reg [63:0] GEN_8;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1025_data;
  wire  ram_payload_data_T_1025_addr;
  wire  ram_payload_data_T_1025_mask;
  wire  ram_payload_data_T_1025_en;
  reg  maybe_full;
  reg [31:0] GEN_9;
  wire  T_1022;
  wire  T_1023;
  wire  do_enq;
  wire  T_1024;
  wire  do_deq;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire [1:0] T_1256;
  wire  ptr_diff;
  wire [1:0] T_1258;
  assign io_enq_ready = T_1022;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_a_type = ram_payload_a_type_T_1144_data;
  assign io_deq_bits_payload_union = ram_payload_union_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1258[0];
  assign ram_header_src_T_1144_addr = 1'h0;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1025_data = io_enq_bits_header_src;
  assign ram_header_src_T_1025_addr = 1'h0;
  assign ram_header_src_T_1025_mask = do_enq;
  assign ram_header_src_T_1025_en = do_enq;
  assign ram_header_dst_T_1144_addr = 1'h0;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1025_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1025_addr = 1'h0;
  assign ram_header_dst_T_1025_mask = do_enq;
  assign ram_header_dst_T_1025_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = 1'h0;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1025_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1025_addr = 1'h0;
  assign ram_payload_addr_block_T_1025_mask = do_enq;
  assign ram_payload_addr_block_T_1025_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1025_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1025_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1025_mask = do_enq;
  assign ram_payload_client_xact_id_T_1025_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = 1'h0;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1025_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1025_addr = 1'h0;
  assign ram_payload_addr_beat_T_1025_mask = do_enq;
  assign ram_payload_addr_beat_T_1025_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1025_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1025_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1025_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1025_en = do_enq;
  assign ram_payload_a_type_T_1144_addr = 1'h0;
  assign ram_payload_a_type_T_1144_en = 1'h1;
  assign ram_payload_a_type_T_1144_data = ram_payload_a_type[ram_payload_a_type_T_1144_addr];
  assign ram_payload_a_type_T_1025_data = io_enq_bits_payload_a_type;
  assign ram_payload_a_type_T_1025_addr = 1'h0;
  assign ram_payload_a_type_T_1025_mask = do_enq;
  assign ram_payload_a_type_T_1025_en = do_enq;
  assign ram_payload_union_T_1144_addr = 1'h0;
  assign ram_payload_union_T_1144_en = 1'h1;
  assign ram_payload_union_T_1144_data = ram_payload_union[ram_payload_union_T_1144_addr];
  assign ram_payload_union_T_1025_data = io_enq_bits_payload_union;
  assign ram_payload_union_T_1025_addr = 1'h0;
  assign ram_payload_union_T_1025_mask = do_enq;
  assign ram_payload_union_T_1025_en = do_enq;
  assign ram_payload_data_T_1144_addr = 1'h0;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1025_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1025_addr = 1'h0;
  assign ram_payload_data_T_1025_mask = do_enq;
  assign ram_payload_data_T_1025_en = do_enq;
  assign T_1022 = maybe_full == 1'h0;
  assign T_1023 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1023;
  assign T_1024 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1024;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = T_1022 == 1'h0;
  assign T_1256 = 1'h0 - 1'h0;
  assign ptr_diff = T_1256[0:0];
  assign T_1258 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_a_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_union[initvar] = GEN_7[10:0];
  `endif
  GEN_8 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_8[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  maybe_full = GEN_9[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1025_en & ram_header_src_T_1025_mask) begin
      ram_header_src[ram_header_src_T_1025_addr] <= ram_header_src_T_1025_data;
    end
    if(ram_header_dst_T_1025_en & ram_header_dst_T_1025_mask) begin
      ram_header_dst[ram_header_dst_T_1025_addr] <= ram_header_dst_T_1025_data;
    end
    if(ram_payload_addr_block_T_1025_en & ram_payload_addr_block_T_1025_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1025_addr] <= ram_payload_addr_block_T_1025_data;
    end
    if(ram_payload_client_xact_id_T_1025_en & ram_payload_client_xact_id_T_1025_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1025_addr] <= ram_payload_client_xact_id_T_1025_data;
    end
    if(ram_payload_addr_beat_T_1025_en & ram_payload_addr_beat_T_1025_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1025_addr] <= ram_payload_addr_beat_T_1025_data;
    end
    if(ram_payload_is_builtin_type_T_1025_en & ram_payload_is_builtin_type_T_1025_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1025_addr] <= ram_payload_is_builtin_type_T_1025_data;
    end
    if(ram_payload_a_type_T_1025_en & ram_payload_a_type_T_1025_mask) begin
      ram_payload_a_type[ram_payload_a_type_T_1025_addr] <= ram_payload_a_type_T_1025_data;
    end
    if(ram_payload_union_T_1025_en & ram_payload_union_T_1025_mask) begin
      ram_payload_union[ram_payload_union_T_1025_addr] <= ram_payload_union_T_1025_data;
    end
    if(ram_payload_data_T_1025_en & ram_payload_data_T_1025_mask) begin
      ram_payload_data[ram_payload_data_T_1025_addr] <= ram_payload_data_T_1025_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_p_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_p_type,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1094_data;
  wire  ram_header_src_T_1094_addr;
  wire  ram_header_src_T_1094_en;
  wire [1:0] ram_header_src_T_980_data;
  wire  ram_header_src_T_980_addr;
  wire  ram_header_src_T_980_mask;
  wire  ram_header_src_T_980_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1094_data;
  wire  ram_header_dst_T_1094_addr;
  wire  ram_header_dst_T_1094_en;
  wire [1:0] ram_header_dst_T_980_data;
  wire  ram_header_dst_T_980_addr;
  wire  ram_header_dst_T_980_mask;
  wire  ram_header_dst_T_980_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1094_data;
  wire  ram_payload_addr_block_T_1094_addr;
  wire  ram_payload_addr_block_T_1094_en;
  wire [25:0] ram_payload_addr_block_T_980_data;
  wire  ram_payload_addr_block_T_980_addr;
  wire  ram_payload_addr_block_T_980_mask;
  wire  ram_payload_addr_block_T_980_en;
  reg [1:0] ram_payload_p_type [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_p_type_T_1094_data;
  wire  ram_payload_p_type_T_1094_addr;
  wire  ram_payload_p_type_T_1094_en;
  wire [1:0] ram_payload_p_type_T_980_data;
  wire  ram_payload_p_type_T_980_addr;
  wire  ram_payload_p_type_T_980_mask;
  wire  ram_payload_p_type_T_980_en;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  T_977;
  wire  T_978;
  wire  do_enq;
  wire  T_979;
  wire  do_deq;
  wire  T_1089;
  wire  GEN_11;
  wire  T_1091;
  wire [1:0] T_1201;
  wire  ptr_diff;
  wire [1:0] T_1203;
  assign io_enq_ready = T_977;
  assign io_deq_valid = T_1091;
  assign io_deq_bits_header_src = ram_header_src_T_1094_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1094_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1094_data;
  assign io_deq_bits_payload_p_type = ram_payload_p_type_T_1094_data;
  assign io_count = T_1203[0];
  assign ram_header_src_T_1094_addr = 1'h0;
  assign ram_header_src_T_1094_en = 1'h1;
  assign ram_header_src_T_1094_data = ram_header_src[ram_header_src_T_1094_addr];
  assign ram_header_src_T_980_data = io_enq_bits_header_src;
  assign ram_header_src_T_980_addr = 1'h0;
  assign ram_header_src_T_980_mask = do_enq;
  assign ram_header_src_T_980_en = do_enq;
  assign ram_header_dst_T_1094_addr = 1'h0;
  assign ram_header_dst_T_1094_en = 1'h1;
  assign ram_header_dst_T_1094_data = ram_header_dst[ram_header_dst_T_1094_addr];
  assign ram_header_dst_T_980_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_980_addr = 1'h0;
  assign ram_header_dst_T_980_mask = do_enq;
  assign ram_header_dst_T_980_en = do_enq;
  assign ram_payload_addr_block_T_1094_addr = 1'h0;
  assign ram_payload_addr_block_T_1094_en = 1'h1;
  assign ram_payload_addr_block_T_1094_data = ram_payload_addr_block[ram_payload_addr_block_T_1094_addr];
  assign ram_payload_addr_block_T_980_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_980_addr = 1'h0;
  assign ram_payload_addr_block_T_980_mask = do_enq;
  assign ram_payload_addr_block_T_980_en = do_enq;
  assign ram_payload_p_type_T_1094_addr = 1'h0;
  assign ram_payload_p_type_T_1094_en = 1'h1;
  assign ram_payload_p_type_T_1094_data = ram_payload_p_type[ram_payload_p_type_T_1094_addr];
  assign ram_payload_p_type_T_980_data = io_enq_bits_payload_p_type;
  assign ram_payload_p_type_T_980_addr = 1'h0;
  assign ram_payload_p_type_T_980_mask = do_enq;
  assign ram_payload_p_type_T_980_en = do_enq;
  assign T_977 = maybe_full == 1'h0;
  assign T_978 = io_enq_ready & io_enq_valid;
  assign do_enq = T_978;
  assign T_979 = io_deq_ready & io_deq_valid;
  assign do_deq = T_979;
  assign T_1089 = do_enq != do_deq;
  assign GEN_11 = T_1089 ? do_enq : maybe_full;
  assign T_1091 = T_977 == 1'h0;
  assign T_1201 = 1'h0 - 1'h0;
  assign ptr_diff = T_1201[0:0];
  assign T_1203 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_p_type[initvar] = GEN_3[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_980_en & ram_header_src_T_980_mask) begin
      ram_header_src[ram_header_src_T_980_addr] <= ram_header_src_T_980_data;
    end
    if(ram_header_dst_T_980_en & ram_header_dst_T_980_mask) begin
      ram_header_dst[ram_header_dst_T_980_addr] <= ram_header_dst_T_980_data;
    end
    if(ram_payload_addr_block_T_980_en & ram_payload_addr_block_T_980_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_980_addr] <= ram_payload_addr_block_T_980_data;
    end
    if(ram_payload_p_type_T_980_en & ram_payload_p_type_T_980_mask) begin
      ram_payload_p_type[ram_payload_p_type_T_980_addr] <= ram_payload_p_type_T_980_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1089) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_4(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input   io_enq_bits_payload_voluntary,
  input  [2:0] io_enq_bits_payload_r_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output  io_deq_bits_payload_voluntary,
  output [2:0] io_deq_bits_payload_r_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg [25:0] ram_payload_addr_block [0:1];
  reg [31:0] GEN_3;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1018_data;
  wire  ram_payload_addr_block_T_1018_addr;
  wire  ram_payload_addr_block_T_1018_mask;
  wire  ram_payload_addr_block_T_1018_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [1:0] ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire [1:0] ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg  ram_payload_voluntary [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_voluntary_T_1144_data;
  wire  ram_payload_voluntary_T_1144_addr;
  wire  ram_payload_voluntary_T_1144_en;
  wire  ram_payload_voluntary_T_1018_data;
  wire  ram_payload_voluntary_T_1018_addr;
  wire  ram_payload_voluntary_T_1018_mask;
  wire  ram_payload_voluntary_T_1018_en;
  reg [2:0] ram_payload_r_type [0:1];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_r_type_T_1144_data;
  wire  ram_payload_r_type_T_1144_addr;
  wire  ram_payload_r_type_T_1144_en;
  wire [2:0] ram_payload_r_type_T_1018_data;
  wire  ram_payload_r_type_T_1018_addr;
  wire  ram_payload_r_type_T_1018_mask;
  wire  ram_payload_r_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_voluntary = ram_payload_voluntary_T_1144_data;
  assign io_deq_bits_payload_r_type = ram_payload_r_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = T_1012;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1018_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1018_addr = T_1010;
  assign ram_payload_addr_block_T_1018_mask = do_enq;
  assign ram_payload_addr_block_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_voluntary_T_1144_addr = T_1012;
  assign ram_payload_voluntary_T_1144_en = 1'h1;
  assign ram_payload_voluntary_T_1144_data = ram_payload_voluntary[ram_payload_voluntary_T_1144_addr];
  assign ram_payload_voluntary_T_1018_data = io_enq_bits_payload_voluntary;
  assign ram_payload_voluntary_T_1018_addr = T_1010;
  assign ram_payload_voluntary_T_1018_mask = do_enq;
  assign ram_payload_voluntary_T_1018_en = do_enq;
  assign ram_payload_r_type_T_1144_addr = T_1012;
  assign ram_payload_r_type_T_1144_en = 1'h1;
  assign ram_payload_r_type_T_1144_data = ram_payload_r_type[ram_payload_r_type_T_1144_addr];
  assign ram_payload_r_type_T_1018_data = io_enq_bits_payload_r_type;
  assign ram_payload_r_type_T_1018_addr = T_1010;
  assign ram_payload_r_type_T_1018_mask = do_enq;
  assign ram_payload_r_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_3[25:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_4[1:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_voluntary[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_r_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_addr_block_T_1018_en & ram_payload_addr_block_T_1018_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1018_addr] <= ram_payload_addr_block_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_voluntary_T_1018_en & ram_payload_voluntary_T_1018_mask) begin
      ram_payload_voluntary[ram_payload_voluntary_T_1018_addr] <= ram_payload_voluntary_T_1018_data;
    end
    if(ram_payload_r_type_T_1018_en & ram_payload_r_type_T_1018_mask) begin
      ram_payload_r_type[ram_payload_r_type_T_1018_addr] <= ram_payload_r_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_5(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_manager_xact_id,
  input   io_enq_bits_payload_is_builtin_type,
  input  [3:0] io_enq_bits_payload_g_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_manager_xact_id,
  output  io_deq_bits_payload_is_builtin_type,
  output [3:0] io_deq_bits_payload_g_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire [1:0] ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg [2:0] ram_payload_manager_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_manager_xact_id_T_1144_data;
  wire  ram_payload_manager_xact_id_T_1144_addr;
  wire  ram_payload_manager_xact_id_T_1144_en;
  wire [2:0] ram_payload_manager_xact_id_T_1018_data;
  wire  ram_payload_manager_xact_id_T_1018_addr;
  wire  ram_payload_manager_xact_id_T_1018_mask;
  wire  ram_payload_manager_xact_id_T_1018_en;
  reg  ram_payload_is_builtin_type [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1018_data;
  wire  ram_payload_is_builtin_type_T_1018_addr;
  wire  ram_payload_is_builtin_type_T_1018_mask;
  wire  ram_payload_is_builtin_type_T_1018_en;
  reg [3:0] ram_payload_g_type [0:1];
  reg [31:0] GEN_6;
  wire [3:0] ram_payload_g_type_T_1144_data;
  wire  ram_payload_g_type_T_1144_addr;
  wire  ram_payload_g_type_T_1144_en;
  wire [3:0] ram_payload_g_type_T_1018_data;
  wire  ram_payload_g_type_T_1018_addr;
  wire  ram_payload_g_type_T_1018_mask;
  wire  ram_payload_g_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_manager_xact_id = ram_payload_manager_xact_id_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_g_type = ram_payload_g_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_manager_xact_id_T_1144_addr = T_1012;
  assign ram_payload_manager_xact_id_T_1144_en = 1'h1;
  assign ram_payload_manager_xact_id_T_1144_data = ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1144_addr];
  assign ram_payload_manager_xact_id_T_1018_data = io_enq_bits_payload_manager_xact_id;
  assign ram_payload_manager_xact_id_T_1018_addr = T_1010;
  assign ram_payload_manager_xact_id_T_1018_mask = do_enq;
  assign ram_payload_manager_xact_id_T_1018_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = T_1012;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1018_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1018_addr = T_1010;
  assign ram_payload_is_builtin_type_T_1018_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1018_en = do_enq;
  assign ram_payload_g_type_T_1144_addr = T_1012;
  assign ram_payload_g_type_T_1144_en = 1'h1;
  assign ram_payload_g_type_T_1144_data = ram_payload_g_type[ram_payload_g_type_T_1144_addr];
  assign ram_payload_g_type_T_1018_data = io_enq_bits_payload_g_type;
  assign ram_payload_g_type_T_1018_addr = T_1010;
  assign ram_payload_g_type_T_1018_mask = do_enq;
  assign ram_payload_g_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_manager_xact_id[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_g_type[initvar] = GEN_6[3:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_manager_xact_id_T_1018_en & ram_payload_manager_xact_id_T_1018_mask) begin
      ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1018_addr] <= ram_payload_manager_xact_id_T_1018_data;
    end
    if(ram_payload_is_builtin_type_T_1018_en & ram_payload_is_builtin_type_T_1018_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1018_addr] <= ram_payload_is_builtin_type_T_1018_data;
    end
    if(ram_payload_g_type_T_1018_en & ram_payload_g_type_T_1018_mask) begin
      ram_payload_g_type[ram_payload_g_type_T_1018_addr] <= ram_payload_g_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_2_1_clk;
  wire  Queue_2_1_reset;
  wire  Queue_2_1_io_enq_ready;
  wire  Queue_2_1_io_enq_valid;
  wire [1:0] Queue_2_1_io_enq_bits_header_src;
  wire [1:0] Queue_2_1_io_enq_bits_header_dst;
  wire [25:0] Queue_2_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_2_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_2_1_io_enq_bits_payload_addr_beat;
  wire  Queue_2_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_2_1_io_enq_bits_payload_a_type;
  wire [10:0] Queue_2_1_io_enq_bits_payload_union;
  wire [63:0] Queue_2_1_io_enq_bits_payload_data;
  wire  Queue_2_1_io_deq_ready;
  wire  Queue_2_1_io_deq_valid;
  wire [1:0] Queue_2_1_io_deq_bits_header_src;
  wire [1:0] Queue_2_1_io_deq_bits_header_dst;
  wire [25:0] Queue_2_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_2_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_2_1_io_deq_bits_payload_addr_beat;
  wire  Queue_2_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_2_1_io_deq_bits_payload_a_type;
  wire [10:0] Queue_2_1_io_deq_bits_payload_union;
  wire [63:0] Queue_2_1_io_deq_bits_payload_data;
  wire  Queue_2_1_io_count;
  wire  Queue_3_1_clk;
  wire  Queue_3_1_reset;
  wire  Queue_3_1_io_enq_ready;
  wire  Queue_3_1_io_enq_valid;
  wire [1:0] Queue_3_1_io_enq_bits_header_src;
  wire [1:0] Queue_3_1_io_enq_bits_header_dst;
  wire [25:0] Queue_3_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_3_1_io_enq_bits_payload_p_type;
  wire  Queue_3_1_io_deq_ready;
  wire  Queue_3_1_io_deq_valid;
  wire [1:0] Queue_3_1_io_deq_bits_header_src;
  wire [1:0] Queue_3_1_io_deq_bits_header_dst;
  wire [25:0] Queue_3_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_3_1_io_deq_bits_payload_p_type;
  wire  Queue_3_1_io_count;
  wire  Queue_4_1_clk;
  wire  Queue_4_1_reset;
  wire  Queue_4_1_io_enq_ready;
  wire  Queue_4_1_io_enq_valid;
  wire [1:0] Queue_4_1_io_enq_bits_header_src;
  wire [1:0] Queue_4_1_io_enq_bits_header_dst;
  wire [2:0] Queue_4_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_4_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_4_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_4_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_4_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_4_1_io_enq_bits_payload_data;
  wire  Queue_4_1_io_deq_ready;
  wire  Queue_4_1_io_deq_valid;
  wire [1:0] Queue_4_1_io_deq_bits_header_src;
  wire [1:0] Queue_4_1_io_deq_bits_header_dst;
  wire [2:0] Queue_4_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_4_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_4_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_4_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_4_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_4_1_io_deq_bits_payload_data;
  wire [1:0] Queue_4_1_io_count;
  wire  Queue_5_1_clk;
  wire  Queue_5_1_reset;
  wire  Queue_5_1_io_enq_ready;
  wire  Queue_5_1_io_enq_valid;
  wire [1:0] Queue_5_1_io_enq_bits_header_src;
  wire [1:0] Queue_5_1_io_enq_bits_header_dst;
  wire [2:0] Queue_5_1_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_5_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_5_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_5_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_5_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_5_1_io_enq_bits_payload_data;
  wire  Queue_5_1_io_deq_ready;
  wire  Queue_5_1_io_deq_valid;
  wire [1:0] Queue_5_1_io_deq_bits_header_src;
  wire [1:0] Queue_5_1_io_deq_bits_header_dst;
  wire [2:0] Queue_5_1_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_5_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_5_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_5_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_5_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_5_1_io_deq_bits_payload_data;
  wire [1:0] Queue_5_1_io_count;
  Queue_2 Queue_2_1 (
    .clk(Queue_2_1_clk),
    .reset(Queue_2_1_reset),
    .io_enq_ready(Queue_2_1_io_enq_ready),
    .io_enq_valid(Queue_2_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_2_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_2_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_2_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_2_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_2_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_2_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_2_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_2_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_2_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_2_1_io_deq_ready),
    .io_deq_valid(Queue_2_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_2_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_2_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_2_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_2_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_2_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_2_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_2_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_2_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_2_1_io_deq_bits_payload_data),
    .io_count(Queue_2_1_io_count)
  );
  Queue_3 Queue_3_1 (
    .clk(Queue_3_1_clk),
    .reset(Queue_3_1_reset),
    .io_enq_ready(Queue_3_1_io_enq_ready),
    .io_enq_valid(Queue_3_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_3_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_3_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_3_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_3_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_3_1_io_deq_ready),
    .io_deq_valid(Queue_3_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_3_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_3_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_3_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_3_1_io_deq_bits_payload_p_type),
    .io_count(Queue_3_1_io_count)
  );
  Queue_4 Queue_4_1 (
    .clk(Queue_4_1_clk),
    .reset(Queue_4_1_reset),
    .io_enq_ready(Queue_4_1_io_enq_ready),
    .io_enq_valid(Queue_4_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_4_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_4_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_4_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_4_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_4_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_4_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_4_1_io_deq_ready),
    .io_deq_valid(Queue_4_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_4_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_4_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_4_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_4_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_4_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_4_1_io_deq_bits_payload_data),
    .io_count(Queue_4_1_io_count)
  );
  Queue_5 Queue_5_1 (
    .clk(Queue_5_1_clk),
    .reset(Queue_5_1_reset),
    .io_enq_ready(Queue_5_1_io_enq_ready),
    .io_enq_valid(Queue_5_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_5_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_5_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_5_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_5_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_5_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_5_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_5_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_5_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_5_1_io_deq_ready),
    .io_deq_valid(Queue_5_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_5_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_5_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_5_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_5_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_5_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_5_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_5_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_5_1_io_deq_bits_payload_data),
    .io_count(Queue_5_1_io_count)
  );
  assign io_client_acquire_ready = Queue_2_1_io_enq_ready;
  assign io_client_grant_valid = Queue_5_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_5_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_5_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_5_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_5_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_5_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_5_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_5_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_5_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_3_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_3_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_3_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_3_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_3_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_4_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_2_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_2_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_2_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_2_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_2_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_2_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_2_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_2_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_2_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_2_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_5_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_3_1_io_enq_ready;
  assign io_manager_release_valid = Queue_4_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_4_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_4_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_4_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_4_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_4_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_4_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_4_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_4_1_io_deq_bits_payload_data;
  assign Queue_2_1_clk = clk;
  assign Queue_2_1_reset = reset;
  assign Queue_2_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_2_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_2_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_2_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_2_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_2_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_2_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_2_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_2_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_2_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_2_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_3_1_clk = clk;
  assign Queue_3_1_reset = reset;
  assign Queue_3_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_3_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_3_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_3_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_3_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_3_1_io_deq_ready = io_client_probe_ready;
  assign Queue_4_1_clk = clk;
  assign Queue_4_1_reset = reset;
  assign Queue_4_1_io_enq_valid = io_client_release_valid;
  assign Queue_4_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_4_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_4_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_4_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_4_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_4_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_4_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_4_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_4_1_io_deq_ready = io_manager_release_ready;
  assign Queue_5_1_clk = clk;
  assign Queue_5_1_reset = reset;
  assign Queue_5_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_5_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_5_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_5_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_5_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_5_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_5_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_5_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_5_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_5_1_io_deq_ready = io_client_grant_ready;
endmodule
module ClientTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [10:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [25:0] io_client_probe_bits_addr_block,
  output [1:0] io_client_probe_bits_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_addr_beat,
  input  [25:0] io_client_release_bits_addr_block,
  input  [1:0] io_client_release_bits_client_xact_id,
  input   io_client_release_bits_voluntary,
  input  [2:0] io_client_release_bits_r_type,
  input  [63:0] io_client_release_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  output  io_client_grant_bits_manager_id,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_manager_xact_id,
  input   io_client_finish_bits_manager_id,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [10:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [10:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3894;
  wire  T_3896;
  wire  T_3898;
  wire  T_3899;
  wire  T_3902;
  wire  rel_with_header_ready;
  wire  rel_with_header_valid;
  wire [1:0] rel_with_header_bits_header_src;
  wire [1:0] rel_with_header_bits_header_dst;
  wire [2:0] rel_with_header_bits_payload_addr_beat;
  wire [25:0] rel_with_header_bits_payload_addr_block;
  wire [1:0] rel_with_header_bits_payload_client_xact_id;
  wire  rel_with_header_bits_payload_voluntary;
  wire [2:0] rel_with_header_bits_payload_r_type;
  wire [63:0] rel_with_header_bits_payload_data;
  wire [31:0] GEN_1;
  wire [31:0] T_4464;
  wire  T_4466;
  wire  T_4468;
  wire  T_4469;
  wire  T_4472;
  wire  fin_with_header_ready;
  wire  fin_with_header_valid;
  wire [1:0] fin_with_header_bits_header_src;
  wire [1:0] fin_with_header_bits_header_dst;
  wire [2:0] fin_with_header_bits_payload_manager_xact_id;
  wire  fin_with_header_bits_payload_manager_id;
  wire  prb_without_header_ready;
  wire  prb_without_header_valid;
  wire [25:0] prb_without_header_bits_addr_block;
  wire [1:0] prb_without_header_bits_p_type;
  wire  gnt_without_header_ready;
  wire  gnt_without_header_valid;
  wire [2:0] gnt_without_header_bits_addr_beat;
  wire [1:0] gnt_without_header_bits_client_xact_id;
  wire [2:0] gnt_without_header_bits_manager_xact_id;
  wire  gnt_without_header_bits_is_builtin_type;
  wire [3:0] gnt_without_header_bits_g_type;
  wire [63:0] gnt_without_header_bits_data;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_probe_valid = prb_without_header_valid;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign io_client_release_ready = rel_with_header_ready;
  assign io_client_grant_valid = gnt_without_header_valid;
  assign io_client_grant_bits_addr_beat = gnt_without_header_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = gnt_without_header_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = gnt_without_header_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = gnt_without_header_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = gnt_without_header_bits_g_type;
  assign io_client_grant_bits_data = gnt_without_header_bits_data;
  assign io_client_grant_bits_manager_id = io_network_grant_bits_header_src[0];
  assign io_client_finish_ready = fin_with_header_ready;
  assign io_network_acquire_valid = acq_with_header_valid;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = gnt_without_header_ready;
  assign io_network_finish_valid = fin_with_header_valid;
  assign io_network_finish_bits_header_src = fin_with_header_bits_header_src;
  assign io_network_finish_bits_header_dst = fin_with_header_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = fin_with_header_bits_payload_manager_xact_id;
  assign io_network_probe_ready = prb_without_header_ready;
  assign io_network_release_valid = rel_with_header_valid;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign acq_with_header_ready = io_network_acquire_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h0;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3902};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3894 = GEN_0 << 6;
  assign T_3896 = 32'h80000000 <= T_3894;
  assign T_3898 = T_3894 < 32'h90000000;
  assign T_3899 = T_3896 & T_3898;
  assign T_3902 = T_3899 ? 1'h0 : 1'h1;
  assign rel_with_header_ready = io_network_release_ready;
  assign rel_with_header_valid = io_client_release_valid;
  assign rel_with_header_bits_header_src = 2'h0;
  assign rel_with_header_bits_header_dst = {{1'd0}, T_4472};
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign GEN_1 = {{6'd0}, io_client_release_bits_addr_block};
  assign T_4464 = GEN_1 << 6;
  assign T_4466 = 32'h80000000 <= T_4464;
  assign T_4468 = T_4464 < 32'h90000000;
  assign T_4469 = T_4466 & T_4468;
  assign T_4472 = T_4469 ? 1'h0 : 1'h1;
  assign fin_with_header_ready = io_network_finish_ready;
  assign fin_with_header_valid = io_client_finish_valid;
  assign fin_with_header_bits_header_src = 2'h0;
  assign fin_with_header_bits_header_dst = {{1'd0}, io_client_finish_bits_manager_id};
  assign fin_with_header_bits_payload_manager_xact_id = io_client_finish_bits_manager_xact_id;
  assign fin_with_header_bits_payload_manager_id = io_client_finish_bits_manager_id;
  assign prb_without_header_ready = io_client_probe_ready;
  assign prb_without_header_valid = io_network_probe_valid;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign gnt_without_header_ready = io_client_grant_ready;
  assign gnt_without_header_valid = io_network_grant_valid;
  assign gnt_without_header_bits_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign gnt_without_header_bits_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign gnt_without_header_bits_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign gnt_without_header_bits_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign gnt_without_header_bits_g_type = io_network_grant_bits_payload_g_type;
  assign gnt_without_header_bits_data = io_network_grant_bits_payload_data;
endmodule
module TileLinkEnqueuer_1(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_6_1_clk;
  wire  Queue_6_1_reset;
  wire  Queue_6_1_io_enq_ready;
  wire  Queue_6_1_io_enq_valid;
  wire [1:0] Queue_6_1_io_enq_bits_header_src;
  wire [1:0] Queue_6_1_io_enq_bits_header_dst;
  wire [25:0] Queue_6_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_6_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_6_1_io_enq_bits_payload_addr_beat;
  wire  Queue_6_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_6_1_io_enq_bits_payload_a_type;
  wire [10:0] Queue_6_1_io_enq_bits_payload_union;
  wire [63:0] Queue_6_1_io_enq_bits_payload_data;
  wire  Queue_6_1_io_deq_ready;
  wire  Queue_6_1_io_deq_valid;
  wire [1:0] Queue_6_1_io_deq_bits_header_src;
  wire [1:0] Queue_6_1_io_deq_bits_header_dst;
  wire [25:0] Queue_6_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_6_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_6_1_io_deq_bits_payload_addr_beat;
  wire  Queue_6_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_6_1_io_deq_bits_payload_a_type;
  wire [10:0] Queue_6_1_io_deq_bits_payload_union;
  wire [63:0] Queue_6_1_io_deq_bits_payload_data;
  wire  Queue_6_1_io_count;
  wire  Queue_7_1_clk;
  wire  Queue_7_1_reset;
  wire  Queue_7_1_io_enq_ready;
  wire  Queue_7_1_io_enq_valid;
  wire [1:0] Queue_7_1_io_enq_bits_header_src;
  wire [1:0] Queue_7_1_io_enq_bits_header_dst;
  wire [25:0] Queue_7_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_7_1_io_enq_bits_payload_p_type;
  wire  Queue_7_1_io_deq_ready;
  wire  Queue_7_1_io_deq_valid;
  wire [1:0] Queue_7_1_io_deq_bits_header_src;
  wire [1:0] Queue_7_1_io_deq_bits_header_dst;
  wire [25:0] Queue_7_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_7_1_io_deq_bits_payload_p_type;
  wire  Queue_7_1_io_count;
  wire  Queue_8_1_clk;
  wire  Queue_8_1_reset;
  wire  Queue_8_1_io_enq_ready;
  wire  Queue_8_1_io_enq_valid;
  wire [1:0] Queue_8_1_io_enq_bits_header_src;
  wire [1:0] Queue_8_1_io_enq_bits_header_dst;
  wire [2:0] Queue_8_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_8_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_8_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_8_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_8_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_8_1_io_enq_bits_payload_data;
  wire  Queue_8_1_io_deq_ready;
  wire  Queue_8_1_io_deq_valid;
  wire [1:0] Queue_8_1_io_deq_bits_header_src;
  wire [1:0] Queue_8_1_io_deq_bits_header_dst;
  wire [2:0] Queue_8_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_8_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_8_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_8_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_8_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_8_1_io_deq_bits_payload_data;
  wire [1:0] Queue_8_1_io_count;
  wire  Queue_9_1_clk;
  wire  Queue_9_1_reset;
  wire  Queue_9_1_io_enq_ready;
  wire  Queue_9_1_io_enq_valid;
  wire [1:0] Queue_9_1_io_enq_bits_header_src;
  wire [1:0] Queue_9_1_io_enq_bits_header_dst;
  wire [2:0] Queue_9_1_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_9_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_9_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_9_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_9_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_9_1_io_enq_bits_payload_data;
  wire  Queue_9_1_io_deq_ready;
  wire  Queue_9_1_io_deq_valid;
  wire [1:0] Queue_9_1_io_deq_bits_header_src;
  wire [1:0] Queue_9_1_io_deq_bits_header_dst;
  wire [2:0] Queue_9_1_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_9_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_9_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_9_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_9_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_9_1_io_deq_bits_payload_data;
  wire [1:0] Queue_9_1_io_count;
  Queue_2 Queue_6_1 (
    .clk(Queue_6_1_clk),
    .reset(Queue_6_1_reset),
    .io_enq_ready(Queue_6_1_io_enq_ready),
    .io_enq_valid(Queue_6_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_6_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_6_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_6_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_6_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_6_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_6_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_6_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_6_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_6_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_6_1_io_deq_ready),
    .io_deq_valid(Queue_6_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_6_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_6_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_6_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_6_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_6_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_6_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_6_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_6_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_6_1_io_deq_bits_payload_data),
    .io_count(Queue_6_1_io_count)
  );
  Queue_3 Queue_7_1 (
    .clk(Queue_7_1_clk),
    .reset(Queue_7_1_reset),
    .io_enq_ready(Queue_7_1_io_enq_ready),
    .io_enq_valid(Queue_7_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_7_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_7_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_7_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_7_1_io_deq_ready),
    .io_deq_valid(Queue_7_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_7_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_7_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_7_1_io_deq_bits_payload_p_type),
    .io_count(Queue_7_1_io_count)
  );
  Queue_4 Queue_8_1 (
    .clk(Queue_8_1_clk),
    .reset(Queue_8_1_reset),
    .io_enq_ready(Queue_8_1_io_enq_ready),
    .io_enq_valid(Queue_8_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_8_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_8_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_8_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_8_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_8_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_8_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_8_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_8_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_8_1_io_deq_ready),
    .io_deq_valid(Queue_8_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_8_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_8_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_8_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_8_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_8_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_8_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_8_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_8_1_io_deq_bits_payload_data),
    .io_count(Queue_8_1_io_count)
  );
  Queue_5 Queue_9_1 (
    .clk(Queue_9_1_clk),
    .reset(Queue_9_1_reset),
    .io_enq_ready(Queue_9_1_io_enq_ready),
    .io_enq_valid(Queue_9_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_9_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_9_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_9_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_9_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_9_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_9_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_9_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_9_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_9_1_io_deq_ready),
    .io_deq_valid(Queue_9_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_9_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_9_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_9_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_9_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_9_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_9_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_9_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_9_1_io_deq_bits_payload_data),
    .io_count(Queue_9_1_io_count)
  );
  assign io_client_acquire_ready = Queue_6_1_io_enq_ready;
  assign io_client_grant_valid = Queue_9_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_9_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_9_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_9_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_9_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_9_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_9_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_9_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_9_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_7_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_7_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_7_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_7_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_7_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_8_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_6_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_6_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_6_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_6_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_6_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_6_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_6_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_6_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_6_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_6_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_9_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_7_1_io_enq_ready;
  assign io_manager_release_valid = Queue_8_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_8_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_8_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_8_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_8_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_8_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_8_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_8_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_8_1_io_deq_bits_payload_data;
  assign Queue_6_1_clk = clk;
  assign Queue_6_1_reset = reset;
  assign Queue_6_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_6_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_6_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_6_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_6_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_6_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_6_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_6_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_6_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_6_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_6_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_7_1_clk = clk;
  assign Queue_7_1_reset = reset;
  assign Queue_7_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_7_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_7_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_7_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_7_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_7_1_io_deq_ready = io_client_probe_ready;
  assign Queue_8_1_clk = clk;
  assign Queue_8_1_reset = reset;
  assign Queue_8_1_io_enq_valid = io_client_release_valid;
  assign Queue_8_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_8_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_8_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_8_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_8_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_8_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_8_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_8_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_8_1_io_deq_ready = io_manager_release_ready;
  assign Queue_9_1_clk = clk;
  assign Queue_9_1_reset = reset;
  assign Queue_9_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_9_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_9_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_9_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_9_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_9_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_9_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_9_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_9_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_9_1_io_deq_ready = io_client_grant_ready;
endmodule
module FinishQueue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output [1:0] io_count
);
  reg [2:0] ram_manager_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [2:0] ram_manager_xact_id_T_264_data;
  wire  ram_manager_xact_id_T_264_addr;
  wire  ram_manager_xact_id_T_264_en;
  wire [2:0] ram_manager_xact_id_T_226_data;
  wire  ram_manager_xact_id_T_226_addr;
  wire  ram_manager_xact_id_T_226_mask;
  wire  ram_manager_xact_id_T_226_en;
  reg  ram_manager_id [0:1];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_264_data;
  wire  ram_manager_id_T_264_addr;
  wire  ram_manager_id_T_264_en;
  wire  ram_manager_id_T_226_data;
  wire  ram_manager_id_T_226_addr;
  wire  ram_manager_id_T_226_mask;
  wire  ram_manager_id_T_226_en;
  reg  T_218;
  reg [31:0] GEN_2;
  reg  T_220;
  reg [31:0] GEN_3;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  ptr_match;
  wire  T_223;
  wire  empty;
  wire  full;
  wire  T_224;
  wire  do_enq;
  wire  T_225;
  wire  do_deq;
  wire [1:0] T_252;
  wire  T_253;
  wire  GEN_7;
  wire [1:0] T_257;
  wire  T_258;
  wire  GEN_8;
  wire  T_259;
  wire  GEN_9;
  wire  T_261;
  wire  T_263;
  wire [1:0] T_287;
  wire  ptr_diff;
  wire  T_288;
  wire [1:0] T_289;
  assign io_enq_ready = T_263;
  assign io_deq_valid = T_261;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_264_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_264_data;
  assign io_count = T_289;
  assign ram_manager_xact_id_T_264_addr = T_220;
  assign ram_manager_xact_id_T_264_en = 1'h1;
  assign ram_manager_xact_id_T_264_data = ram_manager_xact_id[ram_manager_xact_id_T_264_addr];
  assign ram_manager_xact_id_T_226_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_226_addr = T_218;
  assign ram_manager_xact_id_T_226_mask = do_enq;
  assign ram_manager_xact_id_T_226_en = do_enq;
  assign ram_manager_id_T_264_addr = T_220;
  assign ram_manager_id_T_264_en = 1'h1;
  assign ram_manager_id_T_264_data = ram_manager_id[ram_manager_id_T_264_addr];
  assign ram_manager_id_T_226_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_226_addr = T_218;
  assign ram_manager_id_T_226_mask = do_enq;
  assign ram_manager_id_T_226_en = do_enq;
  assign ptr_match = T_218 == T_220;
  assign T_223 = maybe_full == 1'h0;
  assign empty = ptr_match & T_223;
  assign full = ptr_match & maybe_full;
  assign T_224 = io_enq_ready & io_enq_valid;
  assign do_enq = T_224;
  assign T_225 = io_deq_ready & io_deq_valid;
  assign do_deq = T_225;
  assign T_252 = T_218 + 1'h1;
  assign T_253 = T_252[0:0];
  assign GEN_7 = do_enq ? T_253 : T_218;
  assign T_257 = T_220 + 1'h1;
  assign T_258 = T_257[0:0];
  assign GEN_8 = do_deq ? T_258 : T_220;
  assign T_259 = do_enq != do_deq;
  assign GEN_9 = T_259 ? do_enq : maybe_full;
  assign T_261 = empty == 1'h0;
  assign T_263 = full == 1'h0;
  assign T_287 = T_218 - T_220;
  assign ptr_diff = T_287[0:0];
  assign T_288 = maybe_full & ptr_match;
  assign T_289 = {T_288,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[2:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_218 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  T_220 = GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_226_en & ram_manager_xact_id_T_226_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_226_addr] <= ram_manager_xact_id_T_226_data;
    end
    if(ram_manager_id_T_226_en & ram_manager_id_T_226_mask) begin
      ram_manager_id[ram_manager_id_T_226_addr] <= ram_manager_id_T_226_data;
    end
    if(reset) begin
      T_218 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_218 <= T_253;
      end
    end
    if(reset) begin
      T_220 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_220 <= T_258;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_259) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module FinishUnit(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [1:0] io_grant_bits_header_src,
  input  [1:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input  [1:0] io_grant_bits_payload_client_xact_id,
  input  [2:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output [1:0] io_refill_bits_client_xact_id,
  output [2:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [1:0] io_finish_bits_header_src,
  output [1:0] io_finish_bits_header_dst,
  output [2:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1035;
  wire [2:0] T_1044_0;
  wire [3:0] GEN_1;
  wire  T_1046;
  wire  T_1047;
  wire  T_1048;
  wire  T_1050;
  reg [2:0] T_1052;
  reg [31:0] GEN_3;
  wire  T_1054;
  wire [3:0] T_1056;
  wire [2:0] T_1057;
  wire [2:0] GEN_0;
  wire  T_1058;
  wire  T_1060;
  wire  FinishQueue_3_1_clk;
  wire  FinishQueue_3_1_reset;
  wire  FinishQueue_3_1_io_enq_ready;
  wire  FinishQueue_3_1_io_enq_valid;
  wire [2:0] FinishQueue_3_1_io_enq_bits_manager_xact_id;
  wire  FinishQueue_3_1_io_enq_bits_manager_id;
  wire  FinishQueue_3_1_io_deq_ready;
  wire  FinishQueue_3_1_io_deq_valid;
  wire [2:0] FinishQueue_3_1_io_deq_bits_manager_xact_id;
  wire  FinishQueue_3_1_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_3_1_io_count;
  wire  T_1090;
  wire  T_1092;
  wire  T_1094;
  wire [2:0] T_1102_0;
  wire [3:0] GEN_2;
  wire  T_1104;
  wire  T_1106;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire [2:0] T_1134_manager_xact_id;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1182;
  FinishQueue_3 FinishQueue_3_1 (
    .clk(FinishQueue_3_1_clk),
    .reset(FinishQueue_3_1_reset),
    .io_enq_ready(FinishQueue_3_1_io_enq_ready),
    .io_enq_valid(FinishQueue_3_1_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_3_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_3_1_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_3_1_io_deq_ready),
    .io_deq_valid(FinishQueue_3_1_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_3_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_3_1_io_deq_bits_manager_id),
    .io_count(FinishQueue_3_1_io_count)
  );
  assign io_grant_ready = T_1182;
  assign io_refill_valid = T_1169;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_3_1_io_deq_valid;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_bits_header_dst = {{1'd0}, FinishQueue_3_1_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_3_1_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_3_1_io_enq_ready;
  assign T_1035 = io_grant_ready & io_grant_valid;
  assign T_1044_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1044_0};
  assign T_1046 = io_grant_bits_payload_g_type == GEN_1;
  assign T_1047 = io_grant_bits_payload_g_type == 4'h0;
  assign T_1048 = io_grant_bits_payload_is_builtin_type ? T_1046 : T_1047;
  assign T_1050 = T_1035 & T_1048;
  assign T_1054 = T_1052 == 3'h7;
  assign T_1056 = T_1052 + 3'h1;
  assign T_1057 = T_1056[2:0];
  assign GEN_0 = T_1050 ? T_1057 : T_1052;
  assign T_1058 = T_1050 & T_1054;
  assign T_1060 = T_1048 ? T_1058 : T_1035;
  assign FinishQueue_3_1_clk = clk;
  assign FinishQueue_3_1_reset = reset;
  assign FinishQueue_3_1_io_enq_valid = T_1111;
  assign FinishQueue_3_1_io_enq_bits_manager_xact_id = T_1134_manager_xact_id;
  assign FinishQueue_3_1_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_3_1_io_deq_ready = io_finish_ready;
  assign T_1090 = io_grant_bits_payload_is_builtin_type & T_1047;
  assign T_1092 = T_1090 == 1'h0;
  assign T_1094 = T_1035 & T_1092;
  assign T_1102_0 = 3'h5;
  assign GEN_2 = {{1'd0}, T_1102_0};
  assign T_1104 = io_grant_bits_payload_g_type == GEN_2;
  assign T_1106 = io_grant_bits_payload_is_builtin_type ? T_1104 : T_1047;
  assign T_1109 = T_1106 == 1'h0;
  assign T_1110 = T_1109 | T_1060;
  assign T_1111 = T_1094 & T_1110;
  assign T_1134_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1167 = T_1092 == 1'h0;
  assign T_1168 = FinishQueue_3_1_io_enq_ready | T_1167;
  assign T_1169 = T_1168 & io_grant_valid;
  assign T_1182 = T_1168 & io_refill_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  T_1052 = GEN_3[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1052 <= 3'h0;
    end else begin
      if(T_1050) begin
        T_1052 <= T_1057;
      end
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [10:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [10:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [1:0] finisher_io_grant_bits_header_src;
  wire [1:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire [1:0] finisher_io_grant_bits_payload_client_xact_id;
  wire [2:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire [1:0] finisher_io_refill_bits_client_xact_id;
  wire [2:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [1:0] finisher_io_finish_bits_header_src;
  wire [1:0] finisher_io_finish_bits_header_dst;
  wire [2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [10:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3330;
  wire  T_3332;
  wire  T_3334;
  wire  T_3335;
  wire  T_3338;
  wire  T_3339;
  wire  T_3340;
  wire [1:0] GEN_1;
  reg [31:0] GEN_9;
  wire [1:0] GEN_2;
  reg [31:0] GEN_10;
  wire [2:0] GEN_3;
  reg [31:0] GEN_11;
  wire [25:0] GEN_4;
  reg [31:0] GEN_12;
  wire [1:0] GEN_5;
  reg [31:0] GEN_13;
  wire  GEN_6;
  reg [31:0] GEN_14;
  wire [2:0] GEN_7;
  reg [31:0] GEN_15;
  wire [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3339;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3340;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h1;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3338};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3330 = GEN_0 << 6;
  assign T_3332 = 32'h80000000 <= T_3330;
  assign T_3334 = T_3330 < 32'h90000000;
  assign T_3335 = T_3332 & T_3334;
  assign T_3338 = T_3335 ? 1'h0 : 1'h1;
  assign T_3339 = acq_with_header_valid & finisher_io_ready;
  assign T_3340 = io_network_acquire_ready & finisher_io_ready;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_9[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_10[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_12[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_13[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_15[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_16[63:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_9 = {1{$random}};
  GEN_10 = {1{$random}};
  GEN_11 = {1{$random}};
  GEN_12 = {1{$random}};
  GEN_13 = {1{$random}};
  GEN_14 = {1{$random}};
  GEN_15 = {1{$random}};
  GEN_16 = {2{$random}};
  end
`endif
endmodule
module ManagerTileLinkNetworkPort(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [10:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [10:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire [1:0] T_6043_bits_payload_client_xact_id;
  wire [2:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire [1:0] T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [10:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire [1:0] T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [2:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h0;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h0;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module TileLinkEnqueuer_2(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [10:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [10:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  assign io_client_acquire_ready = io_manager_acquire_ready;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
endmodule
module ManagerTileLinkNetworkPort_1(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [10:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [10:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire [1:0] T_6043_bits_payload_client_xact_id;
  wire [2:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire [1:0] T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [10:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire [1:0] T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [2:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h1;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h1;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module LockingRRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [10:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [10:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [10:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [10:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_is_builtin_type,
  output [2:0] io_out_bits_payload_a_type,
  output [10:0] io_out_bits_payload_union,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [2:0] GEN_0_bits_payload_a_type;
  wire [10:0] GEN_0_bits_payload_union;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [25:0] GEN_14;
  wire [1:0] GEN_15;
  wire [2:0] GEN_16;
  wire  GEN_17;
  wire [2:0] GEN_18;
  wire [10:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [25:0] GEN_25;
  wire [1:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire [10:0] GEN_30;
  wire [63:0] GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  wire [25:0] GEN_36;
  wire [1:0] GEN_37;
  wire [2:0] GEN_38;
  wire  GEN_39;
  wire [2:0] GEN_40;
  wire [10:0] GEN_41;
  wire [63:0] GEN_42;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire [1:0] GEN_1_bits_payload_client_xact_id;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire  GEN_1_bits_payload_is_builtin_type;
  wire [2:0] GEN_1_bits_payload_a_type;
  wire [10:0] GEN_1_bits_payload_union;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire [1:0] GEN_2_bits_payload_client_xact_id;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire  GEN_2_bits_payload_is_builtin_type;
  wire [2:0] GEN_2_bits_payload_a_type;
  wire [10:0] GEN_2_bits_payload_union;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire [1:0] GEN_3_bits_payload_client_xact_id;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire  GEN_3_bits_payload_is_builtin_type;
  wire [2:0] GEN_3_bits_payload_a_type;
  wire [10:0] GEN_3_bits_payload_union;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire [1:0] GEN_4_bits_payload_client_xact_id;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire  GEN_4_bits_payload_is_builtin_type;
  wire [2:0] GEN_4_bits_payload_a_type;
  wire [10:0] GEN_4_bits_payload_union;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [25:0] GEN_5_bits_payload_addr_block;
  wire [1:0] GEN_5_bits_payload_client_xact_id;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire  GEN_5_bits_payload_is_builtin_type;
  wire [2:0] GEN_5_bits_payload_a_type;
  wire [10:0] GEN_5_bits_payload_union;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [25:0] GEN_6_bits_payload_addr_block;
  wire [1:0] GEN_6_bits_payload_client_xact_id;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire  GEN_6_bits_payload_is_builtin_type;
  wire [2:0] GEN_6_bits_payload_a_type;
  wire [10:0] GEN_6_bits_payload_union;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [25:0] GEN_7_bits_payload_addr_block;
  wire [1:0] GEN_7_bits_payload_client_xact_id;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire  GEN_7_bits_payload_is_builtin_type;
  wire [2:0] GEN_7_bits_payload_a_type;
  wire [10:0] GEN_7_bits_payload_union;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [25:0] GEN_8_bits_payload_addr_block;
  wire [1:0] GEN_8_bits_payload_client_xact_id;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire  GEN_8_bits_payload_is_builtin_type;
  wire [2:0] GEN_8_bits_payload_a_type;
  wire [10:0] GEN_8_bits_payload_union;
  wire [63:0] GEN_8_bits_payload_data;
  wire  GEN_9_ready;
  wire  GEN_9_valid;
  wire [1:0] GEN_9_bits_header_src;
  wire [1:0] GEN_9_bits_header_dst;
  wire [25:0] GEN_9_bits_payload_addr_block;
  wire [1:0] GEN_9_bits_payload_client_xact_id;
  wire [2:0] GEN_9_bits_payload_addr_beat;
  wire  GEN_9_bits_payload_is_builtin_type;
  wire [2:0] GEN_9_bits_payload_a_type;
  wire [10:0] GEN_9_bits_payload_union;
  wire [63:0] GEN_9_bits_payload_data;
  reg [2:0] T_1134;
  reg [31:0] GEN_0;
  reg [1:0] T_1136;
  reg [31:0] GEN_1;
  wire  T_1138;
  wire [2:0] T_1147_0;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire [3:0] T_1156;
  wire [2:0] T_1157;
  wire [1:0] GEN_340;
  wire [2:0] GEN_341;
  wire [1:0] GEN_342;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_343;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1165;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1173;
  wire  T_1175;
  wire  T_1177;
  wire  T_1179;
  wire  T_1181;
  wire  T_1183;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1190;
  wire  T_1191;
  wire  T_1193;
  wire  T_1194;
  wire  T_1195;
  wire  T_1197;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1205;
  wire  T_1206;
  wire  T_1207;
  wire [1:0] GEN_344;
  wire [1:0] GEN_345;
  wire [1:0] GEN_346;
  wire [1:0] GEN_347;
  wire [1:0] GEN_348;
  wire [1:0] GEN_349;
  assign io_in_0_ready = T_1195;
  assign io_in_1_ready = T_1199;
  assign io_in_2_ready = T_1203;
  assign io_in_3_ready = T_1207;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_block = GEN_3_bits_payload_addr_block;
  assign io_out_bits_payload_client_xact_id = GEN_4_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr_beat = GEN_5_bits_payload_addr_beat;
  assign io_out_bits_payload_is_builtin_type = GEN_6_bits_payload_is_builtin_type;
  assign io_out_bits_payload_a_type = GEN_7_bits_payload_a_type;
  assign io_out_bits_payload_union = GEN_8_bits_payload_union;
  assign io_out_bits_payload_data = GEN_9_bits_payload_data;
  assign io_chosen = GEN_342;
  assign choice = GEN_349;
  assign GEN_0_ready = GEN_32;
  assign GEN_0_valid = GEN_33;
  assign GEN_0_bits_header_src = GEN_34;
  assign GEN_0_bits_header_dst = GEN_35;
  assign GEN_0_bits_payload_addr_block = GEN_36;
  assign GEN_0_bits_payload_client_xact_id = GEN_37;
  assign GEN_0_bits_payload_addr_beat = GEN_38;
  assign GEN_0_bits_payload_is_builtin_type = GEN_39;
  assign GEN_0_bits_payload_a_type = GEN_40;
  assign GEN_0_bits_payload_union = GEN_41;
  assign GEN_0_bits_payload_data = GEN_42;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign GEN_19 = 2'h1 == io_chosen ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign GEN_20 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_ready : GEN_10;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_valid : GEN_11;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_13;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_15;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_16;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_17;
  assign GEN_29 = 2'h2 == io_chosen ? io_in_2_bits_payload_a_type : GEN_18;
  assign GEN_30 = 2'h2 == io_chosen ? io_in_2_bits_payload_union : GEN_19;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_20;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_ready : GEN_21;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_valid : GEN_22;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_23;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_24;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_25;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_26;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_27;
  assign GEN_39 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_28;
  assign GEN_40 = 2'h3 == io_chosen ? io_in_3_bits_payload_a_type : GEN_29;
  assign GEN_41 = 2'h3 == io_chosen ? io_in_3_bits_payload_union : GEN_30;
  assign GEN_42 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_31;
  assign GEN_1_ready = GEN_32;
  assign GEN_1_valid = GEN_33;
  assign GEN_1_bits_header_src = GEN_34;
  assign GEN_1_bits_header_dst = GEN_35;
  assign GEN_1_bits_payload_addr_block = GEN_36;
  assign GEN_1_bits_payload_client_xact_id = GEN_37;
  assign GEN_1_bits_payload_addr_beat = GEN_38;
  assign GEN_1_bits_payload_is_builtin_type = GEN_39;
  assign GEN_1_bits_payload_a_type = GEN_40;
  assign GEN_1_bits_payload_union = GEN_41;
  assign GEN_1_bits_payload_data = GEN_42;
  assign GEN_2_ready = GEN_32;
  assign GEN_2_valid = GEN_33;
  assign GEN_2_bits_header_src = GEN_34;
  assign GEN_2_bits_header_dst = GEN_35;
  assign GEN_2_bits_payload_addr_block = GEN_36;
  assign GEN_2_bits_payload_client_xact_id = GEN_37;
  assign GEN_2_bits_payload_addr_beat = GEN_38;
  assign GEN_2_bits_payload_is_builtin_type = GEN_39;
  assign GEN_2_bits_payload_a_type = GEN_40;
  assign GEN_2_bits_payload_union = GEN_41;
  assign GEN_2_bits_payload_data = GEN_42;
  assign GEN_3_ready = GEN_32;
  assign GEN_3_valid = GEN_33;
  assign GEN_3_bits_header_src = GEN_34;
  assign GEN_3_bits_header_dst = GEN_35;
  assign GEN_3_bits_payload_addr_block = GEN_36;
  assign GEN_3_bits_payload_client_xact_id = GEN_37;
  assign GEN_3_bits_payload_addr_beat = GEN_38;
  assign GEN_3_bits_payload_is_builtin_type = GEN_39;
  assign GEN_3_bits_payload_a_type = GEN_40;
  assign GEN_3_bits_payload_union = GEN_41;
  assign GEN_3_bits_payload_data = GEN_42;
  assign GEN_4_ready = GEN_32;
  assign GEN_4_valid = GEN_33;
  assign GEN_4_bits_header_src = GEN_34;
  assign GEN_4_bits_header_dst = GEN_35;
  assign GEN_4_bits_payload_addr_block = GEN_36;
  assign GEN_4_bits_payload_client_xact_id = GEN_37;
  assign GEN_4_bits_payload_addr_beat = GEN_38;
  assign GEN_4_bits_payload_is_builtin_type = GEN_39;
  assign GEN_4_bits_payload_a_type = GEN_40;
  assign GEN_4_bits_payload_union = GEN_41;
  assign GEN_4_bits_payload_data = GEN_42;
  assign GEN_5_ready = GEN_32;
  assign GEN_5_valid = GEN_33;
  assign GEN_5_bits_header_src = GEN_34;
  assign GEN_5_bits_header_dst = GEN_35;
  assign GEN_5_bits_payload_addr_block = GEN_36;
  assign GEN_5_bits_payload_client_xact_id = GEN_37;
  assign GEN_5_bits_payload_addr_beat = GEN_38;
  assign GEN_5_bits_payload_is_builtin_type = GEN_39;
  assign GEN_5_bits_payload_a_type = GEN_40;
  assign GEN_5_bits_payload_union = GEN_41;
  assign GEN_5_bits_payload_data = GEN_42;
  assign GEN_6_ready = GEN_32;
  assign GEN_6_valid = GEN_33;
  assign GEN_6_bits_header_src = GEN_34;
  assign GEN_6_bits_header_dst = GEN_35;
  assign GEN_6_bits_payload_addr_block = GEN_36;
  assign GEN_6_bits_payload_client_xact_id = GEN_37;
  assign GEN_6_bits_payload_addr_beat = GEN_38;
  assign GEN_6_bits_payload_is_builtin_type = GEN_39;
  assign GEN_6_bits_payload_a_type = GEN_40;
  assign GEN_6_bits_payload_union = GEN_41;
  assign GEN_6_bits_payload_data = GEN_42;
  assign GEN_7_ready = GEN_32;
  assign GEN_7_valid = GEN_33;
  assign GEN_7_bits_header_src = GEN_34;
  assign GEN_7_bits_header_dst = GEN_35;
  assign GEN_7_bits_payload_addr_block = GEN_36;
  assign GEN_7_bits_payload_client_xact_id = GEN_37;
  assign GEN_7_bits_payload_addr_beat = GEN_38;
  assign GEN_7_bits_payload_is_builtin_type = GEN_39;
  assign GEN_7_bits_payload_a_type = GEN_40;
  assign GEN_7_bits_payload_union = GEN_41;
  assign GEN_7_bits_payload_data = GEN_42;
  assign GEN_8_ready = GEN_32;
  assign GEN_8_valid = GEN_33;
  assign GEN_8_bits_header_src = GEN_34;
  assign GEN_8_bits_header_dst = GEN_35;
  assign GEN_8_bits_payload_addr_block = GEN_36;
  assign GEN_8_bits_payload_client_xact_id = GEN_37;
  assign GEN_8_bits_payload_addr_beat = GEN_38;
  assign GEN_8_bits_payload_is_builtin_type = GEN_39;
  assign GEN_8_bits_payload_a_type = GEN_40;
  assign GEN_8_bits_payload_union = GEN_41;
  assign GEN_8_bits_payload_data = GEN_42;
  assign GEN_9_ready = GEN_32;
  assign GEN_9_valid = GEN_33;
  assign GEN_9_bits_header_src = GEN_34;
  assign GEN_9_bits_header_dst = GEN_35;
  assign GEN_9_bits_payload_addr_block = GEN_36;
  assign GEN_9_bits_payload_client_xact_id = GEN_37;
  assign GEN_9_bits_payload_addr_beat = GEN_38;
  assign GEN_9_bits_payload_is_builtin_type = GEN_39;
  assign GEN_9_bits_payload_a_type = GEN_40;
  assign GEN_9_bits_payload_union = GEN_41;
  assign GEN_9_bits_payload_data = GEN_42;
  assign T_1138 = T_1134 != 3'h0;
  assign T_1147_0 = 3'h3;
  assign T_1149 = io_out_bits_payload_a_type == T_1147_0;
  assign T_1150 = io_out_bits_payload_is_builtin_type & T_1149;
  assign T_1151 = io_out_ready & io_out_valid;
  assign T_1152 = T_1151 & T_1150;
  assign T_1156 = T_1134 + 3'h1;
  assign T_1157 = T_1156[2:0];
  assign GEN_340 = T_1152 ? io_chosen : T_1136;
  assign GEN_341 = T_1152 ? T_1157 : T_1134;
  assign GEN_342 = T_1138 ? T_1136 : choice;
  assign GEN_343 = T_1151 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1165 = validMask_1 | validMask_2;
  assign T_1166 = T_1165 | validMask_3;
  assign T_1167 = T_1166 | io_in_0_valid;
  assign T_1168 = T_1167 | io_in_1_valid;
  assign T_1169 = T_1168 | io_in_2_valid;
  assign T_1173 = validMask_1 == 1'h0;
  assign T_1175 = T_1165 == 1'h0;
  assign T_1177 = T_1166 == 1'h0;
  assign T_1179 = T_1167 == 1'h0;
  assign T_1181 = T_1168 == 1'h0;
  assign T_1183 = T_1169 == 1'h0;
  assign T_1187 = grantMask_1 | T_1179;
  assign T_1188 = T_1173 & grantMask_2;
  assign T_1189 = T_1188 | T_1181;
  assign T_1190 = T_1175 & grantMask_3;
  assign T_1191 = T_1190 | T_1183;
  assign T_1193 = T_1136 == 2'h0;
  assign T_1194 = T_1138 ? T_1193 : T_1177;
  assign T_1195 = T_1194 & io_out_ready;
  assign T_1197 = T_1136 == 2'h1;
  assign T_1198 = T_1138 ? T_1197 : T_1187;
  assign T_1199 = T_1198 & io_out_ready;
  assign T_1201 = T_1136 == 2'h2;
  assign T_1202 = T_1138 ? T_1201 : T_1189;
  assign T_1203 = T_1202 & io_out_ready;
  assign T_1205 = T_1136 == 2'h3;
  assign T_1206 = T_1138 ? T_1205 : T_1191;
  assign T_1207 = T_1206 & io_out_ready;
  assign GEN_344 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_345 = io_in_1_valid ? 2'h1 : GEN_344;
  assign GEN_346 = io_in_0_valid ? 2'h0 : GEN_345;
  assign GEN_347 = validMask_3 ? 2'h3 : GEN_346;
  assign GEN_348 = validMask_2 ? 2'h2 : GEN_347;
  assign GEN_349 = validMask_1 ? 2'h1 : GEN_348;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1134 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1136 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1134 <= 3'h0;
    end else begin
      if(T_1152) begin
        T_1134 <= T_1157;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1152) begin
        T_1136 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1151) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [10:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [10:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [10:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [10:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_is_builtin_type,
  output [2:0] io_out_0_bits_payload_a_type,
  output [10:0] io_out_0_bits_payload_union,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_is_builtin_type,
  output [2:0] io_out_1_bits_payload_a_type,
  output [10:0] io_out_1_bits_payload_union,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_is_builtin_type,
  output [2:0] io_out_2_bits_payload_a_type,
  output [10:0] io_out_2_bits_payload_union,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_is_builtin_type,
  output [2:0] io_out_3_bits_payload_a_type,
  output [10:0] io_out_3_bits_payload_union,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_0_bits_payload_a_type;
  wire [10:0] arb_io_in_0_bits_payload_union;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_1_bits_payload_a_type;
  wire [10:0] arb_io_in_1_bits_payload_union;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_2_bits_payload_a_type;
  wire [10:0] arb_io_in_2_bits_payload_union;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_3_bits_payload_a_type;
  wire [10:0] arb_io_in_3_bits_payload_union;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [2:0] arb_io_out_bits_payload_a_type;
  wire [10:0] arb_io_out_bits_payload_union;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [2:0] GEN_0_bits_payload_a_type;
  wire [10:0] GEN_0_bits_payload_union;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [25:0] GEN_5;
  wire [1:0] GEN_6;
  wire [2:0] GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [10:0] GEN_10;
  wire [63:0] GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [25:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_18;
  wire  GEN_19;
  wire [2:0] GEN_20;
  wire [10:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [25:0] GEN_27;
  wire [1:0] GEN_28;
  wire [2:0] GEN_29;
  wire  GEN_30;
  wire [2:0] GEN_31;
  wire [10:0] GEN_32;
  wire [63:0] GEN_33;
  wire  T_1529;
  wire  T_1530;
  wire  T_1532;
  wire  T_1533;
  wire  T_1535;
  wire  T_1536;
  wire  T_1538;
  wire  T_1539;
  LockingRRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(arb_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(arb_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(arb_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(arb_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(arb_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(arb_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(arb_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(arb_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_a_type(arb_io_out_bits_payload_a_type),
    .io_out_bits_payload_union(arb_io_out_bits_payload_union),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1530;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1533;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1536;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1539;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_a_type = io_in_0_bits_payload_a_type;
  assign arb_io_in_0_bits_payload_union = io_in_0_bits_payload_union;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_a_type = io_in_1_bits_payload_a_type;
  assign arb_io_in_1_bits_payload_union = io_in_1_bits_payload_union;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_a_type = io_in_2_bits_payload_a_type;
  assign arb_io_in_2_bits_payload_union = io_in_2_bits_payload_union;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_a_type = io_in_3_bits_payload_a_type;
  assign arb_io_in_3_bits_payload_union = io_in_3_bits_payload_union;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_23;
  assign GEN_0_valid = GEN_24;
  assign GEN_0_bits_header_src = GEN_25;
  assign GEN_0_bits_header_dst = GEN_26;
  assign GEN_0_bits_payload_addr_block = GEN_27;
  assign GEN_0_bits_payload_client_xact_id = GEN_28;
  assign GEN_0_bits_payload_addr_beat = GEN_29;
  assign GEN_0_bits_payload_is_builtin_type = GEN_30;
  assign GEN_0_bits_payload_a_type = GEN_31;
  assign GEN_0_bits_payload_union = GEN_32;
  assign GEN_0_bits_payload_data = GEN_33;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_is_builtin_type : io_out_0_bits_payload_is_builtin_type;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_a_type : io_out_0_bits_payload_a_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_union : io_out_0_bits_payload_union;
  assign GEN_11 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_5;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_6;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_7;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_is_builtin_type : GEN_8;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_a_type : GEN_9;
  assign GEN_21 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_union : GEN_10;
  assign GEN_22 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_11;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_12;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_13;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_14;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_15;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_16;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_17;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_18;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_is_builtin_type : GEN_19;
  assign GEN_31 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_a_type : GEN_20;
  assign GEN_32 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_union : GEN_21;
  assign GEN_33 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_22;
  assign T_1529 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1530 = arb_io_out_valid & T_1529;
  assign T_1532 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1533 = arb_io_out_valid & T_1532;
  assign T_1535 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1536 = arb_io_out_valid & T_1535;
  assign T_1538 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1539 = arb_io_out_valid & T_1538;
endmodule
module LockingRRArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output  io_out_bits_payload_voluntary,
  output [2:0] io_out_bits_payload_r_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire  GEN_0_bits_payload_voluntary;
  wire [2:0] GEN_0_bits_payload_r_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_13;
  wire [25:0] GEN_14;
  wire [1:0] GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [63:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [2:0] GEN_23;
  wire [25:0] GEN_24;
  wire [1:0] GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_27;
  wire [63:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire [2:0] GEN_33;
  wire [25:0] GEN_34;
  wire [1:0] GEN_35;
  wire  GEN_36;
  wire [2:0] GEN_37;
  wire [63:0] GEN_38;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire [1:0] GEN_1_bits_payload_client_xact_id;
  wire  GEN_1_bits_payload_voluntary;
  wire [2:0] GEN_1_bits_payload_r_type;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire [1:0] GEN_2_bits_payload_client_xact_id;
  wire  GEN_2_bits_payload_voluntary;
  wire [2:0] GEN_2_bits_payload_r_type;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire [1:0] GEN_3_bits_payload_client_xact_id;
  wire  GEN_3_bits_payload_voluntary;
  wire [2:0] GEN_3_bits_payload_r_type;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire [1:0] GEN_4_bits_payload_client_xact_id;
  wire  GEN_4_bits_payload_voluntary;
  wire [2:0] GEN_4_bits_payload_r_type;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire [25:0] GEN_5_bits_payload_addr_block;
  wire [1:0] GEN_5_bits_payload_client_xact_id;
  wire  GEN_5_bits_payload_voluntary;
  wire [2:0] GEN_5_bits_payload_r_type;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire [25:0] GEN_6_bits_payload_addr_block;
  wire [1:0] GEN_6_bits_payload_client_xact_id;
  wire  GEN_6_bits_payload_voluntary;
  wire [2:0] GEN_6_bits_payload_r_type;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire [25:0] GEN_7_bits_payload_addr_block;
  wire [1:0] GEN_7_bits_payload_client_xact_id;
  wire  GEN_7_bits_payload_voluntary;
  wire [2:0] GEN_7_bits_payload_r_type;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire [25:0] GEN_8_bits_payload_addr_block;
  wire [1:0] GEN_8_bits_payload_client_xact_id;
  wire  GEN_8_bits_payload_voluntary;
  wire [2:0] GEN_8_bits_payload_r_type;
  wire [63:0] GEN_8_bits_payload_data;
  reg [2:0] T_1100;
  reg [31:0] GEN_0;
  reg [1:0] T_1102;
  reg [31:0] GEN_1;
  wire  T_1104;
  wire  T_1106;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1112;
  wire  T_1113;
  wire [3:0] T_1117;
  wire [2:0] T_1118;
  wire [1:0] GEN_279;
  wire [2:0] GEN_280;
  wire [1:0] GEN_281;
  reg [1:0] lastGrant;
  reg [31:0] GEN_2;
  wire [1:0] GEN_282;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1126;
  wire  T_1127;
  wire  T_1128;
  wire  T_1129;
  wire  T_1130;
  wire  T_1134;
  wire  T_1136;
  wire  T_1138;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1148;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1158;
  wire  T_1159;
  wire  T_1160;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire [1:0] GEN_283;
  wire [1:0] GEN_284;
  wire [1:0] GEN_285;
  wire [1:0] GEN_286;
  wire [1:0] GEN_287;
  wire [1:0] GEN_288;
  assign io_in_0_ready = T_1156;
  assign io_in_1_ready = T_1160;
  assign io_in_2_ready = T_1164;
  assign io_in_3_ready = T_1168;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_beat = GEN_3_bits_payload_addr_beat;
  assign io_out_bits_payload_addr_block = GEN_4_bits_payload_addr_block;
  assign io_out_bits_payload_client_xact_id = GEN_5_bits_payload_client_xact_id;
  assign io_out_bits_payload_voluntary = GEN_6_bits_payload_voluntary;
  assign io_out_bits_payload_r_type = GEN_7_bits_payload_r_type;
  assign io_out_bits_payload_data = GEN_8_bits_payload_data;
  assign io_chosen = GEN_281;
  assign choice = GEN_288;
  assign GEN_0_ready = GEN_29;
  assign GEN_0_valid = GEN_30;
  assign GEN_0_bits_header_src = GEN_31;
  assign GEN_0_bits_header_dst = GEN_32;
  assign GEN_0_bits_payload_addr_beat = GEN_33;
  assign GEN_0_bits_payload_addr_block = GEN_34;
  assign GEN_0_bits_payload_client_xact_id = GEN_35;
  assign GEN_0_bits_payload_voluntary = GEN_36;
  assign GEN_0_bits_payload_r_type = GEN_37;
  assign GEN_0_bits_payload_data = GEN_38;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_ready : GEN_9;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_11;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_12;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_13;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_15;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_voluntary : GEN_16;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_r_type : GEN_17;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_18;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_ready : GEN_19;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_valid : GEN_20;
  assign GEN_31 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_21;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_22;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_23;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_24;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_25;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_voluntary : GEN_26;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_r_type : GEN_27;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_28;
  assign GEN_1_ready = GEN_29;
  assign GEN_1_valid = GEN_30;
  assign GEN_1_bits_header_src = GEN_31;
  assign GEN_1_bits_header_dst = GEN_32;
  assign GEN_1_bits_payload_addr_beat = GEN_33;
  assign GEN_1_bits_payload_addr_block = GEN_34;
  assign GEN_1_bits_payload_client_xact_id = GEN_35;
  assign GEN_1_bits_payload_voluntary = GEN_36;
  assign GEN_1_bits_payload_r_type = GEN_37;
  assign GEN_1_bits_payload_data = GEN_38;
  assign GEN_2_ready = GEN_29;
  assign GEN_2_valid = GEN_30;
  assign GEN_2_bits_header_src = GEN_31;
  assign GEN_2_bits_header_dst = GEN_32;
  assign GEN_2_bits_payload_addr_beat = GEN_33;
  assign GEN_2_bits_payload_addr_block = GEN_34;
  assign GEN_2_bits_payload_client_xact_id = GEN_35;
  assign GEN_2_bits_payload_voluntary = GEN_36;
  assign GEN_2_bits_payload_r_type = GEN_37;
  assign GEN_2_bits_payload_data = GEN_38;
  assign GEN_3_ready = GEN_29;
  assign GEN_3_valid = GEN_30;
  assign GEN_3_bits_header_src = GEN_31;
  assign GEN_3_bits_header_dst = GEN_32;
  assign GEN_3_bits_payload_addr_beat = GEN_33;
  assign GEN_3_bits_payload_addr_block = GEN_34;
  assign GEN_3_bits_payload_client_xact_id = GEN_35;
  assign GEN_3_bits_payload_voluntary = GEN_36;
  assign GEN_3_bits_payload_r_type = GEN_37;
  assign GEN_3_bits_payload_data = GEN_38;
  assign GEN_4_ready = GEN_29;
  assign GEN_4_valid = GEN_30;
  assign GEN_4_bits_header_src = GEN_31;
  assign GEN_4_bits_header_dst = GEN_32;
  assign GEN_4_bits_payload_addr_beat = GEN_33;
  assign GEN_4_bits_payload_addr_block = GEN_34;
  assign GEN_4_bits_payload_client_xact_id = GEN_35;
  assign GEN_4_bits_payload_voluntary = GEN_36;
  assign GEN_4_bits_payload_r_type = GEN_37;
  assign GEN_4_bits_payload_data = GEN_38;
  assign GEN_5_ready = GEN_29;
  assign GEN_5_valid = GEN_30;
  assign GEN_5_bits_header_src = GEN_31;
  assign GEN_5_bits_header_dst = GEN_32;
  assign GEN_5_bits_payload_addr_beat = GEN_33;
  assign GEN_5_bits_payload_addr_block = GEN_34;
  assign GEN_5_bits_payload_client_xact_id = GEN_35;
  assign GEN_5_bits_payload_voluntary = GEN_36;
  assign GEN_5_bits_payload_r_type = GEN_37;
  assign GEN_5_bits_payload_data = GEN_38;
  assign GEN_6_ready = GEN_29;
  assign GEN_6_valid = GEN_30;
  assign GEN_6_bits_header_src = GEN_31;
  assign GEN_6_bits_header_dst = GEN_32;
  assign GEN_6_bits_payload_addr_beat = GEN_33;
  assign GEN_6_bits_payload_addr_block = GEN_34;
  assign GEN_6_bits_payload_client_xact_id = GEN_35;
  assign GEN_6_bits_payload_voluntary = GEN_36;
  assign GEN_6_bits_payload_r_type = GEN_37;
  assign GEN_6_bits_payload_data = GEN_38;
  assign GEN_7_ready = GEN_29;
  assign GEN_7_valid = GEN_30;
  assign GEN_7_bits_header_src = GEN_31;
  assign GEN_7_bits_header_dst = GEN_32;
  assign GEN_7_bits_payload_addr_beat = GEN_33;
  assign GEN_7_bits_payload_addr_block = GEN_34;
  assign GEN_7_bits_payload_client_xact_id = GEN_35;
  assign GEN_7_bits_payload_voluntary = GEN_36;
  assign GEN_7_bits_payload_r_type = GEN_37;
  assign GEN_7_bits_payload_data = GEN_38;
  assign GEN_8_ready = GEN_29;
  assign GEN_8_valid = GEN_30;
  assign GEN_8_bits_header_src = GEN_31;
  assign GEN_8_bits_header_dst = GEN_32;
  assign GEN_8_bits_payload_addr_beat = GEN_33;
  assign GEN_8_bits_payload_addr_block = GEN_34;
  assign GEN_8_bits_payload_client_xact_id = GEN_35;
  assign GEN_8_bits_payload_voluntary = GEN_36;
  assign GEN_8_bits_payload_r_type = GEN_37;
  assign GEN_8_bits_payload_data = GEN_38;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1106 = io_out_bits_payload_r_type == 3'h0;
  assign T_1107 = io_out_bits_payload_r_type == 3'h1;
  assign T_1108 = io_out_bits_payload_r_type == 3'h2;
  assign T_1109 = T_1106 | T_1107;
  assign T_1110 = T_1109 | T_1108;
  assign T_1112 = io_out_ready & io_out_valid;
  assign T_1113 = T_1112 & T_1110;
  assign T_1117 = T_1100 + 3'h1;
  assign T_1118 = T_1117[2:0];
  assign GEN_279 = T_1113 ? io_chosen : T_1102;
  assign GEN_280 = T_1113 ? T_1118 : T_1100;
  assign GEN_281 = T_1104 ? T_1102 : choice;
  assign GEN_282 = T_1112 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1126 = validMask_1 | validMask_2;
  assign T_1127 = T_1126 | validMask_3;
  assign T_1128 = T_1127 | io_in_0_valid;
  assign T_1129 = T_1128 | io_in_1_valid;
  assign T_1130 = T_1129 | io_in_2_valid;
  assign T_1134 = validMask_1 == 1'h0;
  assign T_1136 = T_1126 == 1'h0;
  assign T_1138 = T_1127 == 1'h0;
  assign T_1140 = T_1128 == 1'h0;
  assign T_1142 = T_1129 == 1'h0;
  assign T_1144 = T_1130 == 1'h0;
  assign T_1148 = grantMask_1 | T_1140;
  assign T_1149 = T_1134 & grantMask_2;
  assign T_1150 = T_1149 | T_1142;
  assign T_1151 = T_1136 & grantMask_3;
  assign T_1152 = T_1151 | T_1144;
  assign T_1154 = T_1102 == 2'h0;
  assign T_1155 = T_1104 ? T_1154 : T_1138;
  assign T_1156 = T_1155 & io_out_ready;
  assign T_1158 = T_1102 == 2'h1;
  assign T_1159 = T_1104 ? T_1158 : T_1148;
  assign T_1160 = T_1159 & io_out_ready;
  assign T_1162 = T_1102 == 2'h2;
  assign T_1163 = T_1104 ? T_1162 : T_1150;
  assign T_1164 = T_1163 & io_out_ready;
  assign T_1166 = T_1102 == 2'h3;
  assign T_1167 = T_1104 ? T_1166 : T_1152;
  assign T_1168 = T_1167 & io_out_ready;
  assign GEN_283 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_284 = io_in_1_valid ? 2'h1 : GEN_283;
  assign GEN_285 = io_in_0_valid ? 2'h0 : GEN_284;
  assign GEN_286 = validMask_3 ? 2'h3 : GEN_285;
  assign GEN_287 = validMask_2 ? 2'h2 : GEN_286;
  assign GEN_288 = validMask_1 ? 2'h1 : GEN_287;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1100 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1102 = GEN_1[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1113) begin
        T_1100 <= T_1118;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1113) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1112) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output  io_out_0_bits_payload_voluntary,
  output [2:0] io_out_0_bits_payload_r_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output  io_out_1_bits_payload_voluntary,
  output [2:0] io_out_1_bits_payload_r_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output  io_out_2_bits_payload_voluntary,
  output [2:0] io_out_2_bits_payload_r_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output  io_out_3_bits_payload_voluntary,
  output [2:0] io_out_3_bits_payload_r_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire  arb_io_in_0_bits_payload_voluntary;
  wire [2:0] arb_io_in_0_bits_payload_r_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire  arb_io_in_1_bits_payload_voluntary;
  wire [2:0] arb_io_in_1_bits_payload_r_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire  arb_io_in_2_bits_payload_voluntary;
  wire [2:0] arb_io_in_2_bits_payload_r_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire  arb_io_in_3_bits_payload_voluntary;
  wire [2:0] arb_io_in_3_bits_payload_r_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire  arb_io_out_bits_payload_voluntary;
  wire [2:0] arb_io_out_bits_payload_r_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire  GEN_0_bits_payload_voluntary;
  wire [2:0] GEN_0_bits_payload_r_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [2:0] GEN_5;
  wire [25:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [63:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire [25:0] GEN_16;
  wire [1:0] GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire [25:0] GEN_26;
  wire [1:0] GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire [63:0] GEN_30;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_1 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(arb_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(arb_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(arb_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(arb_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(arb_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(arb_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(arb_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(arb_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_voluntary(arb_io_out_bits_payload_voluntary),
    .io_out_bits_payload_r_type(arb_io_out_bits_payload_r_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_voluntary = io_in_0_bits_payload_voluntary;
  assign arb_io_in_0_bits_payload_r_type = io_in_0_bits_payload_r_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_voluntary = io_in_1_bits_payload_voluntary;
  assign arb_io_in_1_bits_payload_r_type = io_in_1_bits_payload_r_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_voluntary = io_in_2_bits_payload_voluntary;
  assign arb_io_in_2_bits_payload_r_type = io_in_2_bits_payload_r_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_voluntary = io_in_3_bits_payload_voluntary;
  assign arb_io_in_3_bits_payload_r_type = io_in_3_bits_payload_r_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_21;
  assign GEN_0_valid = GEN_22;
  assign GEN_0_bits_header_src = GEN_23;
  assign GEN_0_bits_header_dst = GEN_24;
  assign GEN_0_bits_payload_addr_beat = GEN_25;
  assign GEN_0_bits_payload_addr_block = GEN_26;
  assign GEN_0_bits_payload_client_xact_id = GEN_27;
  assign GEN_0_bits_payload_voluntary = GEN_28;
  assign GEN_0_bits_payload_r_type = GEN_29;
  assign GEN_0_bits_payload_data = GEN_30;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_voluntary : io_out_0_bits_payload_voluntary;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_r_type : io_out_0_bits_payload_r_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_5;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_6;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_7;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_voluntary : GEN_8;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_r_type : GEN_9;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_10;
  assign GEN_21 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_11;
  assign GEN_22 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_12;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_13;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_14;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_15;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_16;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_17;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_voluntary : GEN_18;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_r_type : GEN_19;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_20;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_p_type,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_p_type;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] GEN_7;
  wire [1:0] GEN_8;
  wire [25:0] GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [25:0] GEN_15;
  wire [1:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [1:0] GEN_19;
  wire [1:0] GEN_20;
  wire [25:0] GEN_21;
  wire [1:0] GEN_22;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [25:0] GEN_1_bits_payload_addr_block;
  wire [1:0] GEN_1_bits_payload_p_type;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [25:0] GEN_2_bits_payload_addr_block;
  wire [1:0] GEN_2_bits_payload_p_type;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [25:0] GEN_3_bits_payload_addr_block;
  wire [1:0] GEN_3_bits_payload_p_type;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [25:0] GEN_4_bits_payload_addr_block;
  wire [1:0] GEN_4_bits_payload_p_type;
  wire  T_964;
  reg [1:0] lastGrant;
  reg [31:0] GEN_0;
  wire [1:0] GEN_95;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire  T_978;
  wire  T_980;
  wire  T_982;
  wire  T_984;
  wire  T_986;
  wire  T_988;
  wire  T_992;
  wire  T_993;
  wire  T_994;
  wire  T_995;
  wire  T_996;
  wire  T_997;
  wire  T_998;
  wire  T_999;
  wire  T_1000;
  wire [1:0] GEN_96;
  wire [1:0] GEN_97;
  wire [1:0] GEN_98;
  wire [1:0] GEN_99;
  wire [1:0] GEN_100;
  wire [1:0] GEN_101;
  assign io_in_0_ready = T_997;
  assign io_in_1_ready = T_998;
  assign io_in_2_ready = T_999;
  assign io_in_3_ready = T_1000;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_block = GEN_3_bits_payload_addr_block;
  assign io_out_bits_payload_p_type = GEN_4_bits_payload_p_type;
  assign io_chosen = choice;
  assign choice = GEN_101;
  assign GEN_0_ready = GEN_17;
  assign GEN_0_valid = GEN_18;
  assign GEN_0_bits_header_src = GEN_19;
  assign GEN_0_bits_header_dst = GEN_20;
  assign GEN_0_bits_payload_addr_block = GEN_21;
  assign GEN_0_bits_payload_p_type = GEN_22;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_6 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_ready : GEN_5;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_valid : GEN_6;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_7;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_8;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_9;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_payload_p_type : GEN_10;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_ready : GEN_11;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_valid : GEN_12;
  assign GEN_19 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_14;
  assign GEN_21 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_15;
  assign GEN_22 = 2'h3 == io_chosen ? io_in_3_bits_payload_p_type : GEN_16;
  assign GEN_1_ready = GEN_17;
  assign GEN_1_valid = GEN_18;
  assign GEN_1_bits_header_src = GEN_19;
  assign GEN_1_bits_header_dst = GEN_20;
  assign GEN_1_bits_payload_addr_block = GEN_21;
  assign GEN_1_bits_payload_p_type = GEN_22;
  assign GEN_2_ready = GEN_17;
  assign GEN_2_valid = GEN_18;
  assign GEN_2_bits_header_src = GEN_19;
  assign GEN_2_bits_header_dst = GEN_20;
  assign GEN_2_bits_payload_addr_block = GEN_21;
  assign GEN_2_bits_payload_p_type = GEN_22;
  assign GEN_3_ready = GEN_17;
  assign GEN_3_valid = GEN_18;
  assign GEN_3_bits_header_src = GEN_19;
  assign GEN_3_bits_header_dst = GEN_20;
  assign GEN_3_bits_payload_addr_block = GEN_21;
  assign GEN_3_bits_payload_p_type = GEN_22;
  assign GEN_4_ready = GEN_17;
  assign GEN_4_valid = GEN_18;
  assign GEN_4_bits_header_src = GEN_19;
  assign GEN_4_bits_header_dst = GEN_20;
  assign GEN_4_bits_payload_addr_block = GEN_21;
  assign GEN_4_bits_payload_p_type = GEN_22;
  assign T_964 = io_out_ready & io_out_valid;
  assign GEN_95 = T_964 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_970 = validMask_1 | validMask_2;
  assign T_971 = T_970 | validMask_3;
  assign T_972 = T_971 | io_in_0_valid;
  assign T_973 = T_972 | io_in_1_valid;
  assign T_974 = T_973 | io_in_2_valid;
  assign T_978 = validMask_1 == 1'h0;
  assign T_980 = T_970 == 1'h0;
  assign T_982 = T_971 == 1'h0;
  assign T_984 = T_972 == 1'h0;
  assign T_986 = T_973 == 1'h0;
  assign T_988 = T_974 == 1'h0;
  assign T_992 = grantMask_1 | T_984;
  assign T_993 = T_978 & grantMask_2;
  assign T_994 = T_993 | T_986;
  assign T_995 = T_980 & grantMask_3;
  assign T_996 = T_995 | T_988;
  assign T_997 = T_982 & io_out_ready;
  assign T_998 = T_992 & io_out_ready;
  assign T_999 = T_994 & io_out_ready;
  assign T_1000 = T_996 & io_out_ready;
  assign GEN_96 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_97 = io_in_1_valid ? 2'h1 : GEN_96;
  assign GEN_98 = io_in_0_valid ? 2'h0 : GEN_97;
  assign GEN_99 = validMask_3 ? 2'h3 : GEN_98;
  assign GEN_100 = validMask_2 ? 2'h2 : GEN_99;
  assign GEN_101 = validMask_1 ? 2'h1 : GEN_100;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  lastGrant = GEN_0[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_964) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_p_type,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_p_type,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_p_type,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_p_type
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_p_type;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_p_type;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_p_type;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_p_type;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_p_type;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [25:0] GEN_0_bits_payload_addr_block;
  wire [1:0] GEN_0_bits_payload_p_type;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [25:0] GEN_5;
  wire [1:0] GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [25:0] GEN_17;
  wire [1:0] GEN_18;
  wire  T_1299;
  wire  T_1300;
  wire  T_1302;
  wire  T_1303;
  wire  T_1305;
  wire  T_1306;
  wire  T_1308;
  wire  T_1309;
  LockingRRArbiter_2 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(arb_io_in_0_bits_payload_p_type),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(arb_io_in_1_bits_payload_p_type),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(arb_io_in_2_bits_payload_p_type),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(arb_io_in_3_bits_payload_p_type),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_p_type(arb_io_out_bits_payload_p_type),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1300;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_1_valid = T_1303;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_2_valid = T_1306;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_3_valid = T_1309;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_p_type = io_in_0_bits_payload_p_type;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_p_type = io_in_1_bits_payload_p_type;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_p_type = io_in_2_bits_payload_p_type;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_p_type = io_in_3_bits_payload_p_type;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_13;
  assign GEN_0_valid = GEN_14;
  assign GEN_0_bits_header_src = GEN_15;
  assign GEN_0_bits_header_dst = GEN_16;
  assign GEN_0_bits_payload_addr_block = GEN_17;
  assign GEN_0_bits_payload_p_type = GEN_18;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_block : io_out_0_bits_payload_addr_block;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_p_type : io_out_0_bits_payload_p_type;
  assign GEN_7 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_8 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_9 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_10 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_block : GEN_5;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_p_type : GEN_6;
  assign GEN_13 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_7;
  assign GEN_14 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_8;
  assign GEN_15 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_9;
  assign GEN_16 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_10;
  assign GEN_17 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_block : GEN_11;
  assign GEN_18 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_p_type : GEN_12;
  assign T_1299 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1300 = arb_io_out_valid & T_1299;
  assign T_1302 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1303 = arb_io_out_valid & T_1302;
  assign T_1305 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1306 = arb_io_out_valid & T_1305;
  assign T_1308 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1309 = arb_io_out_valid & T_1308;
endmodule
module LockingRRArbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output  io_out_bits_payload_is_builtin_type,
  output [3:0] io_out_bits_payload_g_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [3:0] GEN_0_bits_payload_g_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire [3:0] GEN_17;
  wire [63:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [2:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire  GEN_26;
  wire [3:0] GEN_27;
  wire [63:0] GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire [2:0] GEN_33;
  wire [1:0] GEN_34;
  wire [2:0] GEN_35;
  wire  GEN_36;
  wire [3:0] GEN_37;
  wire [63:0] GEN_38;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [2:0] GEN_1_bits_payload_addr_beat;
  wire [1:0] GEN_1_bits_payload_client_xact_id;
  wire [2:0] GEN_1_bits_payload_manager_xact_id;
  wire  GEN_1_bits_payload_is_builtin_type;
  wire [3:0] GEN_1_bits_payload_g_type;
  wire [63:0] GEN_1_bits_payload_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [2:0] GEN_2_bits_payload_addr_beat;
  wire [1:0] GEN_2_bits_payload_client_xact_id;
  wire [2:0] GEN_2_bits_payload_manager_xact_id;
  wire  GEN_2_bits_payload_is_builtin_type;
  wire [3:0] GEN_2_bits_payload_g_type;
  wire [63:0] GEN_2_bits_payload_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [2:0] GEN_3_bits_payload_addr_beat;
  wire [1:0] GEN_3_bits_payload_client_xact_id;
  wire [2:0] GEN_3_bits_payload_manager_xact_id;
  wire  GEN_3_bits_payload_is_builtin_type;
  wire [3:0] GEN_3_bits_payload_g_type;
  wire [63:0] GEN_3_bits_payload_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [1:0] GEN_4_bits_header_src;
  wire [1:0] GEN_4_bits_header_dst;
  wire [2:0] GEN_4_bits_payload_addr_beat;
  wire [1:0] GEN_4_bits_payload_client_xact_id;
  wire [2:0] GEN_4_bits_payload_manager_xact_id;
  wire  GEN_4_bits_payload_is_builtin_type;
  wire [3:0] GEN_4_bits_payload_g_type;
  wire [63:0] GEN_4_bits_payload_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [1:0] GEN_5_bits_header_src;
  wire [1:0] GEN_5_bits_header_dst;
  wire [2:0] GEN_5_bits_payload_addr_beat;
  wire [1:0] GEN_5_bits_payload_client_xact_id;
  wire [2:0] GEN_5_bits_payload_manager_xact_id;
  wire  GEN_5_bits_payload_is_builtin_type;
  wire [3:0] GEN_5_bits_payload_g_type;
  wire [63:0] GEN_5_bits_payload_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [1:0] GEN_6_bits_header_src;
  wire [1:0] GEN_6_bits_header_dst;
  wire [2:0] GEN_6_bits_payload_addr_beat;
  wire [1:0] GEN_6_bits_payload_client_xact_id;
  wire [2:0] GEN_6_bits_payload_manager_xact_id;
  wire  GEN_6_bits_payload_is_builtin_type;
  wire [3:0] GEN_6_bits_payload_g_type;
  wire [63:0] GEN_6_bits_payload_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [1:0] GEN_7_bits_header_src;
  wire [1:0] GEN_7_bits_header_dst;
  wire [2:0] GEN_7_bits_payload_addr_beat;
  wire [1:0] GEN_7_bits_payload_client_xact_id;
  wire [2:0] GEN_7_bits_payload_manager_xact_id;
  wire  GEN_7_bits_payload_is_builtin_type;
  wire [3:0] GEN_7_bits_payload_g_type;
  wire [63:0] GEN_7_bits_payload_data;
  wire  GEN_8_ready;
  wire  GEN_8_valid;
  wire [1:0] GEN_8_bits_header_src;
  wire [1:0] GEN_8_bits_header_dst;
  wire [2:0] GEN_8_bits_payload_addr_beat;
  wire [1:0] GEN_8_bits_payload_client_xact_id;
  wire [2:0] GEN_8_bits_payload_manager_xact_id;
  wire  GEN_8_bits_payload_is_builtin_type;
  wire [3:0] GEN_8_bits_payload_g_type;
  wire [63:0] GEN_8_bits_payload_data;
  reg [2:0] T_1100;
  reg [31:0] GEN_1;
  reg [1:0] T_1102;
  reg [31:0] GEN_2;
  wire  T_1104;
  wire [2:0] T_1112_0;
  wire [3:0] GEN_0;
  wire  T_1114;
  wire  T_1115;
  wire  T_1116;
  wire  T_1118;
  wire  T_1119;
  wire [3:0] T_1123;
  wire [2:0] T_1124;
  wire [1:0] GEN_279;
  wire [2:0] GEN_280;
  wire [1:0] GEN_281;
  reg [1:0] lastGrant;
  reg [31:0] GEN_3;
  wire [1:0] GEN_282;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_1132;
  wire  T_1133;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire  T_1140;
  wire  T_1142;
  wire  T_1144;
  wire  T_1146;
  wire  T_1148;
  wire  T_1150;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1162;
  wire  T_1164;
  wire  T_1165;
  wire  T_1166;
  wire  T_1168;
  wire  T_1169;
  wire  T_1170;
  wire  T_1172;
  wire  T_1173;
  wire  T_1174;
  wire [1:0] GEN_283;
  wire [1:0] GEN_284;
  wire [1:0] GEN_285;
  wire [1:0] GEN_286;
  wire [1:0] GEN_287;
  wire [1:0] GEN_288;
  assign io_in_0_ready = T_1162;
  assign io_in_1_ready = T_1166;
  assign io_in_2_ready = T_1170;
  assign io_in_3_ready = T_1174;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_addr_beat = GEN_3_bits_payload_addr_beat;
  assign io_out_bits_payload_client_xact_id = GEN_4_bits_payload_client_xact_id;
  assign io_out_bits_payload_manager_xact_id = GEN_5_bits_payload_manager_xact_id;
  assign io_out_bits_payload_is_builtin_type = GEN_6_bits_payload_is_builtin_type;
  assign io_out_bits_payload_g_type = GEN_7_bits_payload_g_type;
  assign io_out_bits_payload_data = GEN_8_bits_payload_data;
  assign io_chosen = GEN_281;
  assign choice = GEN_288;
  assign GEN_0_ready = GEN_29;
  assign GEN_0_valid = GEN_30;
  assign GEN_0_bits_header_src = GEN_31;
  assign GEN_0_bits_header_dst = GEN_32;
  assign GEN_0_bits_payload_addr_beat = GEN_33;
  assign GEN_0_bits_payload_client_xact_id = GEN_34;
  assign GEN_0_bits_payload_manager_xact_id = GEN_35;
  assign GEN_0_bits_payload_is_builtin_type = GEN_36;
  assign GEN_0_bits_payload_g_type = GEN_37;
  assign GEN_0_bits_payload_data = GEN_38;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_ready : GEN_9;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_11;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_12;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_13;
  assign GEN_24 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_14;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_15;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_16;
  assign GEN_27 = 2'h2 == io_chosen ? io_in_2_bits_payload_g_type : GEN_17;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_18;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_ready : GEN_19;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_valid : GEN_20;
  assign GEN_31 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_21;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_22;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_23;
  assign GEN_34 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_24;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_25;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_26;
  assign GEN_37 = 2'h3 == io_chosen ? io_in_3_bits_payload_g_type : GEN_27;
  assign GEN_38 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_28;
  assign GEN_1_ready = GEN_29;
  assign GEN_1_valid = GEN_30;
  assign GEN_1_bits_header_src = GEN_31;
  assign GEN_1_bits_header_dst = GEN_32;
  assign GEN_1_bits_payload_addr_beat = GEN_33;
  assign GEN_1_bits_payload_client_xact_id = GEN_34;
  assign GEN_1_bits_payload_manager_xact_id = GEN_35;
  assign GEN_1_bits_payload_is_builtin_type = GEN_36;
  assign GEN_1_bits_payload_g_type = GEN_37;
  assign GEN_1_bits_payload_data = GEN_38;
  assign GEN_2_ready = GEN_29;
  assign GEN_2_valid = GEN_30;
  assign GEN_2_bits_header_src = GEN_31;
  assign GEN_2_bits_header_dst = GEN_32;
  assign GEN_2_bits_payload_addr_beat = GEN_33;
  assign GEN_2_bits_payload_client_xact_id = GEN_34;
  assign GEN_2_bits_payload_manager_xact_id = GEN_35;
  assign GEN_2_bits_payload_is_builtin_type = GEN_36;
  assign GEN_2_bits_payload_g_type = GEN_37;
  assign GEN_2_bits_payload_data = GEN_38;
  assign GEN_3_ready = GEN_29;
  assign GEN_3_valid = GEN_30;
  assign GEN_3_bits_header_src = GEN_31;
  assign GEN_3_bits_header_dst = GEN_32;
  assign GEN_3_bits_payload_addr_beat = GEN_33;
  assign GEN_3_bits_payload_client_xact_id = GEN_34;
  assign GEN_3_bits_payload_manager_xact_id = GEN_35;
  assign GEN_3_bits_payload_is_builtin_type = GEN_36;
  assign GEN_3_bits_payload_g_type = GEN_37;
  assign GEN_3_bits_payload_data = GEN_38;
  assign GEN_4_ready = GEN_29;
  assign GEN_4_valid = GEN_30;
  assign GEN_4_bits_header_src = GEN_31;
  assign GEN_4_bits_header_dst = GEN_32;
  assign GEN_4_bits_payload_addr_beat = GEN_33;
  assign GEN_4_bits_payload_client_xact_id = GEN_34;
  assign GEN_4_bits_payload_manager_xact_id = GEN_35;
  assign GEN_4_bits_payload_is_builtin_type = GEN_36;
  assign GEN_4_bits_payload_g_type = GEN_37;
  assign GEN_4_bits_payload_data = GEN_38;
  assign GEN_5_ready = GEN_29;
  assign GEN_5_valid = GEN_30;
  assign GEN_5_bits_header_src = GEN_31;
  assign GEN_5_bits_header_dst = GEN_32;
  assign GEN_5_bits_payload_addr_beat = GEN_33;
  assign GEN_5_bits_payload_client_xact_id = GEN_34;
  assign GEN_5_bits_payload_manager_xact_id = GEN_35;
  assign GEN_5_bits_payload_is_builtin_type = GEN_36;
  assign GEN_5_bits_payload_g_type = GEN_37;
  assign GEN_5_bits_payload_data = GEN_38;
  assign GEN_6_ready = GEN_29;
  assign GEN_6_valid = GEN_30;
  assign GEN_6_bits_header_src = GEN_31;
  assign GEN_6_bits_header_dst = GEN_32;
  assign GEN_6_bits_payload_addr_beat = GEN_33;
  assign GEN_6_bits_payload_client_xact_id = GEN_34;
  assign GEN_6_bits_payload_manager_xact_id = GEN_35;
  assign GEN_6_bits_payload_is_builtin_type = GEN_36;
  assign GEN_6_bits_payload_g_type = GEN_37;
  assign GEN_6_bits_payload_data = GEN_38;
  assign GEN_7_ready = GEN_29;
  assign GEN_7_valid = GEN_30;
  assign GEN_7_bits_header_src = GEN_31;
  assign GEN_7_bits_header_dst = GEN_32;
  assign GEN_7_bits_payload_addr_beat = GEN_33;
  assign GEN_7_bits_payload_client_xact_id = GEN_34;
  assign GEN_7_bits_payload_manager_xact_id = GEN_35;
  assign GEN_7_bits_payload_is_builtin_type = GEN_36;
  assign GEN_7_bits_payload_g_type = GEN_37;
  assign GEN_7_bits_payload_data = GEN_38;
  assign GEN_8_ready = GEN_29;
  assign GEN_8_valid = GEN_30;
  assign GEN_8_bits_header_src = GEN_31;
  assign GEN_8_bits_header_dst = GEN_32;
  assign GEN_8_bits_payload_addr_beat = GEN_33;
  assign GEN_8_bits_payload_client_xact_id = GEN_34;
  assign GEN_8_bits_payload_manager_xact_id = GEN_35;
  assign GEN_8_bits_payload_is_builtin_type = GEN_36;
  assign GEN_8_bits_payload_g_type = GEN_37;
  assign GEN_8_bits_payload_data = GEN_38;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1112_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1112_0};
  assign T_1114 = io_out_bits_payload_g_type == GEN_0;
  assign T_1115 = io_out_bits_payload_g_type == 4'h0;
  assign T_1116 = io_out_bits_payload_is_builtin_type ? T_1114 : T_1115;
  assign T_1118 = io_out_ready & io_out_valid;
  assign T_1119 = T_1118 & T_1116;
  assign T_1123 = T_1100 + 3'h1;
  assign T_1124 = T_1123[2:0];
  assign GEN_279 = T_1119 ? io_chosen : T_1102;
  assign GEN_280 = T_1119 ? T_1124 : T_1100;
  assign GEN_281 = T_1104 ? T_1102 : choice;
  assign GEN_282 = T_1118 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_1132 = validMask_1 | validMask_2;
  assign T_1133 = T_1132 | validMask_3;
  assign T_1134 = T_1133 | io_in_0_valid;
  assign T_1135 = T_1134 | io_in_1_valid;
  assign T_1136 = T_1135 | io_in_2_valid;
  assign T_1140 = validMask_1 == 1'h0;
  assign T_1142 = T_1132 == 1'h0;
  assign T_1144 = T_1133 == 1'h0;
  assign T_1146 = T_1134 == 1'h0;
  assign T_1148 = T_1135 == 1'h0;
  assign T_1150 = T_1136 == 1'h0;
  assign T_1154 = grantMask_1 | T_1146;
  assign T_1155 = T_1140 & grantMask_2;
  assign T_1156 = T_1155 | T_1148;
  assign T_1157 = T_1142 & grantMask_3;
  assign T_1158 = T_1157 | T_1150;
  assign T_1160 = T_1102 == 2'h0;
  assign T_1161 = T_1104 ? T_1160 : T_1144;
  assign T_1162 = T_1161 & io_out_ready;
  assign T_1164 = T_1102 == 2'h1;
  assign T_1165 = T_1104 ? T_1164 : T_1154;
  assign T_1166 = T_1165 & io_out_ready;
  assign T_1168 = T_1102 == 2'h2;
  assign T_1169 = T_1104 ? T_1168 : T_1156;
  assign T_1170 = T_1169 & io_out_ready;
  assign T_1172 = T_1102 == 2'h3;
  assign T_1173 = T_1104 ? T_1172 : T_1158;
  assign T_1174 = T_1173 & io_out_ready;
  assign GEN_283 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_284 = io_in_1_valid ? 2'h1 : GEN_283;
  assign GEN_285 = io_in_0_valid ? 2'h0 : GEN_284;
  assign GEN_286 = validMask_3 ? 2'h3 : GEN_285;
  assign GEN_287 = validMask_2 ? 2'h2 : GEN_286;
  assign GEN_288 = validMask_1 ? 2'h1 : GEN_287;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1100 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_1102 = GEN_2[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1119) begin
        T_1100 <= T_1124;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1119) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1118) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  output  io_out_0_bits_payload_is_builtin_type,
  output [3:0] io_out_0_bits_payload_g_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  output  io_out_1_bits_payload_is_builtin_type,
  output [3:0] io_out_1_bits_payload_g_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  output  io_out_2_bits_payload_is_builtin_type,
  output [3:0] io_out_2_bits_payload_g_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_manager_xact_id,
  output  io_out_3_bits_payload_is_builtin_type,
  output [3:0] io_out_3_bits_payload_g_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_0_bits_payload_g_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_1_bits_payload_g_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_2_bits_payload_g_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_3_bits_payload_g_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [3:0] arb_io_out_bits_payload_g_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_addr_beat;
  wire [1:0] GEN_0_bits_payload_client_xact_id;
  wire [2:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_0_bits_payload_is_builtin_type;
  wire [3:0] GEN_0_bits_payload_g_type;
  wire [63:0] GEN_0_bits_payload_data;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [2:0] GEN_5;
  wire [1:0] GEN_6;
  wire [2:0] GEN_7;
  wire  GEN_8;
  wire [3:0] GEN_9;
  wire [63:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire [1:0] GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  wire [3:0] GEN_19;
  wire [63:0] GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire [1:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [3:0] GEN_29;
  wire [63:0] GEN_30;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_3 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(arb_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(arb_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(arb_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(arb_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_g_type(arb_io_out_bits_payload_g_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_g_type = io_in_1_bits_payload_g_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_g_type = io_in_2_bits_payload_g_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_g_type = io_in_3_bits_payload_g_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_21;
  assign GEN_0_valid = GEN_22;
  assign GEN_0_bits_header_src = GEN_23;
  assign GEN_0_bits_header_dst = GEN_24;
  assign GEN_0_bits_payload_addr_beat = GEN_25;
  assign GEN_0_bits_payload_client_xact_id = GEN_26;
  assign GEN_0_bits_payload_manager_xact_id = GEN_27;
  assign GEN_0_bits_payload_is_builtin_type = GEN_28;
  assign GEN_0_bits_payload_g_type = GEN_29;
  assign GEN_0_bits_payload_data = GEN_30;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_addr_beat : io_out_0_bits_payload_addr_beat;
  assign GEN_6 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_client_xact_id : io_out_0_bits_payload_client_xact_id;
  assign GEN_7 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_manager_xact_id : io_out_0_bits_payload_manager_xact_id;
  assign GEN_8 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_is_builtin_type : io_out_0_bits_payload_is_builtin_type;
  assign GEN_9 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_g_type : io_out_0_bits_payload_g_type;
  assign GEN_10 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_data : io_out_0_bits_payload_data;
  assign GEN_11 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_12 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_13 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_14 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_15 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_addr_beat : GEN_5;
  assign GEN_16 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_client_xact_id : GEN_6;
  assign GEN_17 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_manager_xact_id : GEN_7;
  assign GEN_18 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_is_builtin_type : GEN_8;
  assign GEN_19 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_g_type : GEN_9;
  assign GEN_20 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_data : GEN_10;
  assign GEN_21 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_11;
  assign GEN_22 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_12;
  assign GEN_23 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_13;
  assign GEN_24 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_14;
  assign GEN_25 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_addr_beat : GEN_15;
  assign GEN_26 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_client_xact_id : GEN_16;
  assign GEN_27 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_manager_xact_id : GEN_17;
  assign GEN_28 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_is_builtin_type : GEN_18;
  assign GEN_29 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_g_type : GEN_19;
  assign GEN_30 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_data : GEN_20;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_4;
  wire  GEN_5;
  wire [1:0] GEN_6;
  wire [1:0] GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [2:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_18;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [1:0] GEN_1_bits_header_src;
  wire [1:0] GEN_1_bits_header_dst;
  wire [2:0] GEN_1_bits_payload_manager_xact_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [1:0] GEN_2_bits_header_src;
  wire [1:0] GEN_2_bits_header_dst;
  wire [2:0] GEN_2_bits_payload_manager_xact_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [1:0] GEN_3_bits_header_src;
  wire [1:0] GEN_3_bits_header_dst;
  wire [2:0] GEN_3_bits_payload_manager_xact_id;
  wire  T_930;
  reg [1:0] lastGrant;
  reg [31:0] GEN_0;
  wire [1:0] GEN_64;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_944;
  wire  T_946;
  wire  T_948;
  wire  T_950;
  wire  T_952;
  wire  T_954;
  wire  T_958;
  wire  T_959;
  wire  T_960;
  wire  T_961;
  wire  T_962;
  wire  T_963;
  wire  T_964;
  wire  T_965;
  wire  T_966;
  wire [1:0] GEN_65;
  wire [1:0] GEN_66;
  wire [1:0] GEN_67;
  wire [1:0] GEN_68;
  wire [1:0] GEN_69;
  wire [1:0] GEN_70;
  assign io_in_0_ready = T_963;
  assign io_in_1_ready = T_964;
  assign io_in_2_ready = T_965;
  assign io_in_3_ready = T_966;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_header_src = GEN_1_bits_header_src;
  assign io_out_bits_header_dst = GEN_2_bits_header_dst;
  assign io_out_bits_payload_manager_xact_id = GEN_3_bits_payload_manager_xact_id;
  assign io_chosen = choice;
  assign choice = GEN_70;
  assign GEN_0_ready = GEN_14;
  assign GEN_0_valid = GEN_15;
  assign GEN_0_bits_header_src = GEN_16;
  assign GEN_0_bits_header_dst = GEN_17;
  assign GEN_0_bits_payload_manager_xact_id = GEN_18;
  assign GEN_4 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_ready : GEN_4;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_6;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_7;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_8;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_ready : GEN_9;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_16 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_11;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_12;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_13;
  assign GEN_1_ready = GEN_14;
  assign GEN_1_valid = GEN_15;
  assign GEN_1_bits_header_src = GEN_16;
  assign GEN_1_bits_header_dst = GEN_17;
  assign GEN_1_bits_payload_manager_xact_id = GEN_18;
  assign GEN_2_ready = GEN_14;
  assign GEN_2_valid = GEN_15;
  assign GEN_2_bits_header_src = GEN_16;
  assign GEN_2_bits_header_dst = GEN_17;
  assign GEN_2_bits_payload_manager_xact_id = GEN_18;
  assign GEN_3_ready = GEN_14;
  assign GEN_3_valid = GEN_15;
  assign GEN_3_bits_header_src = GEN_16;
  assign GEN_3_bits_header_dst = GEN_17;
  assign GEN_3_bits_payload_manager_xact_id = GEN_18;
  assign T_930 = io_out_ready & io_out_valid;
  assign GEN_64 = T_930 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_936 = validMask_1 | validMask_2;
  assign T_937 = T_936 | validMask_3;
  assign T_938 = T_937 | io_in_0_valid;
  assign T_939 = T_938 | io_in_1_valid;
  assign T_940 = T_939 | io_in_2_valid;
  assign T_944 = validMask_1 == 1'h0;
  assign T_946 = T_936 == 1'h0;
  assign T_948 = T_937 == 1'h0;
  assign T_950 = T_938 == 1'h0;
  assign T_952 = T_939 == 1'h0;
  assign T_954 = T_940 == 1'h0;
  assign T_958 = grantMask_1 | T_950;
  assign T_959 = T_944 & grantMask_2;
  assign T_960 = T_959 | T_952;
  assign T_961 = T_946 & grantMask_3;
  assign T_962 = T_961 | T_954;
  assign T_963 = T_948 & io_out_ready;
  assign T_964 = T_958 & io_out_ready;
  assign T_965 = T_960 & io_out_ready;
  assign T_966 = T_962 & io_out_ready;
  assign GEN_65 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_66 = io_in_1_valid ? 2'h1 : GEN_65;
  assign GEN_67 = io_in_0_valid ? 2'h0 : GEN_66;
  assign GEN_68 = validMask_3 ? 2'h3 : GEN_67;
  assign GEN_69 = validMask_2 ? 2'h2 : GEN_68;
  assign GEN_70 = validMask_1 ? 2'h1 : GEN_69;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  lastGrant = GEN_0[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_930) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_manager_xact_id
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire [1:0] arb_io_chosen;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [1:0] GEN_0_bits_header_src;
  wire [1:0] GEN_0_bits_header_dst;
  wire [2:0] GEN_0_bits_payload_manager_xact_id;
  wire  GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [1:0] GEN_4;
  wire [2:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [2:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [2:0] GEN_15;
  wire  T_1253;
  wire  T_1254;
  wire  T_1256;
  wire  T_1257;
  wire  T_1259;
  wire  T_1260;
  wire  T_1262;
  wire  T_1263;
  LockingRRArbiter_4 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1254;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_valid = T_1257;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_valid = T_1260;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_valid = T_1263;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_out_ready = GEN_0_ready;
  assign GEN_0_ready = GEN_11;
  assign GEN_0_valid = GEN_12;
  assign GEN_0_bits_header_src = GEN_13;
  assign GEN_0_bits_header_dst = GEN_14;
  assign GEN_0_bits_payload_manager_xact_id = GEN_15;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_valid : io_out_0_valid;
  assign GEN_3 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_src : io_out_0_bits_header_src;
  assign GEN_4 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_header_dst : io_out_0_bits_header_dst;
  assign GEN_5 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_bits_payload_manager_xact_id : io_out_0_bits_payload_manager_xact_id;
  assign GEN_6 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_valid : GEN_2;
  assign GEN_8 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_src : GEN_3;
  assign GEN_9 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_header_dst : GEN_4;
  assign GEN_10 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_bits_payload_manager_xact_id : GEN_5;
  assign GEN_11 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_6;
  assign GEN_12 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_valid : GEN_7;
  assign GEN_13 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_src : GEN_8;
  assign GEN_14 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_header_dst : GEN_9;
  assign GEN_15 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_bits_payload_manager_xact_id : GEN_10;
  assign T_1253 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1254 = arb_io_out_valid & T_1253;
  assign T_1256 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1257 = arb_io_out_valid & T_1256;
  assign T_1259 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1260 = arb_io_out_valid & T_1259;
  assign T_1262 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1263 = arb_io_out_valid & T_1262;
endmodule
module PortedTileLinkCrossbar(
  input   clk,
  input   reset,
  output  io_clients_cached_0_acquire_ready,
  input   io_clients_cached_0_acquire_valid,
  input  [25:0] io_clients_cached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_cached_0_acquire_bits_addr_beat,
  input   io_clients_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_cached_0_acquire_bits_a_type,
  input  [10:0] io_clients_cached_0_acquire_bits_union,
  input  [63:0] io_clients_cached_0_acquire_bits_data,
  input   io_clients_cached_0_probe_ready,
  output  io_clients_cached_0_probe_valid,
  output [25:0] io_clients_cached_0_probe_bits_addr_block,
  output [1:0] io_clients_cached_0_probe_bits_p_type,
  output  io_clients_cached_0_release_ready,
  input   io_clients_cached_0_release_valid,
  input  [2:0] io_clients_cached_0_release_bits_addr_beat,
  input  [25:0] io_clients_cached_0_release_bits_addr_block,
  input  [1:0] io_clients_cached_0_release_bits_client_xact_id,
  input   io_clients_cached_0_release_bits_voluntary,
  input  [2:0] io_clients_cached_0_release_bits_r_type,
  input  [63:0] io_clients_cached_0_release_bits_data,
  input   io_clients_cached_0_grant_ready,
  output  io_clients_cached_0_grant_valid,
  output [2:0] io_clients_cached_0_grant_bits_addr_beat,
  output [1:0] io_clients_cached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_cached_0_grant_bits_manager_xact_id,
  output  io_clients_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_cached_0_grant_bits_g_type,
  output [63:0] io_clients_cached_0_grant_bits_data,
  output  io_clients_cached_0_grant_bits_manager_id,
  output  io_clients_cached_0_finish_ready,
  input   io_clients_cached_0_finish_valid,
  input  [2:0] io_clients_cached_0_finish_bits_manager_xact_id,
  input   io_clients_cached_0_finish_bits_manager_id,
  output  io_clients_uncached_0_acquire_ready,
  input   io_clients_uncached_0_acquire_valid,
  input  [25:0] io_clients_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_0_acquire_bits_addr_beat,
  input   io_clients_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_0_acquire_bits_a_type,
  input  [10:0] io_clients_uncached_0_acquire_bits_union,
  input  [63:0] io_clients_uncached_0_acquire_bits_data,
  input   io_clients_uncached_0_grant_ready,
  output  io_clients_uncached_0_grant_valid,
  output [2:0] io_clients_uncached_0_grant_bits_addr_beat,
  output [1:0] io_clients_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_uncached_0_grant_bits_manager_xact_id,
  output  io_clients_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_0_grant_bits_g_type,
  output [63:0] io_clients_uncached_0_grant_bits_data,
  input   io_managers_0_acquire_ready,
  output  io_managers_0_acquire_valid,
  output [25:0] io_managers_0_acquire_bits_addr_block,
  output [1:0] io_managers_0_acquire_bits_client_xact_id,
  output [2:0] io_managers_0_acquire_bits_addr_beat,
  output  io_managers_0_acquire_bits_is_builtin_type,
  output [2:0] io_managers_0_acquire_bits_a_type,
  output [10:0] io_managers_0_acquire_bits_union,
  output [63:0] io_managers_0_acquire_bits_data,
  output  io_managers_0_acquire_bits_client_id,
  output  io_managers_0_grant_ready,
  input   io_managers_0_grant_valid,
  input  [2:0] io_managers_0_grant_bits_addr_beat,
  input  [1:0] io_managers_0_grant_bits_client_xact_id,
  input  [2:0] io_managers_0_grant_bits_manager_xact_id,
  input   io_managers_0_grant_bits_is_builtin_type,
  input  [3:0] io_managers_0_grant_bits_g_type,
  input  [63:0] io_managers_0_grant_bits_data,
  input   io_managers_0_grant_bits_client_id,
  input   io_managers_0_finish_ready,
  output  io_managers_0_finish_valid,
  output [2:0] io_managers_0_finish_bits_manager_xact_id,
  output  io_managers_0_probe_ready,
  input   io_managers_0_probe_valid,
  input  [25:0] io_managers_0_probe_bits_addr_block,
  input  [1:0] io_managers_0_probe_bits_p_type,
  input   io_managers_0_probe_bits_client_id,
  input   io_managers_0_release_ready,
  output  io_managers_0_release_valid,
  output [2:0] io_managers_0_release_bits_addr_beat,
  output [25:0] io_managers_0_release_bits_addr_block,
  output [1:0] io_managers_0_release_bits_client_xact_id,
  output  io_managers_0_release_bits_voluntary,
  output [2:0] io_managers_0_release_bits_r_type,
  output [63:0] io_managers_0_release_bits_data,
  output  io_managers_0_release_bits_client_id,
  input   io_managers_1_acquire_ready,
  output  io_managers_1_acquire_valid,
  output [25:0] io_managers_1_acquire_bits_addr_block,
  output [1:0] io_managers_1_acquire_bits_client_xact_id,
  output [2:0] io_managers_1_acquire_bits_addr_beat,
  output  io_managers_1_acquire_bits_is_builtin_type,
  output [2:0] io_managers_1_acquire_bits_a_type,
  output [10:0] io_managers_1_acquire_bits_union,
  output [63:0] io_managers_1_acquire_bits_data,
  output  io_managers_1_acquire_bits_client_id,
  output  io_managers_1_grant_ready,
  input   io_managers_1_grant_valid,
  input  [2:0] io_managers_1_grant_bits_addr_beat,
  input  [1:0] io_managers_1_grant_bits_client_xact_id,
  input  [2:0] io_managers_1_grant_bits_manager_xact_id,
  input   io_managers_1_grant_bits_is_builtin_type,
  input  [3:0] io_managers_1_grant_bits_g_type,
  input  [63:0] io_managers_1_grant_bits_data,
  input   io_managers_1_grant_bits_client_id,
  input   io_managers_1_finish_ready,
  output  io_managers_1_finish_valid,
  output [2:0] io_managers_1_finish_bits_manager_xact_id,
  output  io_managers_1_probe_ready,
  input   io_managers_1_probe_valid,
  input  [25:0] io_managers_1_probe_bits_addr_block,
  input  [1:0] io_managers_1_probe_bits_p_type,
  input   io_managers_1_probe_bits_client_id,
  input   io_managers_1_release_ready,
  output  io_managers_1_release_valid,
  output [2:0] io_managers_1_release_bits_addr_beat,
  output [25:0] io_managers_1_release_bits_addr_block,
  output [1:0] io_managers_1_release_bits_client_xact_id,
  output  io_managers_1_release_bits_voluntary,
  output [2:0] io_managers_1_release_bits_r_type,
  output [63:0] io_managers_1_release_bits_data,
  output  io_managers_1_release_bits_client_id
);
  wire  TileLinkEnqueuer_4_clk;
  wire  TileLinkEnqueuer_4_reset;
  wire  TileLinkEnqueuer_4_io_client_acquire_ready;
  wire  TileLinkEnqueuer_4_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_grant_ready;
  wire  TileLinkEnqueuer_4_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_finish_ready;
  wire  TileLinkEnqueuer_4_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_probe_ready;
  wire  TileLinkEnqueuer_4_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_client_release_ready;
  wire  TileLinkEnqueuer_4_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_4_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_grant_ready;
  wire  TileLinkEnqueuer_4_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_finish_ready;
  wire  TileLinkEnqueuer_4_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_probe_ready;
  wire  TileLinkEnqueuer_4_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_manager_release_ready;
  wire  TileLinkEnqueuer_4_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_clk;
  wire  ClientTileLinkNetworkPort_1_reset;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [10:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire  ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_release_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_clk;
  wire  TileLinkEnqueuer_1_1_reset;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_client_release_ready;
  wire  TileLinkEnqueuer_1_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_clk;
  wire  ClientUncachedTileLinkNetworkPort_1_reset;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_clk;
  wire  ManagerTileLinkNetworkPort_2_reset;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_clk;
  wire  TileLinkEnqueuer_2_1_reset;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_client_release_ready;
  wire  TileLinkEnqueuer_2_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_clk;
  wire  ManagerTileLinkNetworkPort_1_1_reset;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type;
  wire [10:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_clk;
  wire  TileLinkEnqueuer_3_1_reset;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_client_release_ready;
  wire  TileLinkEnqueuer_3_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  wire [10:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  wire  acqNet_clk;
  wire  acqNet_reset;
  wire  acqNet_io_in_0_ready;
  wire  acqNet_io_in_0_valid;
  wire [1:0] acqNet_io_in_0_bits_header_src;
  wire [1:0] acqNet_io_in_0_bits_header_dst;
  wire [25:0] acqNet_io_in_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_0_bits_payload_addr_beat;
  wire  acqNet_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_0_bits_payload_a_type;
  wire [10:0] acqNet_io_in_0_bits_payload_union;
  wire [63:0] acqNet_io_in_0_bits_payload_data;
  wire  acqNet_io_in_1_ready;
  wire  acqNet_io_in_1_valid;
  wire [1:0] acqNet_io_in_1_bits_header_src;
  wire [1:0] acqNet_io_in_1_bits_header_dst;
  wire [25:0] acqNet_io_in_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_1_bits_payload_addr_beat;
  wire  acqNet_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_1_bits_payload_a_type;
  wire [10:0] acqNet_io_in_1_bits_payload_union;
  wire [63:0] acqNet_io_in_1_bits_payload_data;
  wire  acqNet_io_in_2_ready;
  wire  acqNet_io_in_2_valid;
  wire [1:0] acqNet_io_in_2_bits_header_src;
  wire [1:0] acqNet_io_in_2_bits_header_dst;
  wire [25:0] acqNet_io_in_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_2_bits_payload_addr_beat;
  wire  acqNet_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_2_bits_payload_a_type;
  wire [10:0] acqNet_io_in_2_bits_payload_union;
  wire [63:0] acqNet_io_in_2_bits_payload_data;
  wire  acqNet_io_in_3_ready;
  wire  acqNet_io_in_3_valid;
  wire [1:0] acqNet_io_in_3_bits_header_src;
  wire [1:0] acqNet_io_in_3_bits_header_dst;
  wire [25:0] acqNet_io_in_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_3_bits_payload_addr_beat;
  wire  acqNet_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_3_bits_payload_a_type;
  wire [10:0] acqNet_io_in_3_bits_payload_union;
  wire [63:0] acqNet_io_in_3_bits_payload_data;
  wire  acqNet_io_out_0_ready;
  wire  acqNet_io_out_0_valid;
  wire [1:0] acqNet_io_out_0_bits_header_src;
  wire [1:0] acqNet_io_out_0_bits_header_dst;
  wire [25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire  acqNet_io_out_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_0_bits_payload_a_type;
  wire [10:0] acqNet_io_out_0_bits_payload_union;
  wire [63:0] acqNet_io_out_0_bits_payload_data;
  wire  acqNet_io_out_1_ready;
  wire  acqNet_io_out_1_valid;
  wire [1:0] acqNet_io_out_1_bits_header_src;
  wire [1:0] acqNet_io_out_1_bits_header_dst;
  wire [25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire  acqNet_io_out_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_1_bits_payload_a_type;
  wire [10:0] acqNet_io_out_1_bits_payload_union;
  wire [63:0] acqNet_io_out_1_bits_payload_data;
  wire  acqNet_io_out_2_ready;
  wire  acqNet_io_out_2_valid;
  wire [1:0] acqNet_io_out_2_bits_header_src;
  wire [1:0] acqNet_io_out_2_bits_header_dst;
  wire [25:0] acqNet_io_out_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_2_bits_payload_addr_beat;
  wire  acqNet_io_out_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_2_bits_payload_a_type;
  wire [10:0] acqNet_io_out_2_bits_payload_union;
  wire [63:0] acqNet_io_out_2_bits_payload_data;
  wire  acqNet_io_out_3_ready;
  wire  acqNet_io_out_3_valid;
  wire [1:0] acqNet_io_out_3_bits_header_src;
  wire [1:0] acqNet_io_out_3_bits_header_dst;
  wire [25:0] acqNet_io_out_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_3_bits_payload_addr_beat;
  wire  acqNet_io_out_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_3_bits_payload_a_type;
  wire [10:0] acqNet_io_out_3_bits_payload_union;
  wire [63:0] acqNet_io_out_3_bits_payload_data;
  wire  relNet_clk;
  wire  relNet_reset;
  wire  relNet_io_in_0_ready;
  wire  relNet_io_in_0_valid;
  wire [1:0] relNet_io_in_0_bits_header_src;
  wire [1:0] relNet_io_in_0_bits_header_dst;
  wire [2:0] relNet_io_in_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_0_bits_payload_addr_block;
  wire [1:0] relNet_io_in_0_bits_payload_client_xact_id;
  wire  relNet_io_in_0_bits_payload_voluntary;
  wire [2:0] relNet_io_in_0_bits_payload_r_type;
  wire [63:0] relNet_io_in_0_bits_payload_data;
  wire  relNet_io_in_1_ready;
  wire  relNet_io_in_1_valid;
  wire [1:0] relNet_io_in_1_bits_header_src;
  wire [1:0] relNet_io_in_1_bits_header_dst;
  wire [2:0] relNet_io_in_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_1_bits_payload_addr_block;
  wire [1:0] relNet_io_in_1_bits_payload_client_xact_id;
  wire  relNet_io_in_1_bits_payload_voluntary;
  wire [2:0] relNet_io_in_1_bits_payload_r_type;
  wire [63:0] relNet_io_in_1_bits_payload_data;
  wire  relNet_io_in_2_ready;
  wire  relNet_io_in_2_valid;
  wire [1:0] relNet_io_in_2_bits_header_src;
  wire [1:0] relNet_io_in_2_bits_header_dst;
  wire [2:0] relNet_io_in_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_2_bits_payload_addr_block;
  wire [1:0] relNet_io_in_2_bits_payload_client_xact_id;
  wire  relNet_io_in_2_bits_payload_voluntary;
  wire [2:0] relNet_io_in_2_bits_payload_r_type;
  wire [63:0] relNet_io_in_2_bits_payload_data;
  wire  relNet_io_in_3_ready;
  wire  relNet_io_in_3_valid;
  wire [1:0] relNet_io_in_3_bits_header_src;
  wire [1:0] relNet_io_in_3_bits_header_dst;
  wire [2:0] relNet_io_in_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_3_bits_payload_addr_block;
  wire [1:0] relNet_io_in_3_bits_payload_client_xact_id;
  wire  relNet_io_in_3_bits_payload_voluntary;
  wire [2:0] relNet_io_in_3_bits_payload_r_type;
  wire [63:0] relNet_io_in_3_bits_payload_data;
  wire  relNet_io_out_0_ready;
  wire  relNet_io_out_0_valid;
  wire [1:0] relNet_io_out_0_bits_header_src;
  wire [1:0] relNet_io_out_0_bits_header_dst;
  wire [2:0] relNet_io_out_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_0_bits_payload_addr_block;
  wire [1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire  relNet_io_out_0_bits_payload_voluntary;
  wire [2:0] relNet_io_out_0_bits_payload_r_type;
  wire [63:0] relNet_io_out_0_bits_payload_data;
  wire  relNet_io_out_1_ready;
  wire  relNet_io_out_1_valid;
  wire [1:0] relNet_io_out_1_bits_header_src;
  wire [1:0] relNet_io_out_1_bits_header_dst;
  wire [2:0] relNet_io_out_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_1_bits_payload_addr_block;
  wire [1:0] relNet_io_out_1_bits_payload_client_xact_id;
  wire  relNet_io_out_1_bits_payload_voluntary;
  wire [2:0] relNet_io_out_1_bits_payload_r_type;
  wire [63:0] relNet_io_out_1_bits_payload_data;
  wire  relNet_io_out_2_ready;
  wire  relNet_io_out_2_valid;
  wire [1:0] relNet_io_out_2_bits_header_src;
  wire [1:0] relNet_io_out_2_bits_header_dst;
  wire [2:0] relNet_io_out_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_2_bits_payload_addr_block;
  wire [1:0] relNet_io_out_2_bits_payload_client_xact_id;
  wire  relNet_io_out_2_bits_payload_voluntary;
  wire [2:0] relNet_io_out_2_bits_payload_r_type;
  wire [63:0] relNet_io_out_2_bits_payload_data;
  wire  relNet_io_out_3_ready;
  wire  relNet_io_out_3_valid;
  wire [1:0] relNet_io_out_3_bits_header_src;
  wire [1:0] relNet_io_out_3_bits_header_dst;
  wire [2:0] relNet_io_out_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_3_bits_payload_addr_block;
  wire [1:0] relNet_io_out_3_bits_payload_client_xact_id;
  wire  relNet_io_out_3_bits_payload_voluntary;
  wire [2:0] relNet_io_out_3_bits_payload_r_type;
  wire [63:0] relNet_io_out_3_bits_payload_data;
  wire  prbNet_clk;
  wire  prbNet_reset;
  wire  prbNet_io_in_0_ready;
  wire  prbNet_io_in_0_valid;
  wire [1:0] prbNet_io_in_0_bits_header_src;
  wire [1:0] prbNet_io_in_0_bits_header_dst;
  wire [25:0] prbNet_io_in_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_0_bits_payload_p_type;
  wire  prbNet_io_in_1_ready;
  wire  prbNet_io_in_1_valid;
  wire [1:0] prbNet_io_in_1_bits_header_src;
  wire [1:0] prbNet_io_in_1_bits_header_dst;
  wire [25:0] prbNet_io_in_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_1_bits_payload_p_type;
  wire  prbNet_io_in_2_ready;
  wire  prbNet_io_in_2_valid;
  wire [1:0] prbNet_io_in_2_bits_header_src;
  wire [1:0] prbNet_io_in_2_bits_header_dst;
  wire [25:0] prbNet_io_in_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_2_bits_payload_p_type;
  wire  prbNet_io_in_3_ready;
  wire  prbNet_io_in_3_valid;
  wire [1:0] prbNet_io_in_3_bits_header_src;
  wire [1:0] prbNet_io_in_3_bits_header_dst;
  wire [25:0] prbNet_io_in_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_3_bits_payload_p_type;
  wire  prbNet_io_out_0_ready;
  wire  prbNet_io_out_0_valid;
  wire [1:0] prbNet_io_out_0_bits_header_src;
  wire [1:0] prbNet_io_out_0_bits_header_dst;
  wire [25:0] prbNet_io_out_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_0_bits_payload_p_type;
  wire  prbNet_io_out_1_ready;
  wire  prbNet_io_out_1_valid;
  wire [1:0] prbNet_io_out_1_bits_header_src;
  wire [1:0] prbNet_io_out_1_bits_header_dst;
  wire [25:0] prbNet_io_out_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_1_bits_payload_p_type;
  wire  prbNet_io_out_2_ready;
  wire  prbNet_io_out_2_valid;
  wire [1:0] prbNet_io_out_2_bits_header_src;
  wire [1:0] prbNet_io_out_2_bits_header_dst;
  wire [25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_2_bits_payload_p_type;
  wire  prbNet_io_out_3_ready;
  wire  prbNet_io_out_3_valid;
  wire [1:0] prbNet_io_out_3_bits_header_src;
  wire [1:0] prbNet_io_out_3_bits_header_dst;
  wire [25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_3_bits_payload_p_type;
  wire  gntNet_clk;
  wire  gntNet_reset;
  wire  gntNet_io_in_0_ready;
  wire  gntNet_io_in_0_valid;
  wire [1:0] gntNet_io_in_0_bits_header_src;
  wire [1:0] gntNet_io_in_0_bits_header_dst;
  wire [2:0] gntNet_io_in_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_0_bits_payload_manager_xact_id;
  wire  gntNet_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_0_bits_payload_g_type;
  wire [63:0] gntNet_io_in_0_bits_payload_data;
  wire  gntNet_io_in_1_ready;
  wire  gntNet_io_in_1_valid;
  wire [1:0] gntNet_io_in_1_bits_header_src;
  wire [1:0] gntNet_io_in_1_bits_header_dst;
  wire [2:0] gntNet_io_in_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_1_bits_payload_manager_xact_id;
  wire  gntNet_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_1_bits_payload_g_type;
  wire [63:0] gntNet_io_in_1_bits_payload_data;
  wire  gntNet_io_in_2_ready;
  wire  gntNet_io_in_2_valid;
  wire [1:0] gntNet_io_in_2_bits_header_src;
  wire [1:0] gntNet_io_in_2_bits_header_dst;
  wire [2:0] gntNet_io_in_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_2_bits_payload_manager_xact_id;
  wire  gntNet_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_2_bits_payload_g_type;
  wire [63:0] gntNet_io_in_2_bits_payload_data;
  wire  gntNet_io_in_3_ready;
  wire  gntNet_io_in_3_valid;
  wire [1:0] gntNet_io_in_3_bits_header_src;
  wire [1:0] gntNet_io_in_3_bits_header_dst;
  wire [2:0] gntNet_io_in_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_3_bits_payload_manager_xact_id;
  wire  gntNet_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_3_bits_payload_g_type;
  wire [63:0] gntNet_io_in_3_bits_payload_data;
  wire  gntNet_io_out_0_ready;
  wire  gntNet_io_out_0_valid;
  wire [1:0] gntNet_io_out_0_bits_header_src;
  wire [1:0] gntNet_io_out_0_bits_header_dst;
  wire [2:0] gntNet_io_out_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_0_bits_payload_manager_xact_id;
  wire  gntNet_io_out_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_0_bits_payload_g_type;
  wire [63:0] gntNet_io_out_0_bits_payload_data;
  wire  gntNet_io_out_1_ready;
  wire  gntNet_io_out_1_valid;
  wire [1:0] gntNet_io_out_1_bits_header_src;
  wire [1:0] gntNet_io_out_1_bits_header_dst;
  wire [2:0] gntNet_io_out_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire  gntNet_io_out_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_1_bits_payload_g_type;
  wire [63:0] gntNet_io_out_1_bits_payload_data;
  wire  gntNet_io_out_2_ready;
  wire  gntNet_io_out_2_valid;
  wire [1:0] gntNet_io_out_2_bits_header_src;
  wire [1:0] gntNet_io_out_2_bits_header_dst;
  wire [2:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire  gntNet_io_out_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_2_bits_payload_g_type;
  wire [63:0] gntNet_io_out_2_bits_payload_data;
  wire  gntNet_io_out_3_ready;
  wire  gntNet_io_out_3_valid;
  wire [1:0] gntNet_io_out_3_bits_header_src;
  wire [1:0] gntNet_io_out_3_bits_header_dst;
  wire [2:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire  gntNet_io_out_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_3_bits_payload_g_type;
  wire [63:0] gntNet_io_out_3_bits_payload_data;
  wire  ackNet_clk;
  wire  ackNet_reset;
  wire  ackNet_io_in_0_ready;
  wire  ackNet_io_in_0_valid;
  wire [1:0] ackNet_io_in_0_bits_header_src;
  wire [1:0] ackNet_io_in_0_bits_header_dst;
  wire [2:0] ackNet_io_in_0_bits_payload_manager_xact_id;
  wire  ackNet_io_in_1_ready;
  wire  ackNet_io_in_1_valid;
  wire [1:0] ackNet_io_in_1_bits_header_src;
  wire [1:0] ackNet_io_in_1_bits_header_dst;
  wire [2:0] ackNet_io_in_1_bits_payload_manager_xact_id;
  wire  ackNet_io_in_2_ready;
  wire  ackNet_io_in_2_valid;
  wire [1:0] ackNet_io_in_2_bits_header_src;
  wire [1:0] ackNet_io_in_2_bits_header_dst;
  wire [2:0] ackNet_io_in_2_bits_payload_manager_xact_id;
  wire  ackNet_io_in_3_ready;
  wire  ackNet_io_in_3_valid;
  wire [1:0] ackNet_io_in_3_bits_header_src;
  wire [1:0] ackNet_io_in_3_bits_header_dst;
  wire [2:0] ackNet_io_in_3_bits_payload_manager_xact_id;
  wire  ackNet_io_out_0_ready;
  wire  ackNet_io_out_0_valid;
  wire [1:0] ackNet_io_out_0_bits_header_src;
  wire [1:0] ackNet_io_out_0_bits_header_dst;
  wire [2:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire  ackNet_io_out_1_ready;
  wire  ackNet_io_out_1_valid;
  wire [1:0] ackNet_io_out_1_bits_header_src;
  wire [1:0] ackNet_io_out_1_bits_header_dst;
  wire [2:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire  ackNet_io_out_2_ready;
  wire  ackNet_io_out_2_valid;
  wire [1:0] ackNet_io_out_2_bits_header_src;
  wire [1:0] ackNet_io_out_2_bits_header_dst;
  wire [2:0] ackNet_io_out_2_bits_payload_manager_xact_id;
  wire  ackNet_io_out_3_ready;
  wire  ackNet_io_out_3_valid;
  wire [1:0] ackNet_io_out_3_bits_header_src;
  wire [1:0] ackNet_io_out_3_bits_header_dst;
  wire [2:0] ackNet_io_out_3_bits_payload_manager_xact_id;
  wire  T_12724_ready;
  wire  T_12724_valid;
  wire [1:0] T_12724_bits_header_src;
  wire [1:0] T_12724_bits_header_dst;
  wire [25:0] T_12724_bits_payload_addr_block;
  wire [1:0] T_12724_bits_payload_client_xact_id;
  wire [2:0] T_12724_bits_payload_addr_beat;
  wire  T_12724_bits_payload_is_builtin_type;
  wire [2:0] T_12724_bits_payload_a_type;
  wire [10:0] T_12724_bits_payload_union;
  wire [63:0] T_12724_bits_payload_data;
  wire [2:0] T_12952;
  wire [1:0] T_12953;
  wire  T_13294_ready;
  wire  T_13294_valid;
  wire [1:0] T_13294_bits_header_src;
  wire [1:0] T_13294_bits_header_dst;
  wire [25:0] T_13294_bits_payload_addr_block;
  wire [1:0] T_13294_bits_payload_client_xact_id;
  wire [2:0] T_13294_bits_payload_addr_beat;
  wire  T_13294_bits_payload_is_builtin_type;
  wire [2:0] T_13294_bits_payload_a_type;
  wire [10:0] T_13294_bits_payload_union;
  wire [63:0] T_13294_bits_payload_data;
  wire [2:0] T_13522;
  wire [1:0] T_13523;
  wire  T_13624_ready;
  wire  T_13624_valid;
  wire [1:0] T_13624_bits_header_src;
  wire [1:0] T_13624_bits_header_dst;
  wire [25:0] T_13624_bits_payload_addr_block;
  wire [1:0] T_13624_bits_payload_client_xact_id;
  wire [2:0] T_13624_bits_payload_addr_beat;
  wire  T_13624_bits_payload_is_builtin_type;
  wire [2:0] T_13624_bits_payload_a_type;
  wire [10:0] T_13624_bits_payload_union;
  wire [63:0] T_13624_bits_payload_data;
  wire [2:0] T_13692;
  wire [1:0] T_13693;
  wire  T_13794_ready;
  wire  T_13794_valid;
  wire [1:0] T_13794_bits_header_src;
  wire [1:0] T_13794_bits_header_dst;
  wire [25:0] T_13794_bits_payload_addr_block;
  wire [1:0] T_13794_bits_payload_client_xact_id;
  wire [2:0] T_13794_bits_payload_addr_beat;
  wire  T_13794_bits_payload_is_builtin_type;
  wire [2:0] T_13794_bits_payload_a_type;
  wire [10:0] T_13794_bits_payload_union;
  wire [63:0] T_13794_bits_payload_data;
  wire [2:0] T_13862;
  wire [1:0] T_13863;
  wire  T_14201_ready;
  wire  T_14201_valid;
  wire [1:0] T_14201_bits_header_src;
  wire [1:0] T_14201_bits_header_dst;
  wire [2:0] T_14201_bits_payload_addr_beat;
  wire [25:0] T_14201_bits_payload_addr_block;
  wire [1:0] T_14201_bits_payload_client_xact_id;
  wire  T_14201_bits_payload_voluntary;
  wire [2:0] T_14201_bits_payload_r_type;
  wire [63:0] T_14201_bits_payload_data;
  wire [2:0] T_14427;
  wire [1:0] T_14428;
  wire  T_14766_ready;
  wire  T_14766_valid;
  wire [1:0] T_14766_bits_header_src;
  wire [1:0] T_14766_bits_header_dst;
  wire [2:0] T_14766_bits_payload_addr_beat;
  wire [25:0] T_14766_bits_payload_addr_block;
  wire [1:0] T_14766_bits_payload_client_xact_id;
  wire  T_14766_bits_payload_voluntary;
  wire [2:0] T_14766_bits_payload_r_type;
  wire [63:0] T_14766_bits_payload_data;
  wire [2:0] T_14992;
  wire [1:0] T_14993;
  wire  T_15091_ready;
  wire  T_15091_valid;
  wire [1:0] T_15091_bits_header_src;
  wire [1:0] T_15091_bits_header_dst;
  wire [2:0] T_15091_bits_payload_addr_beat;
  wire [25:0] T_15091_bits_payload_addr_block;
  wire [1:0] T_15091_bits_payload_client_xact_id;
  wire  T_15091_bits_payload_voluntary;
  wire [2:0] T_15091_bits_payload_r_type;
  wire [63:0] T_15091_bits_payload_data;
  wire [2:0] T_15157;
  wire [1:0] T_15158;
  wire  T_15256_ready;
  wire  T_15256_valid;
  wire [1:0] T_15256_bits_header_src;
  wire [1:0] T_15256_bits_header_dst;
  wire [2:0] T_15256_bits_payload_addr_beat;
  wire [25:0] T_15256_bits_payload_addr_block;
  wire [1:0] T_15256_bits_payload_client_xact_id;
  wire  T_15256_bits_payload_voluntary;
  wire [2:0] T_15256_bits_payload_r_type;
  wire [63:0] T_15256_bits_payload_data;
  wire [2:0] T_15322;
  wire [1:0] T_15323;
  wire  T_15409_ready;
  wire  T_15409_valid;
  wire [1:0] T_15409_bits_header_src;
  wire [1:0] T_15409_bits_header_dst;
  wire [25:0] T_15409_bits_payload_addr_block;
  wire [1:0] T_15409_bits_payload_p_type;
  wire [2:0] T_15467;
  wire [1:0] T_15468;
  wire  T_15554_ready;
  wire  T_15554_valid;
  wire [1:0] T_15554_bits_header_src;
  wire [1:0] T_15554_bits_header_dst;
  wire [25:0] T_15554_bits_payload_addr_block;
  wire [1:0] T_15554_bits_payload_p_type;
  wire [2:0] T_15612;
  wire [1:0] T_15613;
  wire  T_15939_ready;
  wire  T_15939_valid;
  wire [1:0] T_15939_bits_header_src;
  wire [1:0] T_15939_bits_header_dst;
  wire [25:0] T_15939_bits_payload_addr_block;
  wire [1:0] T_15939_bits_payload_p_type;
  wire [2:0] T_16157;
  wire [1:0] T_16158;
  wire  T_16484_ready;
  wire  T_16484_valid;
  wire [1:0] T_16484_bits_header_src;
  wire [1:0] T_16484_bits_header_dst;
  wire [25:0] T_16484_bits_payload_addr_block;
  wire [1:0] T_16484_bits_payload_p_type;
  wire [2:0] T_16702;
  wire [1:0] T_16703;
  wire  T_16801_ready;
  wire  T_16801_valid;
  wire [1:0] T_16801_bits_header_src;
  wire [1:0] T_16801_bits_header_dst;
  wire [2:0] T_16801_bits_payload_addr_beat;
  wire [1:0] T_16801_bits_payload_client_xact_id;
  wire [2:0] T_16801_bits_payload_manager_xact_id;
  wire  T_16801_bits_payload_is_builtin_type;
  wire [3:0] T_16801_bits_payload_g_type;
  wire [63:0] T_16801_bits_payload_data;
  wire [2:0] T_16867;
  wire [1:0] T_16868;
  wire  T_16966_ready;
  wire  T_16966_valid;
  wire [1:0] T_16966_bits_header_src;
  wire [1:0] T_16966_bits_header_dst;
  wire [2:0] T_16966_bits_payload_addr_beat;
  wire [1:0] T_16966_bits_payload_client_xact_id;
  wire [2:0] T_16966_bits_payload_manager_xact_id;
  wire  T_16966_bits_payload_is_builtin_type;
  wire [3:0] T_16966_bits_payload_g_type;
  wire [63:0] T_16966_bits_payload_data;
  wire [2:0] T_17032;
  wire [1:0] T_17033;
  wire  T_17371_ready;
  wire  T_17371_valid;
  wire [1:0] T_17371_bits_header_src;
  wire [1:0] T_17371_bits_header_dst;
  wire [2:0] T_17371_bits_payload_addr_beat;
  wire [1:0] T_17371_bits_payload_client_xact_id;
  wire [2:0] T_17371_bits_payload_manager_xact_id;
  wire  T_17371_bits_payload_is_builtin_type;
  wire [3:0] T_17371_bits_payload_g_type;
  wire [63:0] T_17371_bits_payload_data;
  wire [2:0] T_17597;
  wire [1:0] T_17598;
  wire  T_17936_ready;
  wire  T_17936_valid;
  wire [1:0] T_17936_bits_header_src;
  wire [1:0] T_17936_bits_header_dst;
  wire [2:0] T_17936_bits_payload_addr_beat;
  wire [1:0] T_17936_bits_payload_client_xact_id;
  wire [2:0] T_17936_bits_payload_manager_xact_id;
  wire  T_17936_bits_payload_is_builtin_type;
  wire [3:0] T_17936_bits_payload_g_type;
  wire [63:0] T_17936_bits_payload_data;
  wire [2:0] T_18162;
  wire [1:0] T_18163;
  wire  T_18486_ready;
  wire  T_18486_valid;
  wire [1:0] T_18486_bits_header_src;
  wire [1:0] T_18486_bits_header_dst;
  wire [2:0] T_18486_bits_payload_manager_xact_id;
  wire [2:0] T_18702;
  wire [1:0] T_18703;
  wire  T_19026_ready;
  wire  T_19026_valid;
  wire [1:0] T_19026_bits_header_src;
  wire [1:0] T_19026_bits_header_dst;
  wire [2:0] T_19026_bits_payload_manager_xact_id;
  wire [2:0] T_19242;
  wire [1:0] T_19243;
  wire  T_19326_ready;
  wire  T_19326_valid;
  wire [1:0] T_19326_bits_header_src;
  wire [1:0] T_19326_bits_header_dst;
  wire [2:0] T_19326_bits_payload_manager_xact_id;
  wire [2:0] T_19382;
  wire [1:0] T_19383;
  wire  T_19466_ready;
  wire  T_19466_valid;
  wire [1:0] T_19466_bits_header_src;
  wire [1:0] T_19466_bits_header_dst;
  wire [2:0] T_19466_bits_payload_manager_xact_id;
  wire [2:0] T_19522;
  wire [1:0] T_19523;
  wire [1:0] GEN_0;
  reg [31:0] GEN_64;
  wire [1:0] GEN_1;
  reg [31:0] GEN_65;
  wire [25:0] GEN_2;
  reg [31:0] GEN_66;
  wire [1:0] GEN_3;
  reg [31:0] GEN_67;
  wire [2:0] GEN_4;
  reg [31:0] GEN_68;
  wire  GEN_5;
  reg [31:0] GEN_69;
  wire [2:0] GEN_6;
  reg [31:0] GEN_70;
  wire [10:0] GEN_7;
  reg [31:0] GEN_71;
  wire [63:0] GEN_8;
  reg [63:0] GEN_72;
  wire [1:0] GEN_9;
  reg [31:0] GEN_73;
  wire [1:0] GEN_10;
  reg [31:0] GEN_74;
  wire [25:0] GEN_11;
  reg [31:0] GEN_75;
  wire [1:0] GEN_12;
  reg [31:0] GEN_76;
  wire [2:0] GEN_13;
  reg [31:0] GEN_77;
  wire  GEN_14;
  reg [31:0] GEN_78;
  wire [2:0] GEN_15;
  reg [31:0] GEN_79;
  wire [10:0] GEN_16;
  reg [31:0] GEN_80;
  wire [63:0] GEN_17;
  reg [63:0] GEN_81;
  wire [1:0] GEN_18;
  reg [31:0] GEN_82;
  wire [1:0] GEN_19;
  reg [31:0] GEN_83;
  wire [2:0] GEN_20;
  reg [31:0] GEN_84;
  wire [25:0] GEN_21;
  reg [31:0] GEN_85;
  wire [1:0] GEN_22;
  reg [31:0] GEN_86;
  wire  GEN_23;
  reg [31:0] GEN_87;
  wire [2:0] GEN_24;
  reg [31:0] GEN_88;
  wire [63:0] GEN_25;
  reg [63:0] GEN_89;
  wire [1:0] GEN_26;
  reg [31:0] GEN_90;
  wire [1:0] GEN_27;
  reg [31:0] GEN_91;
  wire [2:0] GEN_28;
  reg [31:0] GEN_92;
  wire [25:0] GEN_29;
  reg [31:0] GEN_93;
  wire [1:0] GEN_30;
  reg [31:0] GEN_94;
  wire  GEN_31;
  reg [31:0] GEN_95;
  wire [2:0] GEN_32;
  reg [31:0] GEN_96;
  wire [63:0] GEN_33;
  reg [63:0] GEN_97;
  wire [1:0] GEN_34;
  reg [31:0] GEN_98;
  wire [1:0] GEN_35;
  reg [31:0] GEN_99;
  wire [25:0] GEN_36;
  reg [31:0] GEN_100;
  wire [1:0] GEN_37;
  reg [31:0] GEN_101;
  wire [1:0] GEN_38;
  reg [31:0] GEN_102;
  wire [1:0] GEN_39;
  reg [31:0] GEN_103;
  wire [25:0] GEN_40;
  reg [31:0] GEN_104;
  wire [1:0] GEN_41;
  reg [31:0] GEN_105;
  wire [1:0] GEN_42;
  reg [31:0] GEN_106;
  wire [1:0] GEN_43;
  reg [31:0] GEN_107;
  wire [2:0] GEN_44;
  reg [31:0] GEN_108;
  wire [1:0] GEN_45;
  reg [31:0] GEN_109;
  wire [2:0] GEN_46;
  reg [31:0] GEN_110;
  wire  GEN_47;
  reg [31:0] GEN_111;
  wire [3:0] GEN_48;
  reg [31:0] GEN_112;
  wire [63:0] GEN_49;
  reg [63:0] GEN_113;
  wire [1:0] GEN_50;
  reg [31:0] GEN_114;
  wire [1:0] GEN_51;
  reg [31:0] GEN_115;
  wire [2:0] GEN_52;
  reg [31:0] GEN_116;
  wire [1:0] GEN_53;
  reg [31:0] GEN_117;
  wire [2:0] GEN_54;
  reg [31:0] GEN_118;
  wire  GEN_55;
  reg [31:0] GEN_119;
  wire [3:0] GEN_56;
  reg [31:0] GEN_120;
  wire [63:0] GEN_57;
  reg [63:0] GEN_121;
  wire [1:0] GEN_58;
  reg [31:0] GEN_122;
  wire [1:0] GEN_59;
  reg [31:0] GEN_123;
  wire [2:0] GEN_60;
  reg [31:0] GEN_124;
  wire [1:0] GEN_61;
  reg [31:0] GEN_125;
  wire [1:0] GEN_62;
  reg [31:0] GEN_126;
  wire [2:0] GEN_63;
  reg [31:0] GEN_127;
  TileLinkEnqueuer TileLinkEnqueuer_4 (
    .clk(TileLinkEnqueuer_4_clk),
    .reset(TileLinkEnqueuer_4_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_4_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_4_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_4_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_4_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_4_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_4_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_4_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_4_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_4_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_4_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_4_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_4_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_4_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_4_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_4_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_4_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_4_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_4_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_4_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_4_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_4_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_4_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_4_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_4_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_4_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_4_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_4_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_4_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_4_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_4_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_4_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_4_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_4_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_4_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_4_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_4_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_4_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_4_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_4_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_4_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_4_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_4_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_4_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_4_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_4_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_4_io_manager_release_bits_payload_data)
  );
  ClientTileLinkNetworkPort ClientTileLinkNetworkPort_1 (
    .clk(ClientTileLinkNetworkPort_1_clk),
    .reset(ClientTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_probe_ready(ClientTileLinkNetworkPort_1_io_client_probe_ready),
    .io_client_probe_valid(ClientTileLinkNetworkPort_1_io_client_probe_valid),
    .io_client_probe_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block),
    .io_client_probe_bits_p_type(ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type),
    .io_client_release_ready(ClientTileLinkNetworkPort_1_io_client_release_ready),
    .io_client_release_valid(ClientTileLinkNetworkPort_1_io_client_release_valid),
    .io_client_release_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat),
    .io_client_release_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block),
    .io_client_release_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id),
    .io_client_release_bits_voluntary(ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary),
    .io_client_release_bits_r_type(ClientTileLinkNetworkPort_1_io_client_release_bits_r_type),
    .io_client_release_bits_data(ClientTileLinkNetworkPort_1_io_client_release_bits_data),
    .io_client_grant_ready(ClientTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_client_grant_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id),
    .io_client_finish_ready(ClientTileLinkNetworkPort_1_io_client_finish_ready),
    .io_client_finish_valid(ClientTileLinkNetworkPort_1_io_client_finish_valid),
    .io_client_finish_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id),
    .io_client_finish_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id),
    .io_network_acquire_ready(ClientTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_1_1 (
    .clk(TileLinkEnqueuer_1_1_clk),
    .reset(TileLinkEnqueuer_1_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_1_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_1_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_1_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_1_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_1_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_1_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_1_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_1_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_1_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_1_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_1_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_1_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_1_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_1_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_1_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_1_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_1_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_1_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_1_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort ClientUncachedTileLinkNetworkPort_1 (
    .clk(ClientUncachedTileLinkNetworkPort_1_clk),
    .reset(ClientUncachedTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort_2 (
    .clk(ManagerTileLinkNetworkPort_2_clk),
    .reset(ManagerTileLinkNetworkPort_2_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_2_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_2_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_2_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_2_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_2_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_2_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_2_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_2_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_2_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_2_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_2_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_2_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_2_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_2_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_2_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_2_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_2_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_2_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_2_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_2_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_2_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_2_1 (
    .clk(TileLinkEnqueuer_2_1_clk),
    .reset(TileLinkEnqueuer_2_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_2_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_2_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_2_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_2_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_2_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_2_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_2_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_2_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_2_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_2_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_2_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_2_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_2_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_2_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_2_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_2_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_2_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_2_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_2_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_2_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_2_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_2_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_2_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_2_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_2_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_2_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_2_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort_1_1 (
    .clk(ManagerTileLinkNetworkPort_1_1_clk),
    .reset(ManagerTileLinkNetworkPort_1_1_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_1_1_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_1_1_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_1_1_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_1_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_1_1_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_1_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_1_1_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_1_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_1_1_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_1_1_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_3_1 (
    .clk(TileLinkEnqueuer_3_1_clk),
    .reset(TileLinkEnqueuer_3_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_3_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_3_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_3_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_3_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_3_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_3_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_3_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_3_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_3_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_3_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_3_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_3_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_3_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_3_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_3_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_3_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_3_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_3_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_3_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_3_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_3_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_3_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_3_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_3_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_3_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_3_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_3_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data)
  );
  BasicBus acqNet (
    .clk(acqNet_clk),
    .reset(acqNet_reset),
    .io_in_0_ready(acqNet_io_in_0_ready),
    .io_in_0_valid(acqNet_io_in_0_valid),
    .io_in_0_bits_header_src(acqNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(acqNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(acqNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(acqNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(acqNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(acqNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(acqNet_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(acqNet_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(acqNet_io_in_0_bits_payload_data),
    .io_in_1_ready(acqNet_io_in_1_ready),
    .io_in_1_valid(acqNet_io_in_1_valid),
    .io_in_1_bits_header_src(acqNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(acqNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(acqNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(acqNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(acqNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(acqNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(acqNet_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(acqNet_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(acqNet_io_in_1_bits_payload_data),
    .io_in_2_ready(acqNet_io_in_2_ready),
    .io_in_2_valid(acqNet_io_in_2_valid),
    .io_in_2_bits_header_src(acqNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(acqNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(acqNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(acqNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(acqNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(acqNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(acqNet_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(acqNet_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(acqNet_io_in_2_bits_payload_data),
    .io_in_3_ready(acqNet_io_in_3_ready),
    .io_in_3_valid(acqNet_io_in_3_valid),
    .io_in_3_bits_header_src(acqNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(acqNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(acqNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(acqNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(acqNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(acqNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(acqNet_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(acqNet_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(acqNet_io_in_3_bits_payload_data),
    .io_out_0_ready(acqNet_io_out_0_ready),
    .io_out_0_valid(acqNet_io_out_0_valid),
    .io_out_0_bits_header_src(acqNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(acqNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(acqNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(acqNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_addr_beat(acqNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_is_builtin_type(acqNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_a_type(acqNet_io_out_0_bits_payload_a_type),
    .io_out_0_bits_payload_union(acqNet_io_out_0_bits_payload_union),
    .io_out_0_bits_payload_data(acqNet_io_out_0_bits_payload_data),
    .io_out_1_ready(acqNet_io_out_1_ready),
    .io_out_1_valid(acqNet_io_out_1_valid),
    .io_out_1_bits_header_src(acqNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(acqNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(acqNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(acqNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_addr_beat(acqNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_is_builtin_type(acqNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_a_type(acqNet_io_out_1_bits_payload_a_type),
    .io_out_1_bits_payload_union(acqNet_io_out_1_bits_payload_union),
    .io_out_1_bits_payload_data(acqNet_io_out_1_bits_payload_data),
    .io_out_2_ready(acqNet_io_out_2_ready),
    .io_out_2_valid(acqNet_io_out_2_valid),
    .io_out_2_bits_header_src(acqNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(acqNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(acqNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(acqNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_addr_beat(acqNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_is_builtin_type(acqNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_a_type(acqNet_io_out_2_bits_payload_a_type),
    .io_out_2_bits_payload_union(acqNet_io_out_2_bits_payload_union),
    .io_out_2_bits_payload_data(acqNet_io_out_2_bits_payload_data),
    .io_out_3_ready(acqNet_io_out_3_ready),
    .io_out_3_valid(acqNet_io_out_3_valid),
    .io_out_3_bits_header_src(acqNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(acqNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(acqNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(acqNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_addr_beat(acqNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_is_builtin_type(acqNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_a_type(acqNet_io_out_3_bits_payload_a_type),
    .io_out_3_bits_payload_union(acqNet_io_out_3_bits_payload_union),
    .io_out_3_bits_payload_data(acqNet_io_out_3_bits_payload_data)
  );
  BasicBus_1 relNet (
    .clk(relNet_clk),
    .reset(relNet_reset),
    .io_in_0_ready(relNet_io_in_0_ready),
    .io_in_0_valid(relNet_io_in_0_valid),
    .io_in_0_bits_header_src(relNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(relNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(relNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(relNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(relNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(relNet_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(relNet_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(relNet_io_in_0_bits_payload_data),
    .io_in_1_ready(relNet_io_in_1_ready),
    .io_in_1_valid(relNet_io_in_1_valid),
    .io_in_1_bits_header_src(relNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(relNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(relNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(relNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(relNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(relNet_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(relNet_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(relNet_io_in_1_bits_payload_data),
    .io_in_2_ready(relNet_io_in_2_ready),
    .io_in_2_valid(relNet_io_in_2_valid),
    .io_in_2_bits_header_src(relNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(relNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(relNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(relNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(relNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(relNet_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(relNet_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(relNet_io_in_2_bits_payload_data),
    .io_in_3_ready(relNet_io_in_3_ready),
    .io_in_3_valid(relNet_io_in_3_valid),
    .io_in_3_bits_header_src(relNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(relNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(relNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(relNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(relNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(relNet_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(relNet_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(relNet_io_in_3_bits_payload_data),
    .io_out_0_ready(relNet_io_out_0_ready),
    .io_out_0_valid(relNet_io_out_0_valid),
    .io_out_0_bits_header_src(relNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(relNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(relNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_addr_block(relNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(relNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_voluntary(relNet_io_out_0_bits_payload_voluntary),
    .io_out_0_bits_payload_r_type(relNet_io_out_0_bits_payload_r_type),
    .io_out_0_bits_payload_data(relNet_io_out_0_bits_payload_data),
    .io_out_1_ready(relNet_io_out_1_ready),
    .io_out_1_valid(relNet_io_out_1_valid),
    .io_out_1_bits_header_src(relNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(relNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(relNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_addr_block(relNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(relNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_voluntary(relNet_io_out_1_bits_payload_voluntary),
    .io_out_1_bits_payload_r_type(relNet_io_out_1_bits_payload_r_type),
    .io_out_1_bits_payload_data(relNet_io_out_1_bits_payload_data),
    .io_out_2_ready(relNet_io_out_2_ready),
    .io_out_2_valid(relNet_io_out_2_valid),
    .io_out_2_bits_header_src(relNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(relNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(relNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_addr_block(relNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(relNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_voluntary(relNet_io_out_2_bits_payload_voluntary),
    .io_out_2_bits_payload_r_type(relNet_io_out_2_bits_payload_r_type),
    .io_out_2_bits_payload_data(relNet_io_out_2_bits_payload_data),
    .io_out_3_ready(relNet_io_out_3_ready),
    .io_out_3_valid(relNet_io_out_3_valid),
    .io_out_3_bits_header_src(relNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(relNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(relNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_addr_block(relNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(relNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_voluntary(relNet_io_out_3_bits_payload_voluntary),
    .io_out_3_bits_payload_r_type(relNet_io_out_3_bits_payload_r_type),
    .io_out_3_bits_payload_data(relNet_io_out_3_bits_payload_data)
  );
  BasicBus_2 prbNet (
    .clk(prbNet_clk),
    .reset(prbNet_reset),
    .io_in_0_ready(prbNet_io_in_0_ready),
    .io_in_0_valid(prbNet_io_in_0_valid),
    .io_in_0_bits_header_src(prbNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(prbNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(prbNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(prbNet_io_in_0_bits_payload_p_type),
    .io_in_1_ready(prbNet_io_in_1_ready),
    .io_in_1_valid(prbNet_io_in_1_valid),
    .io_in_1_bits_header_src(prbNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(prbNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(prbNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(prbNet_io_in_1_bits_payload_p_type),
    .io_in_2_ready(prbNet_io_in_2_ready),
    .io_in_2_valid(prbNet_io_in_2_valid),
    .io_in_2_bits_header_src(prbNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(prbNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(prbNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(prbNet_io_in_2_bits_payload_p_type),
    .io_in_3_ready(prbNet_io_in_3_ready),
    .io_in_3_valid(prbNet_io_in_3_valid),
    .io_in_3_bits_header_src(prbNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(prbNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(prbNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(prbNet_io_in_3_bits_payload_p_type),
    .io_out_0_ready(prbNet_io_out_0_ready),
    .io_out_0_valid(prbNet_io_out_0_valid),
    .io_out_0_bits_header_src(prbNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(prbNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(prbNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_p_type(prbNet_io_out_0_bits_payload_p_type),
    .io_out_1_ready(prbNet_io_out_1_ready),
    .io_out_1_valid(prbNet_io_out_1_valid),
    .io_out_1_bits_header_src(prbNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(prbNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(prbNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_p_type(prbNet_io_out_1_bits_payload_p_type),
    .io_out_2_ready(prbNet_io_out_2_ready),
    .io_out_2_valid(prbNet_io_out_2_valid),
    .io_out_2_bits_header_src(prbNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(prbNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(prbNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_p_type(prbNet_io_out_2_bits_payload_p_type),
    .io_out_3_ready(prbNet_io_out_3_ready),
    .io_out_3_valid(prbNet_io_out_3_valid),
    .io_out_3_bits_header_src(prbNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(prbNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(prbNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_p_type(prbNet_io_out_3_bits_payload_p_type)
  );
  BasicBus_3 gntNet (
    .clk(gntNet_clk),
    .reset(gntNet_reset),
    .io_in_0_ready(gntNet_io_in_0_ready),
    .io_in_0_valid(gntNet_io_in_0_valid),
    .io_in_0_bits_header_src(gntNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(gntNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(gntNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(gntNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(gntNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(gntNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(gntNet_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(gntNet_io_in_0_bits_payload_data),
    .io_in_1_ready(gntNet_io_in_1_ready),
    .io_in_1_valid(gntNet_io_in_1_valid),
    .io_in_1_bits_header_src(gntNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(gntNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(gntNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(gntNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(gntNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(gntNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(gntNet_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(gntNet_io_in_1_bits_payload_data),
    .io_in_2_ready(gntNet_io_in_2_ready),
    .io_in_2_valid(gntNet_io_in_2_valid),
    .io_in_2_bits_header_src(gntNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(gntNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(gntNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(gntNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(gntNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(gntNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(gntNet_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(gntNet_io_in_2_bits_payload_data),
    .io_in_3_ready(gntNet_io_in_3_ready),
    .io_in_3_valid(gntNet_io_in_3_valid),
    .io_in_3_bits_header_src(gntNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(gntNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(gntNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(gntNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(gntNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(gntNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(gntNet_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(gntNet_io_in_3_bits_payload_data),
    .io_out_0_ready(gntNet_io_out_0_ready),
    .io_out_0_valid(gntNet_io_out_0_valid),
    .io_out_0_bits_header_src(gntNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(gntNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(gntNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_client_xact_id(gntNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_manager_xact_id(gntNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_0_bits_payload_is_builtin_type(gntNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_g_type(gntNet_io_out_0_bits_payload_g_type),
    .io_out_0_bits_payload_data(gntNet_io_out_0_bits_payload_data),
    .io_out_1_ready(gntNet_io_out_1_ready),
    .io_out_1_valid(gntNet_io_out_1_valid),
    .io_out_1_bits_header_src(gntNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(gntNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(gntNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_client_xact_id(gntNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_manager_xact_id(gntNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_1_bits_payload_is_builtin_type(gntNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_g_type(gntNet_io_out_1_bits_payload_g_type),
    .io_out_1_bits_payload_data(gntNet_io_out_1_bits_payload_data),
    .io_out_2_ready(gntNet_io_out_2_ready),
    .io_out_2_valid(gntNet_io_out_2_valid),
    .io_out_2_bits_header_src(gntNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(gntNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(gntNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_client_xact_id(gntNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_manager_xact_id(gntNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_2_bits_payload_is_builtin_type(gntNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_g_type(gntNet_io_out_2_bits_payload_g_type),
    .io_out_2_bits_payload_data(gntNet_io_out_2_bits_payload_data),
    .io_out_3_ready(gntNet_io_out_3_ready),
    .io_out_3_valid(gntNet_io_out_3_valid),
    .io_out_3_bits_header_src(gntNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(gntNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(gntNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_client_xact_id(gntNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_manager_xact_id(gntNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_3_bits_payload_is_builtin_type(gntNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_g_type(gntNet_io_out_3_bits_payload_g_type),
    .io_out_3_bits_payload_data(gntNet_io_out_3_bits_payload_data)
  );
  BasicBus_4 ackNet (
    .clk(ackNet_clk),
    .reset(ackNet_reset),
    .io_in_0_ready(ackNet_io_in_0_ready),
    .io_in_0_valid(ackNet_io_in_0_valid),
    .io_in_0_bits_header_src(ackNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(ackNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(ackNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(ackNet_io_in_1_ready),
    .io_in_1_valid(ackNet_io_in_1_valid),
    .io_in_1_bits_header_src(ackNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(ackNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(ackNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(ackNet_io_in_2_ready),
    .io_in_2_valid(ackNet_io_in_2_valid),
    .io_in_2_bits_header_src(ackNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(ackNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(ackNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(ackNet_io_in_3_ready),
    .io_in_3_valid(ackNet_io_in_3_valid),
    .io_in_3_bits_header_src(ackNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(ackNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(ackNet_io_in_3_bits_payload_manager_xact_id),
    .io_out_0_ready(ackNet_io_out_0_ready),
    .io_out_0_valid(ackNet_io_out_0_valid),
    .io_out_0_bits_header_src(ackNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(ackNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_manager_xact_id(ackNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_1_ready(ackNet_io_out_1_ready),
    .io_out_1_valid(ackNet_io_out_1_valid),
    .io_out_1_bits_header_src(ackNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(ackNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_manager_xact_id(ackNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_2_ready(ackNet_io_out_2_ready),
    .io_out_2_valid(ackNet_io_out_2_valid),
    .io_out_2_bits_header_src(ackNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(ackNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_manager_xact_id(ackNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_3_ready(ackNet_io_out_3_ready),
    .io_out_3_valid(ackNet_io_out_3_valid),
    .io_out_3_bits_header_src(ackNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(ackNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_manager_xact_id(ackNet_io_out_3_bits_payload_manager_xact_id)
  );
  assign io_clients_cached_0_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_cached_0_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_cached_0_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_cached_0_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_cached_0_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_cached_0_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_cached_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_cached_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_cached_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_cached_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_cached_0_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_cached_0_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_cached_0_grant_bits_manager_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  assign io_clients_cached_0_finish_ready = ClientTileLinkNetworkPort_1_io_client_finish_ready;
  assign io_clients_uncached_0_acquire_ready = ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_uncached_0_grant_valid = ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_uncached_0_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_0_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_0_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_0_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_0_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_uncached_0_grant_bits_data = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  assign TileLinkEnqueuer_4_clk = clk;
  assign TileLinkEnqueuer_4_reset = reset;
  assign TileLinkEnqueuer_4_io_client_acquire_valid = ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_src = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_union = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_4_io_client_grant_ready = ClientTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_4_io_client_finish_valid = ClientTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_src = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id = ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_client_probe_ready = ClientTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_4_io_client_release_valid = ClientTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_src = ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_r_type = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_acquire_ready = T_13624_ready;
  assign TileLinkEnqueuer_4_io_manager_grant_valid = T_17371_valid;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_src = T_17371_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_dst = T_17371_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat = T_17371_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id = T_17371_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id = T_17371_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type = T_17371_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type = T_17371_bits_payload_g_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_data = T_17371_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_finish_ready = T_19326_ready;
  assign TileLinkEnqueuer_4_io_manager_probe_valid = T_15939_valid;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_src = T_15939_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_dst = T_15939_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block = T_15939_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type = T_15939_bits_payload_p_type;
  assign TileLinkEnqueuer_4_io_manager_release_ready = T_15091_ready;
  assign ClientTileLinkNetworkPort_1_clk = clk;
  assign ClientTileLinkNetworkPort_1_reset = reset;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_cached_0_acquire_valid;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_cached_0_acquire_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_cached_0_acquire_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_cached_0_acquire_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_cached_0_acquire_bits_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_cached_0_acquire_bits_a_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_cached_0_acquire_bits_union;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_cached_0_acquire_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_probe_ready = io_clients_cached_0_probe_ready;
  assign ClientTileLinkNetworkPort_1_io_client_release_valid = io_clients_cached_0_release_valid;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat = io_clients_cached_0_release_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block = io_clients_cached_0_release_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id = io_clients_cached_0_release_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary = io_clients_cached_0_release_bits_voluntary;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_r_type = io_clients_cached_0_release_bits_r_type;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_data = io_clients_cached_0_release_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_grant_ready = io_clients_cached_0_grant_ready;
  assign ClientTileLinkNetworkPort_1_io_client_finish_valid = io_clients_cached_0_finish_valid;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id = io_clients_cached_0_finish_bits_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id = io_clients_cached_0_finish_bits_manager_id;
  assign ClientTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_4_io_client_acquire_ready;
  assign ClientTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_4_io_client_grant_valid;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  assign ClientTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_4_io_client_finish_ready;
  assign ClientTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_4_io_client_probe_valid;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  assign ClientTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_4_io_client_release_ready;
  assign TileLinkEnqueuer_1_1_clk = clk;
  assign TileLinkEnqueuer_1_1_reset = reset;
  assign TileLinkEnqueuer_1_1_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_1_1_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_1_1_io_client_release_valid = ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_acquire_ready = T_13794_ready;
  assign TileLinkEnqueuer_1_1_io_manager_grant_valid = T_17936_valid;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src = T_17936_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst = T_17936_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat = T_17936_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id = T_17936_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id = T_17936_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type = T_17936_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type = T_17936_bits_payload_g_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data = T_17936_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_finish_ready = T_19466_ready;
  assign TileLinkEnqueuer_1_1_io_manager_probe_valid = T_16484_valid;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src = T_16484_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst = T_16484_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block = T_16484_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type = T_16484_bits_payload_p_type;
  assign TileLinkEnqueuer_1_1_io_manager_release_ready = T_15256_ready;
  assign ClientUncachedTileLinkNetworkPort_1_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_1_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_uncached_0_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_uncached_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_uncached_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_uncached_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_uncached_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_uncached_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_uncached_0_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_uncached_0_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready = io_clients_uncached_0_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_1_1_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_1_1_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_1_1_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_1_1_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_1_1_io_client_release_ready;
  assign ManagerTileLinkNetworkPort_2_clk = clk;
  assign ManagerTileLinkNetworkPort_2_reset = reset;
  assign ManagerTileLinkNetworkPort_2_io_manager_acquire_ready = io_managers_0_acquire_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_valid = io_managers_0_grant_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat = io_managers_0_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id = io_managers_0_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id = io_managers_0_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type = io_managers_0_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type = io_managers_0_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data = io_managers_0_grant_bits_data;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id = io_managers_0_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_finish_ready = io_managers_0_finish_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_valid = io_managers_0_probe_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block = io_managers_0_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type = io_managers_0_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id = io_managers_0_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_release_ready = io_managers_0_release_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_valid = TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_2_io_network_grant_ready = TileLinkEnqueuer_2_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_valid = TileLinkEnqueuer_2_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_probe_ready = TileLinkEnqueuer_2_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_release_valid = TileLinkEnqueuer_2_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src = TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_2_1_clk = clk;
  assign TileLinkEnqueuer_2_1_reset = reset;
  assign TileLinkEnqueuer_2_1_io_client_acquire_valid = T_12724_valid;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src = T_12724_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst = T_12724_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block = T_12724_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id = T_12724_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat = T_12724_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type = T_12724_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type = T_12724_bits_payload_a_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union = T_12724_bits_payload_union;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data = T_12724_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_client_grant_ready = T_16801_ready;
  assign TileLinkEnqueuer_2_1_io_client_finish_valid = T_18486_valid;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_src = T_18486_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst = T_18486_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id = T_18486_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_probe_ready = T_15409_ready;
  assign TileLinkEnqueuer_2_1_io_client_release_valid = T_14201_valid;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_src = T_14201_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_dst = T_14201_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat = T_14201_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block = T_14201_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id = T_14201_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary = T_14201_bits_payload_voluntary;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type = T_14201_bits_payload_r_type;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_data = T_14201_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  assign TileLinkEnqueuer_2_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  assign TileLinkEnqueuer_2_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_2_1_io_manager_release_ready = ManagerTileLinkNetworkPort_2_io_network_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_clk = clk;
  assign ManagerTileLinkNetworkPort_1_1_reset = reset;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready = io_managers_1_acquire_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid = io_managers_1_grant_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat = io_managers_1_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id = io_managers_1_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id = io_managers_1_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type = io_managers_1_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type = io_managers_1_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data = io_managers_1_grant_bits_data;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id = io_managers_1_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready = io_managers_1_finish_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid = io_managers_1_probe_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block = io_managers_1_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type = io_managers_1_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id = io_managers_1_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_release_ready = io_managers_1_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid = TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_1_1_io_network_grant_ready = TileLinkEnqueuer_3_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_valid = TileLinkEnqueuer_3_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_probe_ready = TileLinkEnqueuer_3_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_valid = TileLinkEnqueuer_3_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src = TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_3_1_clk = clk;
  assign TileLinkEnqueuer_3_1_reset = reset;
  assign TileLinkEnqueuer_3_1_io_client_acquire_valid = T_13294_valid;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src = T_13294_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst = T_13294_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block = T_13294_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id = T_13294_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat = T_13294_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type = T_13294_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type = T_13294_bits_payload_a_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union = T_13294_bits_payload_union;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data = T_13294_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_client_grant_ready = T_16966_ready;
  assign TileLinkEnqueuer_3_1_io_client_finish_valid = T_19026_valid;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_src = T_19026_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst = T_19026_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id = T_19026_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_probe_ready = T_15554_ready;
  assign TileLinkEnqueuer_3_1_io_client_release_valid = T_14766_valid;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_src = T_14766_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_dst = T_14766_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat = T_14766_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block = T_14766_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id = T_14766_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary = T_14766_bits_payload_voluntary;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type = T_14766_bits_payload_r_type;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_data = T_14766_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  assign TileLinkEnqueuer_3_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  assign TileLinkEnqueuer_3_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_3_1_io_manager_release_ready = ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  assign acqNet_clk = clk;
  assign acqNet_reset = reset;
  assign acqNet_io_in_0_valid = 1'h0;
  assign acqNet_io_in_0_bits_header_src = GEN_0;
  assign acqNet_io_in_0_bits_header_dst = GEN_1;
  assign acqNet_io_in_0_bits_payload_addr_block = GEN_2;
  assign acqNet_io_in_0_bits_payload_client_xact_id = GEN_3;
  assign acqNet_io_in_0_bits_payload_addr_beat = GEN_4;
  assign acqNet_io_in_0_bits_payload_is_builtin_type = GEN_5;
  assign acqNet_io_in_0_bits_payload_a_type = GEN_6;
  assign acqNet_io_in_0_bits_payload_union = GEN_7;
  assign acqNet_io_in_0_bits_payload_data = GEN_8;
  assign acqNet_io_in_1_valid = 1'h0;
  assign acqNet_io_in_1_bits_header_src = GEN_9;
  assign acqNet_io_in_1_bits_header_dst = GEN_10;
  assign acqNet_io_in_1_bits_payload_addr_block = GEN_11;
  assign acqNet_io_in_1_bits_payload_client_xact_id = GEN_12;
  assign acqNet_io_in_1_bits_payload_addr_beat = GEN_13;
  assign acqNet_io_in_1_bits_payload_is_builtin_type = GEN_14;
  assign acqNet_io_in_1_bits_payload_a_type = GEN_15;
  assign acqNet_io_in_1_bits_payload_union = GEN_16;
  assign acqNet_io_in_1_bits_payload_data = GEN_17;
  assign acqNet_io_in_2_valid = T_13624_valid;
  assign acqNet_io_in_2_bits_header_src = T_13624_bits_header_src;
  assign acqNet_io_in_2_bits_header_dst = T_13624_bits_header_dst;
  assign acqNet_io_in_2_bits_payload_addr_block = T_13624_bits_payload_addr_block;
  assign acqNet_io_in_2_bits_payload_client_xact_id = T_13624_bits_payload_client_xact_id;
  assign acqNet_io_in_2_bits_payload_addr_beat = T_13624_bits_payload_addr_beat;
  assign acqNet_io_in_2_bits_payload_is_builtin_type = T_13624_bits_payload_is_builtin_type;
  assign acqNet_io_in_2_bits_payload_a_type = T_13624_bits_payload_a_type;
  assign acqNet_io_in_2_bits_payload_union = T_13624_bits_payload_union;
  assign acqNet_io_in_2_bits_payload_data = T_13624_bits_payload_data;
  assign acqNet_io_in_3_valid = T_13794_valid;
  assign acqNet_io_in_3_bits_header_src = T_13794_bits_header_src;
  assign acqNet_io_in_3_bits_header_dst = T_13794_bits_header_dst;
  assign acqNet_io_in_3_bits_payload_addr_block = T_13794_bits_payload_addr_block;
  assign acqNet_io_in_3_bits_payload_client_xact_id = T_13794_bits_payload_client_xact_id;
  assign acqNet_io_in_3_bits_payload_addr_beat = T_13794_bits_payload_addr_beat;
  assign acqNet_io_in_3_bits_payload_is_builtin_type = T_13794_bits_payload_is_builtin_type;
  assign acqNet_io_in_3_bits_payload_a_type = T_13794_bits_payload_a_type;
  assign acqNet_io_in_3_bits_payload_union = T_13794_bits_payload_union;
  assign acqNet_io_in_3_bits_payload_data = T_13794_bits_payload_data;
  assign acqNet_io_out_0_ready = T_12724_ready;
  assign acqNet_io_out_1_ready = T_13294_ready;
  assign acqNet_io_out_2_ready = 1'h0;
  assign acqNet_io_out_3_ready = 1'h0;
  assign relNet_clk = clk;
  assign relNet_reset = reset;
  assign relNet_io_in_0_valid = 1'h0;
  assign relNet_io_in_0_bits_header_src = GEN_18;
  assign relNet_io_in_0_bits_header_dst = GEN_19;
  assign relNet_io_in_0_bits_payload_addr_beat = GEN_20;
  assign relNet_io_in_0_bits_payload_addr_block = GEN_21;
  assign relNet_io_in_0_bits_payload_client_xact_id = GEN_22;
  assign relNet_io_in_0_bits_payload_voluntary = GEN_23;
  assign relNet_io_in_0_bits_payload_r_type = GEN_24;
  assign relNet_io_in_0_bits_payload_data = GEN_25;
  assign relNet_io_in_1_valid = 1'h0;
  assign relNet_io_in_1_bits_header_src = GEN_26;
  assign relNet_io_in_1_bits_header_dst = GEN_27;
  assign relNet_io_in_1_bits_payload_addr_beat = GEN_28;
  assign relNet_io_in_1_bits_payload_addr_block = GEN_29;
  assign relNet_io_in_1_bits_payload_client_xact_id = GEN_30;
  assign relNet_io_in_1_bits_payload_voluntary = GEN_31;
  assign relNet_io_in_1_bits_payload_r_type = GEN_32;
  assign relNet_io_in_1_bits_payload_data = GEN_33;
  assign relNet_io_in_2_valid = T_15091_valid;
  assign relNet_io_in_2_bits_header_src = T_15091_bits_header_src;
  assign relNet_io_in_2_bits_header_dst = T_15091_bits_header_dst;
  assign relNet_io_in_2_bits_payload_addr_beat = T_15091_bits_payload_addr_beat;
  assign relNet_io_in_2_bits_payload_addr_block = T_15091_bits_payload_addr_block;
  assign relNet_io_in_2_bits_payload_client_xact_id = T_15091_bits_payload_client_xact_id;
  assign relNet_io_in_2_bits_payload_voluntary = T_15091_bits_payload_voluntary;
  assign relNet_io_in_2_bits_payload_r_type = T_15091_bits_payload_r_type;
  assign relNet_io_in_2_bits_payload_data = T_15091_bits_payload_data;
  assign relNet_io_in_3_valid = T_15256_valid;
  assign relNet_io_in_3_bits_header_src = T_15256_bits_header_src;
  assign relNet_io_in_3_bits_header_dst = T_15256_bits_header_dst;
  assign relNet_io_in_3_bits_payload_addr_beat = T_15256_bits_payload_addr_beat;
  assign relNet_io_in_3_bits_payload_addr_block = T_15256_bits_payload_addr_block;
  assign relNet_io_in_3_bits_payload_client_xact_id = T_15256_bits_payload_client_xact_id;
  assign relNet_io_in_3_bits_payload_voluntary = T_15256_bits_payload_voluntary;
  assign relNet_io_in_3_bits_payload_r_type = T_15256_bits_payload_r_type;
  assign relNet_io_in_3_bits_payload_data = T_15256_bits_payload_data;
  assign relNet_io_out_0_ready = T_14201_ready;
  assign relNet_io_out_1_ready = T_14766_ready;
  assign relNet_io_out_2_ready = 1'h0;
  assign relNet_io_out_3_ready = 1'h0;
  assign prbNet_clk = clk;
  assign prbNet_reset = reset;
  assign prbNet_io_in_0_valid = T_15409_valid;
  assign prbNet_io_in_0_bits_header_src = T_15409_bits_header_src;
  assign prbNet_io_in_0_bits_header_dst = T_15409_bits_header_dst;
  assign prbNet_io_in_0_bits_payload_addr_block = T_15409_bits_payload_addr_block;
  assign prbNet_io_in_0_bits_payload_p_type = T_15409_bits_payload_p_type;
  assign prbNet_io_in_1_valid = T_15554_valid;
  assign prbNet_io_in_1_bits_header_src = T_15554_bits_header_src;
  assign prbNet_io_in_1_bits_header_dst = T_15554_bits_header_dst;
  assign prbNet_io_in_1_bits_payload_addr_block = T_15554_bits_payload_addr_block;
  assign prbNet_io_in_1_bits_payload_p_type = T_15554_bits_payload_p_type;
  assign prbNet_io_in_2_valid = 1'h0;
  assign prbNet_io_in_2_bits_header_src = GEN_34;
  assign prbNet_io_in_2_bits_header_dst = GEN_35;
  assign prbNet_io_in_2_bits_payload_addr_block = GEN_36;
  assign prbNet_io_in_2_bits_payload_p_type = GEN_37;
  assign prbNet_io_in_3_valid = 1'h0;
  assign prbNet_io_in_3_bits_header_src = GEN_38;
  assign prbNet_io_in_3_bits_header_dst = GEN_39;
  assign prbNet_io_in_3_bits_payload_addr_block = GEN_40;
  assign prbNet_io_in_3_bits_payload_p_type = GEN_41;
  assign prbNet_io_out_0_ready = 1'h0;
  assign prbNet_io_out_1_ready = 1'h0;
  assign prbNet_io_out_2_ready = T_15939_ready;
  assign prbNet_io_out_3_ready = T_16484_ready;
  assign gntNet_clk = clk;
  assign gntNet_reset = reset;
  assign gntNet_io_in_0_valid = T_16801_valid;
  assign gntNet_io_in_0_bits_header_src = T_16801_bits_header_src;
  assign gntNet_io_in_0_bits_header_dst = T_16801_bits_header_dst;
  assign gntNet_io_in_0_bits_payload_addr_beat = T_16801_bits_payload_addr_beat;
  assign gntNet_io_in_0_bits_payload_client_xact_id = T_16801_bits_payload_client_xact_id;
  assign gntNet_io_in_0_bits_payload_manager_xact_id = T_16801_bits_payload_manager_xact_id;
  assign gntNet_io_in_0_bits_payload_is_builtin_type = T_16801_bits_payload_is_builtin_type;
  assign gntNet_io_in_0_bits_payload_g_type = T_16801_bits_payload_g_type;
  assign gntNet_io_in_0_bits_payload_data = T_16801_bits_payload_data;
  assign gntNet_io_in_1_valid = T_16966_valid;
  assign gntNet_io_in_1_bits_header_src = T_16966_bits_header_src;
  assign gntNet_io_in_1_bits_header_dst = T_16966_bits_header_dst;
  assign gntNet_io_in_1_bits_payload_addr_beat = T_16966_bits_payload_addr_beat;
  assign gntNet_io_in_1_bits_payload_client_xact_id = T_16966_bits_payload_client_xact_id;
  assign gntNet_io_in_1_bits_payload_manager_xact_id = T_16966_bits_payload_manager_xact_id;
  assign gntNet_io_in_1_bits_payload_is_builtin_type = T_16966_bits_payload_is_builtin_type;
  assign gntNet_io_in_1_bits_payload_g_type = T_16966_bits_payload_g_type;
  assign gntNet_io_in_1_bits_payload_data = T_16966_bits_payload_data;
  assign gntNet_io_in_2_valid = 1'h0;
  assign gntNet_io_in_2_bits_header_src = GEN_42;
  assign gntNet_io_in_2_bits_header_dst = GEN_43;
  assign gntNet_io_in_2_bits_payload_addr_beat = GEN_44;
  assign gntNet_io_in_2_bits_payload_client_xact_id = GEN_45;
  assign gntNet_io_in_2_bits_payload_manager_xact_id = GEN_46;
  assign gntNet_io_in_2_bits_payload_is_builtin_type = GEN_47;
  assign gntNet_io_in_2_bits_payload_g_type = GEN_48;
  assign gntNet_io_in_2_bits_payload_data = GEN_49;
  assign gntNet_io_in_3_valid = 1'h0;
  assign gntNet_io_in_3_bits_header_src = GEN_50;
  assign gntNet_io_in_3_bits_header_dst = GEN_51;
  assign gntNet_io_in_3_bits_payload_addr_beat = GEN_52;
  assign gntNet_io_in_3_bits_payload_client_xact_id = GEN_53;
  assign gntNet_io_in_3_bits_payload_manager_xact_id = GEN_54;
  assign gntNet_io_in_3_bits_payload_is_builtin_type = GEN_55;
  assign gntNet_io_in_3_bits_payload_g_type = GEN_56;
  assign gntNet_io_in_3_bits_payload_data = GEN_57;
  assign gntNet_io_out_0_ready = 1'h0;
  assign gntNet_io_out_1_ready = 1'h0;
  assign gntNet_io_out_2_ready = T_17371_ready;
  assign gntNet_io_out_3_ready = T_17936_ready;
  assign ackNet_clk = clk;
  assign ackNet_reset = reset;
  assign ackNet_io_in_0_valid = 1'h0;
  assign ackNet_io_in_0_bits_header_src = GEN_58;
  assign ackNet_io_in_0_bits_header_dst = GEN_59;
  assign ackNet_io_in_0_bits_payload_manager_xact_id = GEN_60;
  assign ackNet_io_in_1_valid = 1'h0;
  assign ackNet_io_in_1_bits_header_src = GEN_61;
  assign ackNet_io_in_1_bits_header_dst = GEN_62;
  assign ackNet_io_in_1_bits_payload_manager_xact_id = GEN_63;
  assign ackNet_io_in_2_valid = T_19326_valid;
  assign ackNet_io_in_2_bits_header_src = T_19326_bits_header_src;
  assign ackNet_io_in_2_bits_header_dst = T_19326_bits_header_dst;
  assign ackNet_io_in_2_bits_payload_manager_xact_id = T_19326_bits_payload_manager_xact_id;
  assign ackNet_io_in_3_valid = T_19466_valid;
  assign ackNet_io_in_3_bits_header_src = T_19466_bits_header_src;
  assign ackNet_io_in_3_bits_header_dst = T_19466_bits_header_dst;
  assign ackNet_io_in_3_bits_payload_manager_xact_id = T_19466_bits_payload_manager_xact_id;
  assign ackNet_io_out_0_ready = T_18486_ready;
  assign ackNet_io_out_1_ready = T_19026_ready;
  assign ackNet_io_out_2_ready = 1'h0;
  assign ackNet_io_out_3_ready = 1'h0;
  assign T_12724_ready = TileLinkEnqueuer_2_1_io_client_acquire_ready;
  assign T_12724_valid = acqNet_io_out_0_valid;
  assign T_12724_bits_header_src = T_12953;
  assign T_12724_bits_header_dst = acqNet_io_out_0_bits_header_dst;
  assign T_12724_bits_payload_addr_block = acqNet_io_out_0_bits_payload_addr_block;
  assign T_12724_bits_payload_client_xact_id = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T_12724_bits_payload_addr_beat = acqNet_io_out_0_bits_payload_addr_beat;
  assign T_12724_bits_payload_is_builtin_type = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T_12724_bits_payload_a_type = acqNet_io_out_0_bits_payload_a_type;
  assign T_12724_bits_payload_union = acqNet_io_out_0_bits_payload_union;
  assign T_12724_bits_payload_data = acqNet_io_out_0_bits_payload_data;
  assign T_12952 = acqNet_io_out_0_bits_header_src - 2'h2;
  assign T_12953 = T_12952[1:0];
  assign T_13294_ready = TileLinkEnqueuer_3_1_io_client_acquire_ready;
  assign T_13294_valid = acqNet_io_out_1_valid;
  assign T_13294_bits_header_src = T_13523;
  assign T_13294_bits_header_dst = acqNet_io_out_1_bits_header_dst;
  assign T_13294_bits_payload_addr_block = acqNet_io_out_1_bits_payload_addr_block;
  assign T_13294_bits_payload_client_xact_id = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T_13294_bits_payload_addr_beat = acqNet_io_out_1_bits_payload_addr_beat;
  assign T_13294_bits_payload_is_builtin_type = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T_13294_bits_payload_a_type = acqNet_io_out_1_bits_payload_a_type;
  assign T_13294_bits_payload_union = acqNet_io_out_1_bits_payload_union;
  assign T_13294_bits_payload_data = acqNet_io_out_1_bits_payload_data;
  assign T_13522 = acqNet_io_out_1_bits_header_src - 2'h2;
  assign T_13523 = T_13522[1:0];
  assign T_13624_ready = acqNet_io_in_2_ready;
  assign T_13624_valid = TileLinkEnqueuer_4_io_manager_acquire_valid;
  assign T_13624_bits_header_src = T_13693;
  assign T_13624_bits_header_dst = TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  assign T_13624_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  assign T_13624_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13624_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  assign T_13624_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13624_bits_payload_a_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  assign T_13624_bits_payload_union = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  assign T_13624_bits_payload_data = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  assign T_13692 = TileLinkEnqueuer_4_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13693 = T_13692[1:0];
  assign T_13794_ready = acqNet_io_in_3_ready;
  assign T_13794_valid = TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  assign T_13794_bits_header_src = T_13863;
  assign T_13794_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  assign T_13794_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  assign T_13794_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13794_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  assign T_13794_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13794_bits_payload_a_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  assign T_13794_bits_payload_union = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  assign T_13794_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  assign T_13862 = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13863 = T_13862[1:0];
  assign T_14201_ready = TileLinkEnqueuer_2_1_io_client_release_ready;
  assign T_14201_valid = relNet_io_out_0_valid;
  assign T_14201_bits_header_src = T_14428;
  assign T_14201_bits_header_dst = relNet_io_out_0_bits_header_dst;
  assign T_14201_bits_payload_addr_beat = relNet_io_out_0_bits_payload_addr_beat;
  assign T_14201_bits_payload_addr_block = relNet_io_out_0_bits_payload_addr_block;
  assign T_14201_bits_payload_client_xact_id = relNet_io_out_0_bits_payload_client_xact_id;
  assign T_14201_bits_payload_voluntary = relNet_io_out_0_bits_payload_voluntary;
  assign T_14201_bits_payload_r_type = relNet_io_out_0_bits_payload_r_type;
  assign T_14201_bits_payload_data = relNet_io_out_0_bits_payload_data;
  assign T_14427 = relNet_io_out_0_bits_header_src - 2'h2;
  assign T_14428 = T_14427[1:0];
  assign T_14766_ready = TileLinkEnqueuer_3_1_io_client_release_ready;
  assign T_14766_valid = relNet_io_out_1_valid;
  assign T_14766_bits_header_src = T_14993;
  assign T_14766_bits_header_dst = relNet_io_out_1_bits_header_dst;
  assign T_14766_bits_payload_addr_beat = relNet_io_out_1_bits_payload_addr_beat;
  assign T_14766_bits_payload_addr_block = relNet_io_out_1_bits_payload_addr_block;
  assign T_14766_bits_payload_client_xact_id = relNet_io_out_1_bits_payload_client_xact_id;
  assign T_14766_bits_payload_voluntary = relNet_io_out_1_bits_payload_voluntary;
  assign T_14766_bits_payload_r_type = relNet_io_out_1_bits_payload_r_type;
  assign T_14766_bits_payload_data = relNet_io_out_1_bits_payload_data;
  assign T_14992 = relNet_io_out_1_bits_header_src - 2'h2;
  assign T_14993 = T_14992[1:0];
  assign T_15091_ready = relNet_io_in_2_ready;
  assign T_15091_valid = TileLinkEnqueuer_4_io_manager_release_valid;
  assign T_15091_bits_header_src = T_15158;
  assign T_15091_bits_header_dst = TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  assign T_15091_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  assign T_15091_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  assign T_15091_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  assign T_15091_bits_payload_voluntary = TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  assign T_15091_bits_payload_r_type = TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  assign T_15091_bits_payload_data = TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  assign T_15157 = TileLinkEnqueuer_4_io_manager_release_bits_header_src + 2'h2;
  assign T_15158 = T_15157[1:0];
  assign T_15256_ready = relNet_io_in_3_ready;
  assign T_15256_valid = TileLinkEnqueuer_1_1_io_manager_release_valid;
  assign T_15256_bits_header_src = T_15323;
  assign T_15256_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  assign T_15256_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  assign T_15256_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  assign T_15256_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  assign T_15256_bits_payload_voluntary = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  assign T_15256_bits_payload_r_type = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  assign T_15256_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  assign T_15322 = TileLinkEnqueuer_1_1_io_manager_release_bits_header_src + 2'h2;
  assign T_15323 = T_15322[1:0];
  assign T_15409_ready = prbNet_io_in_0_ready;
  assign T_15409_valid = TileLinkEnqueuer_2_1_io_client_probe_valid;
  assign T_15409_bits_header_src = TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  assign T_15409_bits_header_dst = T_15468;
  assign T_15409_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  assign T_15409_bits_payload_p_type = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  assign T_15467 = TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15468 = T_15467[1:0];
  assign T_15554_ready = prbNet_io_in_1_ready;
  assign T_15554_valid = TileLinkEnqueuer_3_1_io_client_probe_valid;
  assign T_15554_bits_header_src = TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  assign T_15554_bits_header_dst = T_15613;
  assign T_15554_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  assign T_15554_bits_payload_p_type = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  assign T_15612 = TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15613 = T_15612[1:0];
  assign T_15939_ready = TileLinkEnqueuer_4_io_manager_probe_ready;
  assign T_15939_valid = prbNet_io_out_2_valid;
  assign T_15939_bits_header_src = prbNet_io_out_2_bits_header_src;
  assign T_15939_bits_header_dst = T_16158;
  assign T_15939_bits_payload_addr_block = prbNet_io_out_2_bits_payload_addr_block;
  assign T_15939_bits_payload_p_type = prbNet_io_out_2_bits_payload_p_type;
  assign T_16157 = prbNet_io_out_2_bits_header_dst - 2'h2;
  assign T_16158 = T_16157[1:0];
  assign T_16484_ready = TileLinkEnqueuer_1_1_io_manager_probe_ready;
  assign T_16484_valid = prbNet_io_out_3_valid;
  assign T_16484_bits_header_src = prbNet_io_out_3_bits_header_src;
  assign T_16484_bits_header_dst = T_16703;
  assign T_16484_bits_payload_addr_block = prbNet_io_out_3_bits_payload_addr_block;
  assign T_16484_bits_payload_p_type = prbNet_io_out_3_bits_payload_p_type;
  assign T_16702 = prbNet_io_out_3_bits_header_dst - 2'h2;
  assign T_16703 = T_16702[1:0];
  assign T_16801_ready = gntNet_io_in_0_ready;
  assign T_16801_valid = TileLinkEnqueuer_2_1_io_client_grant_valid;
  assign T_16801_bits_header_src = TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  assign T_16801_bits_header_dst = T_16868;
  assign T_16801_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  assign T_16801_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16801_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16801_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16801_bits_payload_g_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  assign T_16801_bits_payload_data = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  assign T_16867 = TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_16868 = T_16867[1:0];
  assign T_16966_ready = gntNet_io_in_1_ready;
  assign T_16966_valid = TileLinkEnqueuer_3_1_io_client_grant_valid;
  assign T_16966_bits_header_src = TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  assign T_16966_bits_header_dst = T_17033;
  assign T_16966_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  assign T_16966_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16966_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16966_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16966_bits_payload_g_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  assign T_16966_bits_payload_data = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  assign T_17032 = TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_17033 = T_17032[1:0];
  assign T_17371_ready = TileLinkEnqueuer_4_io_manager_grant_ready;
  assign T_17371_valid = gntNet_io_out_2_valid;
  assign T_17371_bits_header_src = gntNet_io_out_2_bits_header_src;
  assign T_17371_bits_header_dst = T_17598;
  assign T_17371_bits_payload_addr_beat = gntNet_io_out_2_bits_payload_addr_beat;
  assign T_17371_bits_payload_client_xact_id = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T_17371_bits_payload_manager_xact_id = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T_17371_bits_payload_is_builtin_type = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T_17371_bits_payload_g_type = gntNet_io_out_2_bits_payload_g_type;
  assign T_17371_bits_payload_data = gntNet_io_out_2_bits_payload_data;
  assign T_17597 = gntNet_io_out_2_bits_header_dst - 2'h2;
  assign T_17598 = T_17597[1:0];
  assign T_17936_ready = TileLinkEnqueuer_1_1_io_manager_grant_ready;
  assign T_17936_valid = gntNet_io_out_3_valid;
  assign T_17936_bits_header_src = gntNet_io_out_3_bits_header_src;
  assign T_17936_bits_header_dst = T_18163;
  assign T_17936_bits_payload_addr_beat = gntNet_io_out_3_bits_payload_addr_beat;
  assign T_17936_bits_payload_client_xact_id = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T_17936_bits_payload_manager_xact_id = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T_17936_bits_payload_is_builtin_type = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T_17936_bits_payload_g_type = gntNet_io_out_3_bits_payload_g_type;
  assign T_17936_bits_payload_data = gntNet_io_out_3_bits_payload_data;
  assign T_18162 = gntNet_io_out_3_bits_header_dst - 2'h2;
  assign T_18163 = T_18162[1:0];
  assign T_18486_ready = TileLinkEnqueuer_2_1_io_client_finish_ready;
  assign T_18486_valid = ackNet_io_out_0_valid;
  assign T_18486_bits_header_src = T_18703;
  assign T_18486_bits_header_dst = ackNet_io_out_0_bits_header_dst;
  assign T_18486_bits_payload_manager_xact_id = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T_18702 = ackNet_io_out_0_bits_header_src - 2'h2;
  assign T_18703 = T_18702[1:0];
  assign T_19026_ready = TileLinkEnqueuer_3_1_io_client_finish_ready;
  assign T_19026_valid = ackNet_io_out_1_valid;
  assign T_19026_bits_header_src = T_19243;
  assign T_19026_bits_header_dst = ackNet_io_out_1_bits_header_dst;
  assign T_19026_bits_payload_manager_xact_id = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T_19242 = ackNet_io_out_1_bits_header_src - 2'h2;
  assign T_19243 = T_19242[1:0];
  assign T_19326_ready = ackNet_io_in_2_ready;
  assign T_19326_valid = TileLinkEnqueuer_4_io_manager_finish_valid;
  assign T_19326_bits_header_src = T_19383;
  assign T_19326_bits_header_dst = TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  assign T_19326_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19382 = TileLinkEnqueuer_4_io_manager_finish_bits_header_src + 2'h2;
  assign T_19383 = T_19382[1:0];
  assign T_19466_ready = ackNet_io_in_3_ready;
  assign T_19466_valid = TileLinkEnqueuer_1_1_io_manager_finish_valid;
  assign T_19466_bits_header_src = T_19523;
  assign T_19466_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  assign T_19466_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19522 = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src + 2'h2;
  assign T_19523 = T_19522[1:0];
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_64[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_65[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_66[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_67[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_68[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_5 = GEN_69[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_6 = GEN_70[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_7 = GEN_71[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_8 = GEN_72[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_73[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_74[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_75[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_12 = GEN_76[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_77[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_78[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_80[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_81[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_18 = GEN_82[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_19 = GEN_83[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_20 = GEN_84[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_21 = GEN_85[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_22 = GEN_86[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_23 = GEN_87[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_24 = GEN_88[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_25 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_26 = GEN_90[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_27 = GEN_91[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_28 = GEN_92[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_93[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_94[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_95[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_32 = GEN_96[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_33 = GEN_97[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_34 = GEN_98[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_35 = GEN_99[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_36 = GEN_100[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_37 = GEN_101[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_38 = GEN_102[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_39 = GEN_103[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_40 = GEN_104[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_41 = GEN_105[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_42 = GEN_106[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_43 = GEN_107[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_44 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_45 = GEN_109[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_46 = GEN_110[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_47 = GEN_111[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_48 = GEN_112[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_49 = GEN_113[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_50 = GEN_114[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_51 = GEN_115[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_52 = GEN_116[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_53 = GEN_117[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_54 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_55 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_56 = GEN_120[3:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_57 = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_58 = GEN_122[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_123[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_124[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_126[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_127[2:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_64 = {1{$random}};
  GEN_65 = {1{$random}};
  GEN_66 = {1{$random}};
  GEN_67 = {1{$random}};
  GEN_68 = {1{$random}};
  GEN_69 = {1{$random}};
  GEN_70 = {1{$random}};
  GEN_71 = {1{$random}};
  GEN_72 = {2{$random}};
  GEN_73 = {1{$random}};
  GEN_74 = {1{$random}};
  GEN_75 = {1{$random}};
  GEN_76 = {1{$random}};
  GEN_77 = {1{$random}};
  GEN_78 = {1{$random}};
  GEN_79 = {1{$random}};
  GEN_80 = {1{$random}};
  GEN_81 = {2{$random}};
  GEN_82 = {1{$random}};
  GEN_83 = {1{$random}};
  GEN_84 = {1{$random}};
  GEN_85 = {1{$random}};
  GEN_86 = {1{$random}};
  GEN_87 = {1{$random}};
  GEN_88 = {1{$random}};
  GEN_89 = {2{$random}};
  GEN_90 = {1{$random}};
  GEN_91 = {1{$random}};
  GEN_92 = {1{$random}};
  GEN_93 = {1{$random}};
  GEN_94 = {1{$random}};
  GEN_95 = {1{$random}};
  GEN_96 = {1{$random}};
  GEN_97 = {2{$random}};
  GEN_98 = {1{$random}};
  GEN_99 = {1{$random}};
  GEN_100 = {1{$random}};
  GEN_101 = {1{$random}};
  GEN_102 = {1{$random}};
  GEN_103 = {1{$random}};
  GEN_104 = {1{$random}};
  GEN_105 = {1{$random}};
  GEN_106 = {1{$random}};
  GEN_107 = {1{$random}};
  GEN_108 = {1{$random}};
  GEN_109 = {1{$random}};
  GEN_110 = {1{$random}};
  GEN_111 = {1{$random}};
  GEN_112 = {1{$random}};
  GEN_113 = {2{$random}};
  GEN_114 = {1{$random}};
  GEN_115 = {1{$random}};
  GEN_116 = {1{$random}};
  GEN_117 = {1{$random}};
  GEN_118 = {1{$random}};
  GEN_119 = {1{$random}};
  GEN_120 = {1{$random}};
  GEN_121 = {2{$random}};
  GEN_122 = {1{$random}};
  GEN_123 = {1{$random}};
  GEN_124 = {1{$random}};
  GEN_125 = {1{$random}};
  GEN_126 = {1{$random}};
  GEN_127 = {1{$random}};
  end
`endif
endmodule
module BufferedBroadcastVoluntaryReleaseTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_69;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_70;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_71;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_72;
  reg [1:0] xact_vol_ir_client_xact_id;
  reg [31:0] GEN_73;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_74;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  reg  pending_orel_send;
  reg [31:0] GEN_75;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_76;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_78;
  wire  T_79;
  wire  scoreboard_2;
  reg  sending_orel;
  reg [31:0] GEN_77;
  wire  T_103_sharers;
  wire [1:0] T_149_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1519;
  wire  T_1520;
  wire  T_1521;
  wire  T_1522;
  wire  T_1524;
  wire  T_1525;
  wire  T_1527;
  wire  T_1528;
  wire  T_1530;
  wire [63:0] T_1544_0;
  wire [63:0] T_1544_1;
  wire [63:0] T_1544_2;
  wire [63:0] T_1544_3;
  wire [63:0] T_1544_4;
  wire [63:0] T_1544_5;
  wire [63:0] T_1544_6;
  wire [63:0] T_1544_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_78;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_79;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_80;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_81;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_82;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_83;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_84;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_85;
  wire  T_1552;
  wire  T_1553;
  wire  T_1554;
  wire  T_1556;
  wire  T_1557;
  wire  T_1559;
  wire  T_1560;
  wire  T_1568;
  wire  T_1572;
  wire  T_1573;
  wire  T_1578;
  wire  T_1580;
  wire  T_1581;
  wire  T_1582;
  wire  T_1583;
  wire  T_1584;
  wire  T_1586;
  reg [2:0] T_1588;
  reg [31:0] GEN_86;
  wire  T_1590;
  wire [3:0] T_1592;
  wire [2:0] T_1593;
  wire [2:0] GEN_2;
  wire  T_1594;
  wire [2:0] T_1595;
  wire  T_1596;
  wire  T_1597;
  wire  T_1600;
  wire  T_1601;
  wire  T_1602;
  wire  T_1603;
  wire [2:0] T_1611_0;
  wire [3:0] GEN_57;
  wire  T_1613;
  wire  T_1615;
  wire  T_1617;
  reg [2:0] T_1619;
  reg [31:0] GEN_87;
  wire  T_1621;
  wire [3:0] T_1623;
  wire [2:0] T_1624;
  wire [2:0] GEN_3;
  wire  T_1625;
  wire [2:0] T_1626;
  wire  T_1627;
  reg  T_1629;
  reg [31:0] GEN_88;
  wire  T_1631;
  wire  T_1632;
  wire [1:0] T_1634;
  wire  T_1635;
  wire  GEN_4;
  wire  T_1637;
  wire  T_1638;
  wire [1:0] T_1640;
  wire  T_1641;
  wire  GEN_5;
  wire  T_1643;
  wire  T_1645;
  wire  T_1646;
  wire [25:0] GEN_6;
  wire [7:0] GEN_7;
  wire [3:0] GEN_8;
  wire  T_1654;
  wire  T_1656;
  wire  T_1657;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1670;
  wire  T_1672;
  wire  T_1673;
  wire [2:0] GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_11;
  wire  T_1687;
  wire [7:0] T_1691;
  wire [7:0] T_1692;
  wire [7:0] T_1694;
  wire [7:0] T_1695;
  wire [7:0] T_1696;
  wire [7:0] T_1698;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [1:0] GEN_14;
  wire [7:0] GEN_15;
  wire  T_1700;
  wire [7:0] T_1717;
  wire [7:0] GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  wire [1:0] GEN_19;
  wire [7:0] GEN_20;
  wire  T_1718;
  wire  T_1719;
  wire  T_1720;
  wire  T_1721;
  wire  T_1722;
  wire  T_1723;
  wire  T_1724;
  wire  T_1725;
  wire  T_1728;
  wire  T_1730;
  wire  T_1731;
  wire [2:0] T_1763_addr_beat;
  wire [25:0] T_1763_addr_block;
  wire [1:0] T_1763_client_xact_id;
  wire  T_1763_voluntary;
  wire [2:0] T_1763_r_type;
  wire [63:0] T_1763_data;
  wire  T_1763_client_id;
  wire [2:0] T_1824_addr_beat;
  wire [1:0] T_1824_client_xact_id;
  wire [2:0] T_1824_manager_xact_id;
  wire  T_1824_is_builtin_type;
  wire [3:0] T_1824_g_type;
  wire [63:0] T_1824_data;
  wire  T_1824_client_id;
  wire  T_1861;
  wire [63:0] GEN_0;
  wire [63:0] GEN_21;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [1:0] T_1893_state;
  wire  T_1922;
  wire [7:0] T_1938;
  wire [7:0] T_1939;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1954;
  wire [7:0] T_1955;
  wire [7:0] T_1956;
  wire [7:0] T_1957;
  wire [7:0] GEN_38;
  wire  GEN_39;
  wire  T_1968;
  wire  T_1970;
  wire  T_1971;
  wire  GEN_40;
  wire  T_1983;
  wire  T_1984;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_1993;
  wire  T_2001;
  reg [2:0] T_2003;
  reg [31:0] GEN_89;
  wire  T_2005;
  wire [3:0] T_2007;
  wire [2:0] T_2008;
  wire [2:0] GEN_44;
  wire  T_2009;
  wire [2:0] T_2010;
  wire  T_2011;
  wire  T_2012;
  wire  T_2014;
  wire  T_2015;
  wire  T_2016;
  wire [2:0] T_2024_0;
  wire [3:0] GEN_58;
  wire  T_2026;
  wire  T_2028;
  wire  T_2030;
  reg [2:0] T_2032;
  reg [31:0] GEN_90;
  wire  T_2034;
  wire [3:0] T_2036;
  wire [2:0] T_2037;
  wire [2:0] GEN_45;
  wire  T_2038;
  wire [2:0] T_2039;
  wire  T_2040;
  reg  T_2042;
  reg [31:0] GEN_91;
  wire  T_2044;
  wire  T_2045;
  wire [1:0] T_2047;
  wire  T_2048;
  wire  GEN_46;
  wire  T_2050;
  wire  T_2051;
  wire [1:0] T_2053;
  wire  T_2054;
  wire  GEN_47;
  wire  T_2056;
  wire [7:0] T_2065;
  wire  T_2066;
  wire  T_2067;
  wire  T_2068;
  wire  T_2082;
  wire [2:0] T_2083;
  wire [2:0] T_2119_addr_beat;
  wire [25:0] T_2119_addr_block;
  wire [2:0] T_2119_client_xact_id;
  wire  T_2119_voluntary;
  wire [2:0] T_2119_r_type;
  wire [63:0] T_2119_data;
  wire [63:0] GEN_1;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire  T_2149;
  wire  T_2150;
  wire  T_2151;
  wire  T_2153;
  wire  T_2155;
  wire [3:0] GEN_56;
  wire [25:0] GEN_29;
  reg [31:0] GEN_92;
  wire [1:0] GEN_55;
  reg [31:0] GEN_93;
  wire  GEN_59;
  reg [31:0] GEN_94;
  wire [25:0] GEN_60;
  reg [31:0] GEN_95;
  wire [2:0] GEN_61;
  reg [31:0] GEN_96;
  wire [2:0] GEN_62;
  reg [31:0] GEN_97;
  wire  GEN_63;
  reg [31:0] GEN_98;
  wire [2:0] GEN_64;
  reg [31:0] GEN_99;
  wire [10:0] GEN_65;
  reg [31:0] GEN_100;
  wire [63:0] GEN_66;
  reg [63:0] GEN_101;
  wire  GEN_67;
  reg [31:0] GEN_102;
  wire  GEN_68;
  reg [31:0] GEN_103;
  assign io_inner_acquire_ready = 1'h0;
  assign io_inner_grant_valid = T_1731;
  assign io_inner_grant_bits_addr_beat = T_1824_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1824_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1824_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1824_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1824_g_type;
  assign io_inner_grant_bits_data = T_1824_data;
  assign io_inner_grant_bits_client_id = T_1824_client_id;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_29;
  assign io_inner_probe_bits_p_type = GEN_55;
  assign io_inner_probe_bits_client_id = GEN_59;
  assign io_inner_release_ready = T_1861;
  assign io_outer_acquire_valid = 1'h0;
  assign io_outer_acquire_bits_addr_block = GEN_60;
  assign io_outer_acquire_bits_client_xact_id = GEN_61;
  assign io_outer_acquire_bits_addr_beat = GEN_62;
  assign io_outer_acquire_bits_is_builtin_type = GEN_63;
  assign io_outer_acquire_bits_a_type = GEN_64;
  assign io_outer_acquire_bits_union = GEN_65;
  assign io_outer_acquire_bits_data = GEN_66;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2068;
  assign io_outer_release_bits_addr_beat = T_2119_addr_beat;
  assign io_outer_release_bits_addr_block = T_2119_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2119_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2119_voluntary;
  assign io_outer_release_bits_r_type = T_2119_r_type;
  assign io_outer_release_bits_data = T_2119_data;
  assign io_outer_grant_ready = vol_ognt_counter_pending;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_67;
  assign io_outer_finish_bits_manager_id = GEN_68;
  assign io_alloc_iacq_matches = T_1554;
  assign io_alloc_iacq_can = 1'h0;
  assign io_alloc_irel_matches = T_1557;
  assign io_alloc_irel_can = T_1519;
  assign io_alloc_oprb_matches = T_1560;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1519;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_2153;
  assign vol_ignt_counter_pending = T_1643;
  assign vol_ignt_counter_up_idx = T_1595;
  assign vol_ignt_counter_up_done = T_1596;
  assign vol_ignt_counter_down_idx = T_1626;
  assign vol_ignt_counter_down_done = T_1627;
  assign vol_ognt_counter_pending = T_2056;
  assign vol_ognt_counter_up_idx = T_2010;
  assign vol_ognt_counter_up_done = T_2011;
  assign vol_ognt_counter_down_idx = T_2039;
  assign vol_ognt_counter_down_done = T_2040;
  assign T_78 = pending_orel_data != 8'h0;
  assign T_79 = pending_orel_send | T_78;
  assign scoreboard_2 = T_79 | vol_ognt_counter_pending;
  assign T_103_sharers = 1'h0;
  assign T_149_state = 2'h0;
  assign coh_inner_sharers = T_103_sharers;
  assign coh_outer_state = T_149_state;
  assign T_1519 = state == 4'h0;
  assign T_1520 = io_inner_release_ready & io_inner_release_valid;
  assign T_1521 = T_1519 & T_1520;
  assign T_1522 = T_1521 & io_alloc_irel_should;
  assign T_1524 = io_inner_release_bits_voluntary == 1'h0;
  assign T_1525 = T_1522 & T_1524;
  assign T_1527 = T_1525 == 1'h0;
  assign T_1528 = T_1527 | reset;
  assign T_1530 = T_1528 == 1'h0;
  assign T_1544_0 = 64'h0;
  assign T_1544_1 = 64'h0;
  assign T_1544_2 = 64'h0;
  assign T_1544_3 = 64'h0;
  assign T_1544_4 = 64'h0;
  assign T_1544_5 = 64'h0;
  assign T_1544_6 = 64'h0;
  assign T_1544_7 = 64'h0;
  assign T_1552 = state != 4'h0;
  assign T_1553 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1554 = T_1552 & T_1553;
  assign T_1556 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1557 = T_1552 & T_1556;
  assign T_1559 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1560 = T_1552 & T_1559;
  assign T_1568 = scoreboard_2 | vol_ognt_counter_pending;
  assign T_1572 = T_1519 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_1573 = T_1572 & io_inner_release_bits_voluntary;
  assign T_1578 = T_1520 & T_1573;
  assign T_1580 = io_inner_release_bits_r_type == 3'h0;
  assign T_1581 = io_inner_release_bits_r_type == 3'h1;
  assign T_1582 = io_inner_release_bits_r_type == 3'h2;
  assign T_1583 = T_1580 | T_1581;
  assign T_1584 = T_1583 | T_1582;
  assign T_1586 = T_1578 & T_1584;
  assign T_1590 = T_1588 == 3'h7;
  assign T_1592 = T_1588 + 3'h1;
  assign T_1593 = T_1592[2:0];
  assign GEN_2 = T_1586 ? T_1593 : T_1588;
  assign T_1594 = T_1586 & T_1590;
  assign T_1595 = T_1584 ? T_1588 : 3'h0;
  assign T_1596 = T_1584 ? T_1594 : T_1578;
  assign T_1597 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1600 = io_inner_grant_bits_g_type == 4'h0;
  assign T_1601 = io_inner_grant_bits_is_builtin_type & T_1600;
  assign T_1602 = T_1552 & T_1601;
  assign T_1603 = T_1597 & T_1602;
  assign T_1611_0 = 3'h5;
  assign GEN_57 = {{1'd0}, T_1611_0};
  assign T_1613 = io_inner_grant_bits_g_type == GEN_57;
  assign T_1615 = io_inner_grant_bits_is_builtin_type ? T_1613 : T_1600;
  assign T_1617 = T_1603 & T_1615;
  assign T_1621 = T_1619 == 3'h7;
  assign T_1623 = T_1619 + 3'h1;
  assign T_1624 = T_1623[2:0];
  assign GEN_3 = T_1617 ? T_1624 : T_1619;
  assign T_1625 = T_1617 & T_1621;
  assign T_1626 = T_1615 ? T_1619 : 3'h0;
  assign T_1627 = T_1615 ? T_1625 : T_1603;
  assign T_1631 = T_1627 == 1'h0;
  assign T_1632 = T_1596 & T_1631;
  assign T_1634 = T_1629 + 1'h1;
  assign T_1635 = T_1634[0:0];
  assign GEN_4 = T_1632 ? T_1635 : T_1629;
  assign T_1637 = T_1596 == 1'h0;
  assign T_1638 = T_1627 & T_1637;
  assign T_1640 = T_1629 - 1'h1;
  assign T_1641 = T_1640[0:0];
  assign GEN_5 = T_1638 ? T_1641 : GEN_4;
  assign T_1643 = T_1629 > 1'h0;
  assign T_1645 = T_1519 & io_alloc_irel_should;
  assign T_1646 = T_1645 & io_inner_release_valid;
  assign GEN_6 = T_1646 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign GEN_7 = T_1646 ? 8'hff : pending_irel_data;
  assign GEN_8 = T_1646 ? 4'h7 : state;
  assign T_1654 = T_1556 & io_inner_release_bits_voluntary;
  assign T_1656 = pending_irel_data != 8'h0;
  assign T_1657 = T_1654 & T_1656;
  assign T_1659 = T_1657 & io_inner_release_valid;
  assign T_1660 = T_1646 | T_1659;
  assign T_1661 = T_1660 & io_inner_release_ready;
  assign T_1670 = T_1584 == 1'h0;
  assign T_1672 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_1673 = T_1670 | T_1672;
  assign GEN_9 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_10 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_11 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_1687 = T_1520 & T_1584;
  assign T_1691 = T_1687 ? 8'hff : 8'h0;
  assign T_1692 = ~ T_1691;
  assign T_1694 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_1695 = ~ T_1694;
  assign T_1696 = T_1692 | T_1695;
  assign T_1698 = T_1584 ? T_1696 : 8'h0;
  assign GEN_12 = T_1673 ? GEN_9 : xact_vol_ir_r_type;
  assign GEN_13 = T_1673 ? GEN_10 : xact_vol_ir_src;
  assign GEN_14 = T_1673 ? GEN_11 : xact_vol_ir_client_xact_id;
  assign GEN_15 = T_1673 ? T_1698 : GEN_7;
  assign T_1700 = T_1673 == 1'h0;
  assign T_1717 = pending_irel_data & T_1696;
  assign GEN_16 = T_1700 ? T_1717 : GEN_15;
  assign GEN_17 = T_1661 ? GEN_12 : xact_vol_ir_r_type;
  assign GEN_18 = T_1661 ? GEN_13 : xact_vol_ir_src;
  assign GEN_19 = T_1661 ? GEN_14 : xact_vol_ir_client_xact_id;
  assign GEN_20 = T_1661 ? GEN_16 : GEN_7;
  assign T_1718 = state == 4'h3;
  assign T_1719 = state == 4'h4;
  assign T_1720 = state == 4'h5;
  assign T_1721 = state == 4'h7;
  assign T_1722 = T_1718 | T_1719;
  assign T_1723 = T_1722 | T_1720;
  assign T_1724 = T_1723 | T_1721;
  assign T_1725 = T_1724 & vol_ignt_counter_pending;
  assign T_1728 = T_1656 | T_1568;
  assign T_1730 = T_1728 == 1'h0;
  assign T_1731 = T_1725 & T_1730;
  assign T_1763_addr_beat = 3'h0;
  assign T_1763_addr_block = xact_addr_block;
  assign T_1763_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_1763_voluntary = 1'h1;
  assign T_1763_r_type = xact_vol_ir_r_type;
  assign T_1763_data = 64'h0;
  assign T_1763_client_id = xact_vol_ir_src;
  assign T_1824_addr_beat = 3'h0;
  assign T_1824_client_xact_id = T_1763_client_xact_id;
  assign T_1824_manager_xact_id = 3'h0;
  assign T_1824_is_builtin_type = 1'h1;
  assign T_1824_g_type = 4'h0;
  assign T_1824_data = 64'h0;
  assign T_1824_client_id = T_1763_client_id;
  assign T_1861 = T_1519 | T_1657;
  assign GEN_0 = io_inner_release_bits_data;
  assign GEN_21 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_0;
  assign GEN_22 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_1;
  assign GEN_23 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_2;
  assign GEN_24 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_3;
  assign GEN_25 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_4;
  assign GEN_26 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_5;
  assign GEN_27 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_6;
  assign GEN_28 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_0 : data_buffer_7;
  assign GEN_30 = T_1520 ? GEN_21 : data_buffer_0;
  assign GEN_31 = T_1520 ? GEN_22 : data_buffer_1;
  assign GEN_32 = T_1520 ? GEN_23 : data_buffer_2;
  assign GEN_33 = T_1520 ? GEN_24 : data_buffer_3;
  assign GEN_34 = T_1520 ? GEN_25 : data_buffer_4;
  assign GEN_35 = T_1520 ? GEN_26 : data_buffer_5;
  assign GEN_36 = T_1520 ? GEN_27 : data_buffer_6;
  assign GEN_37 = T_1520 ? GEN_28 : data_buffer_7;
  assign T_1893_state = 2'h2;
  assign T_1922 = T_1552 | io_alloc_irel_should;
  assign T_1938 = T_1691 & T_1694;
  assign T_1939 = pending_orel_data | T_1938;
  assign T_1941 = io_outer_release_ready & io_outer_release_valid;
  assign T_1942 = io_outer_release_bits_r_type == 3'h0;
  assign T_1943 = io_outer_release_bits_r_type == 3'h1;
  assign T_1944 = io_outer_release_bits_r_type == 3'h2;
  assign T_1945 = T_1942 | T_1943;
  assign T_1946 = T_1945 | T_1944;
  assign T_1947 = T_1941 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1954 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_1955 = ~ T_1954;
  assign T_1956 = T_1952 | T_1955;
  assign T_1957 = T_1939 & T_1956;
  assign GEN_38 = T_1922 ? T_1957 : pending_orel_data;
  assign GEN_39 = T_1646 ? 1'h1 : pending_orel_send;
  assign T_1968 = T_1946 == 1'h0;
  assign T_1970 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_1971 = T_1968 | T_1970;
  assign GEN_40 = T_1971 ? 1'h1 : sending_orel;
  assign T_1983 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_1984 = T_1968 | T_1983;
  assign GEN_41 = T_1984 ? 1'h0 : GEN_40;
  assign GEN_42 = T_1941 ? GEN_41 : sending_orel;
  assign GEN_43 = T_1941 ? 1'h0 : GEN_39;
  assign T_1993 = T_1941 & io_outer_release_bits_voluntary;
  assign T_2001 = T_1993 & T_1946;
  assign T_2005 = T_2003 == 3'h7;
  assign T_2007 = T_2003 + 3'h1;
  assign T_2008 = T_2007[2:0];
  assign GEN_44 = T_2001 ? T_2008 : T_2003;
  assign T_2009 = T_2001 & T_2005;
  assign T_2010 = T_1946 ? T_2003 : 3'h0;
  assign T_2011 = T_1946 ? T_2009 : T_1993;
  assign T_2012 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2014 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2015 = io_outer_grant_bits_is_builtin_type & T_2014;
  assign T_2016 = T_2012 & T_2015;
  assign T_2024_0 = 3'h5;
  assign GEN_58 = {{1'd0}, T_2024_0};
  assign T_2026 = io_outer_grant_bits_g_type == GEN_58;
  assign T_2028 = io_outer_grant_bits_is_builtin_type ? T_2026 : T_2014;
  assign T_2030 = T_2016 & T_2028;
  assign T_2034 = T_2032 == 3'h7;
  assign T_2036 = T_2032 + 3'h1;
  assign T_2037 = T_2036[2:0];
  assign GEN_45 = T_2030 ? T_2037 : T_2032;
  assign T_2038 = T_2030 & T_2034;
  assign T_2039 = T_2028 ? T_2032 : 3'h0;
  assign T_2040 = T_2028 ? T_2038 : T_2016;
  assign T_2044 = T_2040 == 1'h0;
  assign T_2045 = T_2011 & T_2044;
  assign T_2047 = T_2042 + 1'h1;
  assign T_2048 = T_2047[0:0];
  assign GEN_46 = T_2045 ? T_2048 : T_2042;
  assign T_2050 = T_2011 == 1'h0;
  assign T_2051 = T_2040 & T_2050;
  assign T_2053 = T_2042 - 1'h1;
  assign T_2054 = T_2053[0:0];
  assign GEN_47 = T_2051 ? T_2054 : GEN_46;
  assign T_2056 = T_2042 > 1'h0;
  assign T_2065 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2066 = T_2065[0];
  assign T_2067 = T_1946 ? T_2066 : pending_orel_send;
  assign T_2068 = T_1721 & T_2067;
  assign T_2082 = T_1893_state == 2'h2;
  assign T_2083 = T_2082 ? 3'h0 : 3'h3;
  assign T_2119_addr_beat = vol_ognt_counter_up_idx;
  assign T_2119_addr_block = xact_addr_block;
  assign T_2119_client_xact_id = 3'h0;
  assign T_2119_voluntary = 1'h1;
  assign T_2119_r_type = T_2083;
  assign T_2119_data = GEN_1;
  assign GEN_1 = GEN_54;
  assign GEN_48 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_49 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_48;
  assign GEN_50 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_49;
  assign GEN_51 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_50;
  assign GEN_52 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_51;
  assign GEN_53 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_52;
  assign GEN_54 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_53;
  assign T_2149 = T_1656 | vol_ignt_counter_pending;
  assign T_2150 = T_2149 | scoreboard_2;
  assign T_2151 = T_2150 | vol_ognt_counter_pending;
  assign T_2153 = T_2151 == 1'h0;
  assign T_2155 = T_1721 & all_pending_done;
  assign GEN_56 = T_2155 ? 4'h0 : GEN_8;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_29 = GEN_92[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_55 = GEN_93[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_59 = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_60 = GEN_95[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_61 = GEN_96[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_62 = GEN_97[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_63 = GEN_98[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_64 = GEN_99[2:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_65 = GEN_100[10:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_66 = GEN_101[63:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_67 = GEN_102[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_68 = GEN_103[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_69 = {1{$random}};
  state = GEN_69[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_70 = {1{$random}};
  xact_addr_block = GEN_70[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_71 = {1{$random}};
  xact_vol_ir_r_type = GEN_71[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_72 = {1{$random}};
  xact_vol_ir_src = GEN_72[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_73 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_73[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_74 = {1{$random}};
  pending_irel_data = GEN_74[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_75 = {1{$random}};
  pending_orel_send = GEN_75[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_76 = {1{$random}};
  pending_orel_data = GEN_76[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_77 = {1{$random}};
  sending_orel = GEN_77[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {2{$random}};
  data_buffer_0 = GEN_78[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {2{$random}};
  data_buffer_1 = GEN_79[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {2{$random}};
  data_buffer_2 = GEN_80[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {2{$random}};
  data_buffer_3 = GEN_81[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {2{$random}};
  data_buffer_4 = GEN_82[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {2{$random}};
  data_buffer_5 = GEN_83[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {2{$random}};
  data_buffer_6 = GEN_84[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {2{$random}};
  data_buffer_7 = GEN_85[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  T_1588 = GEN_86[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  T_1619 = GEN_87[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  T_1629 = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {1{$random}};
  T_2003 = GEN_89[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  T_2032 = GEN_90[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {1{$random}};
  T_2042 = GEN_91[0:0];
  `endif
  GEN_92 = {1{$random}};
  GEN_93 = {1{$random}};
  GEN_94 = {1{$random}};
  GEN_95 = {1{$random}};
  GEN_96 = {1{$random}};
  GEN_97 = {1{$random}};
  GEN_98 = {1{$random}};
  GEN_99 = {1{$random}};
  GEN_100 = {1{$random}};
  GEN_101 = {2{$random}};
  GEN_102 = {1{$random}};
  GEN_103 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_2155) begin
        state <= 4'h0;
      end else begin
        if(T_1646) begin
          state <= 4'h7;
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_1646) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1661) begin
        if(T_1673) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_1661) begin
        if(T_1700) begin
          pending_irel_data <= T_1717;
        end else begin
          if(T_1673) begin
            if(T_1584) begin
              pending_irel_data <= T_1696;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_1646) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_1646) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_1941) begin
        pending_orel_send <= 1'h0;
      end else begin
        if(T_1646) begin
          pending_orel_send <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_1922) begin
        pending_orel_data <= T_1957;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_1941) begin
        if(T_1984) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_1971) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1544_0;
    end else begin
      if(T_1520) begin
        if(3'h0 == io_inner_release_bits_addr_beat) begin
          data_buffer_0 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1544_1;
    end else begin
      if(T_1520) begin
        if(3'h1 == io_inner_release_bits_addr_beat) begin
          data_buffer_1 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1544_2;
    end else begin
      if(T_1520) begin
        if(3'h2 == io_inner_release_bits_addr_beat) begin
          data_buffer_2 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1544_3;
    end else begin
      if(T_1520) begin
        if(3'h3 == io_inner_release_bits_addr_beat) begin
          data_buffer_3 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1544_4;
    end else begin
      if(T_1520) begin
        if(3'h4 == io_inner_release_bits_addr_beat) begin
          data_buffer_4 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1544_5;
    end else begin
      if(T_1520) begin
        if(3'h5 == io_inner_release_bits_addr_beat) begin
          data_buffer_5 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1544_6;
    end else begin
      if(T_1520) begin
        if(3'h6 == io_inner_release_bits_addr_beat) begin
          data_buffer_6 <= GEN_0;
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1544_7;
    end else begin
      if(T_1520) begin
        if(3'h7 == io_inner_release_bits_addr_beat) begin
          data_buffer_7 <= GEN_0;
        end
      end
    end
    if(reset) begin
      T_1588 <= 3'h0;
    end else begin
      if(T_1586) begin
        T_1588 <= T_1593;
      end
    end
    if(reset) begin
      T_1619 <= 3'h0;
    end else begin
      if(T_1617) begin
        T_1619 <= T_1624;
      end
    end
    if(reset) begin
      T_1629 <= 1'h0;
    end else begin
      if(T_1638) begin
        T_1629 <= T_1641;
      end else begin
        if(T_1632) begin
          T_1629 <= T_1635;
        end
      end
    end
    if(reset) begin
      T_2003 <= 3'h0;
    end else begin
      if(T_2001) begin
        T_2003 <= T_2008;
      end
    end
    if(reset) begin
      T_2032 <= 3'h0;
    end else begin
      if(T_2030) begin
        T_2032 <= T_2037;
      end
    end
    if(reset) begin
      T_2042 <= 1'h0;
    end else begin
      if(T_2051) begin
        T_2042 <= T_2054;
      end else begin
        if(T_2045) begin
          T_2042 <= T_2048;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1530) begin
          $fwrite(32'h80000002,"Assertion failed: VoluntaryReleaseTracker accepted Release that wasn't voluntary!\n    at Broadcast.scala:81 assert(!(state === s_idle && io.inner.release.fire() && io.alloc.irel.should && !io.irel().isVoluntary()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1530) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_10(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_client_id,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_client_id,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [1:0] io_count
);
  reg [1:0] ram_client_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_client_xact_id_T_294_data;
  wire  ram_client_xact_id_T_294_addr;
  wire  ram_client_xact_id_T_294_en;
  wire [1:0] ram_client_xact_id_T_253_data;
  wire  ram_client_xact_id_T_253_addr;
  wire  ram_client_xact_id_T_253_mask;
  wire  ram_client_xact_id_T_253_en;
  reg [2:0] ram_addr_beat [0:1];
  reg [31:0] GEN_1;
  wire [2:0] ram_addr_beat_T_294_data;
  wire  ram_addr_beat_T_294_addr;
  wire  ram_addr_beat_T_294_en;
  wire [2:0] ram_addr_beat_T_253_data;
  wire  ram_addr_beat_T_253_addr;
  wire  ram_addr_beat_T_253_mask;
  wire  ram_addr_beat_T_253_en;
  reg  ram_client_id [0:1];
  reg [31:0] GEN_2;
  wire  ram_client_id_T_294_data;
  wire  ram_client_id_T_294_addr;
  wire  ram_client_id_T_294_en;
  wire  ram_client_id_T_253_data;
  wire  ram_client_id_T_253_addr;
  wire  ram_client_id_T_253_mask;
  wire  ram_client_id_T_253_en;
  reg  ram_is_builtin_type [0:1];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_294_data;
  wire  ram_is_builtin_type_T_294_addr;
  wire  ram_is_builtin_type_T_294_en;
  wire  ram_is_builtin_type_T_253_data;
  wire  ram_is_builtin_type_T_253_addr;
  wire  ram_is_builtin_type_T_253_mask;
  wire  ram_is_builtin_type_T_253_en;
  reg [2:0] ram_a_type [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_294_data;
  wire  ram_a_type_T_294_addr;
  wire  ram_a_type_T_294_en;
  wire [2:0] ram_a_type_T_253_data;
  wire  ram_a_type_T_253_addr;
  wire  ram_a_type_T_253_mask;
  wire  ram_a_type_T_253_en;
  reg  T_245;
  reg [31:0] GEN_5;
  reg  T_247;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_250;
  wire  empty;
  wire  full;
  wire  T_251;
  wire  do_enq;
  wire  T_252;
  wire  do_deq;
  wire [1:0] T_282;
  wire  T_283;
  wire  GEN_13;
  wire [1:0] T_287;
  wire  T_288;
  wire  GEN_14;
  wire  T_289;
  wire  GEN_15;
  wire  T_291;
  wire  T_293;
  wire [1:0] T_320;
  wire  ptr_diff;
  wire  T_321;
  wire [1:0] T_322;
  assign io_enq_ready = T_293;
  assign io_deq_valid = T_291;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_294_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_294_data;
  assign io_deq_bits_client_id = ram_client_id_T_294_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_294_data;
  assign io_deq_bits_a_type = ram_a_type_T_294_data;
  assign io_count = T_322;
  assign ram_client_xact_id_T_294_addr = T_247;
  assign ram_client_xact_id_T_294_en = 1'h1;
  assign ram_client_xact_id_T_294_data = ram_client_xact_id[ram_client_xact_id_T_294_addr];
  assign ram_client_xact_id_T_253_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_253_addr = T_245;
  assign ram_client_xact_id_T_253_mask = do_enq;
  assign ram_client_xact_id_T_253_en = do_enq;
  assign ram_addr_beat_T_294_addr = T_247;
  assign ram_addr_beat_T_294_en = 1'h1;
  assign ram_addr_beat_T_294_data = ram_addr_beat[ram_addr_beat_T_294_addr];
  assign ram_addr_beat_T_253_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_253_addr = T_245;
  assign ram_addr_beat_T_253_mask = do_enq;
  assign ram_addr_beat_T_253_en = do_enq;
  assign ram_client_id_T_294_addr = T_247;
  assign ram_client_id_T_294_en = 1'h1;
  assign ram_client_id_T_294_data = ram_client_id[ram_client_id_T_294_addr];
  assign ram_client_id_T_253_data = io_enq_bits_client_id;
  assign ram_client_id_T_253_addr = T_245;
  assign ram_client_id_T_253_mask = do_enq;
  assign ram_client_id_T_253_en = do_enq;
  assign ram_is_builtin_type_T_294_addr = T_247;
  assign ram_is_builtin_type_T_294_en = 1'h1;
  assign ram_is_builtin_type_T_294_data = ram_is_builtin_type[ram_is_builtin_type_T_294_addr];
  assign ram_is_builtin_type_T_253_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_253_addr = T_245;
  assign ram_is_builtin_type_T_253_mask = do_enq;
  assign ram_is_builtin_type_T_253_en = do_enq;
  assign ram_a_type_T_294_addr = T_247;
  assign ram_a_type_T_294_en = 1'h1;
  assign ram_a_type_T_294_data = ram_a_type[ram_a_type_T_294_addr];
  assign ram_a_type_T_253_data = io_enq_bits_a_type;
  assign ram_a_type_T_253_addr = T_245;
  assign ram_a_type_T_253_mask = do_enq;
  assign ram_a_type_T_253_en = do_enq;
  assign ptr_match = T_245 == T_247;
  assign T_250 = maybe_full == 1'h0;
  assign empty = ptr_match & T_250;
  assign full = ptr_match & maybe_full;
  assign T_251 = io_enq_ready & io_enq_valid;
  assign do_enq = T_251;
  assign T_252 = io_deq_ready & io_deq_valid;
  assign do_deq = T_252;
  assign T_282 = T_245 + 1'h1;
  assign T_283 = T_282[0:0];
  assign GEN_13 = do_enq ? T_283 : T_245;
  assign T_287 = T_247 + 1'h1;
  assign T_288 = T_287[0:0];
  assign GEN_14 = do_deq ? T_288 : T_247;
  assign T_289 = do_enq != do_deq;
  assign GEN_15 = T_289 ? do_enq : maybe_full;
  assign T_291 = empty == 1'h0;
  assign T_293 = full == 1'h0;
  assign T_320 = T_245 - T_247;
  assign ptr_diff = T_320[0:0];
  assign T_321 = maybe_full & ptr_match;
  assign T_322 = {T_321,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_1[2:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_client_id[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_245 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_247 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_client_xact_id_T_253_en & ram_client_xact_id_T_253_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_253_addr] <= ram_client_xact_id_T_253_data;
    end
    if(ram_addr_beat_T_253_en & ram_addr_beat_T_253_mask) begin
      ram_addr_beat[ram_addr_beat_T_253_addr] <= ram_addr_beat_T_253_data;
    end
    if(ram_client_id_T_253_en & ram_client_id_T_253_mask) begin
      ram_client_id[ram_client_id_T_253_addr] <= ram_client_id_T_253_data;
    end
    if(ram_is_builtin_type_T_253_en & ram_is_builtin_type_T_253_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_253_addr] <= ram_is_builtin_type_T_253_data;
    end
    if(ram_a_type_T_253_en & ram_a_type_T_253_mask) begin
      ram_a_type[ram_a_type_T_253_addr] <= ram_a_type_T_253_data;
    end
    if(reset) begin
      T_245 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_245 <= T_283;
      end
    end
    if(reset) begin
      T_247 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_247 <= T_288;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module BufferedBroadcastAcquireTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire [1:0] xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg [1:0] xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire [1:0] ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire [1:0] ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire [1:0] T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire [1:0] GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire [1:0] GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire [1:0] T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire [1:0] T_2440_client_xact_id;
  wire [2:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [2:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [2:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [2:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [2:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire [1:0] T_3455_client_xact_id;
  wire [2:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire [1:0] GEN_341;
  wire [2:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_10 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 3'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 3'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 3'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 3'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 3'h1;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_1(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire [1:0] xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg [1:0] xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire [1:0] ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire [1:0] ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire [1:0] T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire [1:0] GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire [1:0] GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire [1:0] T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire [1:0] T_2440_client_xact_id;
  wire [2:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [2:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [2:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [2:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [2:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire [1:0] T_3455_client_xact_id;
  wire [2:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire [1:0] GEN_341;
  wire [2:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_10 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 3'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 3'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 3'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 3'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 3'h2;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_2(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire [1:0] xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg [1:0] xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire [1:0] ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire [1:0] ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire [1:0] T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire [1:0] GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire [1:0] GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire [1:0] T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire [1:0] T_2440_client_xact_id;
  wire [2:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [2:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [2:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [2:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [2:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire [1:0] T_3455_client_xact_id;
  wire [2:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire [1:0] GEN_341;
  wire [2:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_10 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 3'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 3'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 3'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 3'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 3'h3;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BufferedBroadcastAcquireTracker_3(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id,
  output  io_alloc_iacq_matches,
  output  io_alloc_iacq_can,
  input   io_alloc_iacq_should,
  output  io_alloc_irel_matches,
  output  io_alloc_irel_can,
  input   io_alloc_irel_should,
  output  io_alloc_oprb_matches,
  output  io_alloc_oprb_can,
  input   io_alloc_oprb_should,
  output  io_alloc_idle,
  output [25:0] io_alloc_addr_block
);
  wire  all_pending_done;
  reg [3:0] state;
  reg [31:0] GEN_32;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_33;
  reg  xact_allocate;
  reg [31:0] GEN_41;
  reg [4:0] xact_amo_shift_bytes;
  reg [31:0] GEN_42;
  reg [4:0] xact_op_code;
  reg [31:0] GEN_43;
  reg [2:0] xact_addr_byte;
  reg [31:0] GEN_47;
  reg [1:0] xact_op_size;
  reg [31:0] GEN_78;
  wire [2:0] xact_addr_beat;
  wire [1:0] xact_iacq_client_xact_id;
  wire [2:0] xact_iacq_addr_beat;
  wire  xact_iacq_client_id;
  wire  xact_iacq_is_builtin_type;
  wire [2:0] xact_iacq_a_type;
  reg [2:0] xact_vol_ir_r_type;
  reg [31:0] GEN_79;
  reg  xact_vol_ir_src;
  reg [31:0] GEN_80;
  reg [1:0] xact_vol_ir_client_xact_id;
  reg [31:0] GEN_81;
  reg [7:0] pending_irel_data;
  reg [31:0] GEN_82;
  wire  vol_ignt_counter_pending;
  wire [2:0] vol_ignt_counter_up_idx;
  wire  vol_ignt_counter_up_done;
  wire [2:0] vol_ignt_counter_down_idx;
  wire  vol_ignt_counter_down_done;
  wire  scoreboard_6;
  wire [2:0] ignt_data_idx;
  wire  ignt_data_done;
  wire  ifin_counter_pending;
  wire [2:0] ifin_counter_up_idx;
  wire  ifin_counter_up_done;
  wire [2:0] ifin_counter_down_idx;
  wire  ifin_counter_down_done;
  reg [7:0] pending_put_data;
  reg [31:0] GEN_83;
  reg [7:0] pending_ignt_data;
  reg [31:0] GEN_84;
  wire  ognt_counter_pending;
  wire [2:0] ognt_counter_up_idx;
  wire  ognt_counter_up_done;
  wire [2:0] ognt_counter_down_idx;
  wire  ognt_counter_down_done;
  reg  pending_iprbs;
  reg [31:0] GEN_85;
  reg  pending_orel_send;
  reg [31:0] GEN_86;
  reg [7:0] pending_orel_data;
  reg [31:0] GEN_87;
  wire  vol_ognt_counter_pending;
  wire [2:0] vol_ognt_counter_up_idx;
  wire  vol_ognt_counter_up_done;
  wire [2:0] vol_ognt_counter_down_idx;
  wire  vol_ognt_counter_down_done;
  wire  T_170;
  wire  T_171;
  wire  scoreboard_3;
  reg  sending_orel;
  reg [31:0] GEN_88;
  wire  T_195_sharers;
  wire [1:0] T_241_state;
  wire  coh_inner_sharers;
  wire [1:0] coh_outer_state;
  wire  T_1611;
  wire  T_1612;
  wire  T_1613;
  wire  T_1614;
  wire [2:0] T_1623_0;
  wire  T_1625;
  wire  T_1626;
  wire  T_1627;
  wire [2:0] T_1636_0;
  wire  T_1638;
  wire  T_1639;
  wire  T_1641;
  wire  T_1643;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire  T_1649;
  wire  T_1650;
  wire  T_1652;
  wire  T_1653;
  wire  T_1654;
  wire  T_1656;
  wire  T_1658;
  wire  T_1659;
  wire  T_1660;
  wire  T_1661;
  wire  T_1663;
  wire  T_1664;
  wire  T_1666;
  wire  T_1670;
  wire  T_1671;
  wire  T_1672;
  wire  T_1674;
  wire  T_1675;
  wire  T_1677;
  wire [63:0] T_1691_0;
  wire [63:0] T_1691_1;
  wire [63:0] T_1691_2;
  wire [63:0] T_1691_3;
  wire [63:0] T_1691_4;
  wire [63:0] T_1691_5;
  wire [63:0] T_1691_6;
  wire [63:0] T_1691_7;
  reg [63:0] data_buffer_0;
  reg [63:0] GEN_89;
  reg [63:0] data_buffer_1;
  reg [63:0] GEN_90;
  reg [63:0] data_buffer_2;
  reg [63:0] GEN_91;
  reg [63:0] data_buffer_3;
  reg [63:0] GEN_92;
  reg [63:0] data_buffer_4;
  reg [63:0] GEN_93;
  reg [63:0] data_buffer_5;
  reg [63:0] GEN_94;
  reg [63:0] data_buffer_6;
  reg [63:0] GEN_95;
  reg [63:0] data_buffer_7;
  reg [63:0] GEN_96;
  wire [7:0] T_1709_0;
  wire [7:0] T_1709_1;
  wire [7:0] T_1709_2;
  wire [7:0] T_1709_3;
  wire [7:0] T_1709_4;
  wire [7:0] T_1709_5;
  wire [7:0] T_1709_6;
  wire [7:0] T_1709_7;
  reg [7:0] wmask_buffer_0;
  reg [31:0] GEN_97;
  reg [7:0] wmask_buffer_1;
  reg [31:0] GEN_98;
  reg [7:0] wmask_buffer_2;
  reg [31:0] GEN_99;
  reg [7:0] wmask_buffer_3;
  reg [31:0] GEN_100;
  reg [7:0] wmask_buffer_4;
  reg [31:0] GEN_101;
  reg [7:0] wmask_buffer_5;
  reg [31:0] GEN_102;
  reg [7:0] wmask_buffer_6;
  reg [31:0] GEN_103;
  reg [7:0] wmask_buffer_7;
  reg [31:0] GEN_104;
  wire [7:0] T_1714;
  wire  T_1716;
  wire [7:0] T_1717;
  wire  T_1719;
  wire [7:0] T_1720;
  wire  T_1722;
  wire [7:0] T_1723;
  wire  T_1725;
  wire [7:0] T_1726;
  wire  T_1728;
  wire [7:0] T_1729;
  wire  T_1731;
  wire [7:0] T_1732;
  wire  T_1734;
  wire [7:0] T_1735;
  wire  T_1737;
  wire  data_valid_0;
  wire  data_valid_1;
  wire  data_valid_2;
  wire  data_valid_3;
  wire  data_valid_4;
  wire  data_valid_5;
  wire  data_valid_6;
  wire  data_valid_7;
  wire  T_1748;
  wire  T_1749;
  wire  T_1751;
  wire  T_1752;
  wire  T_1754;
  wire  T_1755;
  wire  T_1764;
  wire  T_1765;
  wire  T_1766;
  wire  T_1767;
  wire  T_1768;
  wire  T_1769;
  wire  ignt_q_clk;
  wire  ignt_q_reset;
  wire  ignt_q_io_enq_ready;
  wire  ignt_q_io_enq_valid;
  wire [1:0] ignt_q_io_enq_bits_client_xact_id;
  wire [2:0] ignt_q_io_enq_bits_addr_beat;
  wire  ignt_q_io_enq_bits_client_id;
  wire  ignt_q_io_enq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_enq_bits_a_type;
  wire  ignt_q_io_deq_ready;
  wire  ignt_q_io_deq_valid;
  wire [1:0] ignt_q_io_deq_bits_client_xact_id;
  wire [2:0] ignt_q_io_deq_bits_addr_beat;
  wire  ignt_q_io_deq_bits_client_id;
  wire  ignt_q_io_deq_bits_is_builtin_type;
  wire [2:0] ignt_q_io_deq_bits_a_type;
  wire [1:0] ignt_q_io_count;
  wire  T_1797;
  wire  T_1798;
  wire  T_1800;
  wire  T_1801;
  wire  T_1803;
  wire [2:0] T_1812_0;
  wire  T_1814;
  wire  T_1815;
  wire  T_1817;
  wire  T_1820;
  wire  T_1821;
  wire  T_1822;
  wire [1:0] T_1823_client_xact_id;
  wire [2:0] T_1823_addr_beat;
  wire  T_1823_client_id;
  wire  T_1823_is_builtin_type;
  wire [2:0] T_1823_a_type;
  wire  T_1850;
  wire  T_1852;
  wire [2:0] T_1862_0;
  wire [2:0] T_1862_1;
  wire [2:0] T_1862_2;
  wire  T_1864;
  wire  T_1865;
  wire  T_1866;
  wire  T_1867;
  wire  T_1868;
  wire  T_1869;
  wire  T_1870;
  wire [7:0] T_1874;
  wire [7:0] T_1875;
  wire [7:0] T_1877;
  wire [7:0] T_1878;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [2:0] T_1890_0;
  wire  T_1892;
  wire  T_1893;
  wire  T_1894;
  wire  T_1897;
  wire [7:0] T_1906;
  wire [7:0] T_1907;
  wire [7:0] GEN_34;
  wire [4:0] T_1915;
  wire  T_1917;
  wire  T_1918;
  wire  T_1920;
  wire  T_1921;
  wire  T_1922;
  wire [4:0] T_1923;
  wire [4:0] T_1924;
  wire [2:0] T_1925;
  wire [1:0] T_1926;
  wire [2:0] T_1939_0;
  wire [2:0] T_1939_1;
  wire [2:0] T_1939_2;
  wire  T_1941;
  wire  T_1942;
  wire  T_1943;
  wire  T_1944;
  wire  T_1945;
  wire  T_1946;
  wire  T_1947;
  wire [7:0] T_1951;
  wire [7:0] T_1952;
  wire [7:0] T_1956;
  wire [7:0] T_1958;
  wire [25:0] GEN_35;
  wire  GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [2:0] GEN_39;
  wire [1:0] GEN_40;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire [3:0] GEN_46;
  wire  scoreboard_0;
  wire [2:0] T_1976_0;
  wire  T_1978;
  wire  T_1979;
  wire  T_1980;
  wire  T_1981;
  wire [7:0] T_1982;
  wire  skip_outer_acquire;
  wire  T_1991;
  wire [1:0] T_1992;
  wire  T_1993;
  wire [1:0] T_1994;
  wire  T_1995;
  wire [1:0] T_1996;
  wire  T_1997;
  wire [1:0] T_1998;
  wire  T_1999;
  wire [1:0] T_2000;
  wire  T_2001;
  wire [1:0] T_2002;
  wire  T_2003;
  wire [1:0] T_2004;
  wire [1:0] T_2005;
  wire [25:0] T_2030_addr_block;
  wire [1:0] T_2030_p_type;
  wire  T_2030_client_id;
  wire  T_2055;
  wire [3:0] T_2056;
  wire  T_2065_pending;
  wire [2:0] T_2065_up_idx;
  wire  T_2065_up_done;
  wire [2:0] T_2065_down_idx;
  wire  T_2065_down_done;
  wire  T_2073;
  wire  T_2074;
  wire [1:0] T_2076;
  wire [1:0] T_2077;
  wire [1:0] GEN_410;
  wire [1:0] T_2078;
  wire [1:0] GEN_411;
  wire [1:0] T_2079;
  wire  T_2080;
  wire  T_2083;
  reg [2:0] T_2091;
  reg [31:0] GEN_105;
  wire  T_2100;
  wire  T_2103;
  wire  T_2104;
  wire  T_2105;
  wire  T_2107;
  wire  T_2108;
  wire  T_2109;
  wire  T_2110;
  wire  T_2111;
  wire  T_2113;
  reg [2:0] T_2115;
  reg [31:0] GEN_106;
  wire  T_2117;
  wire [3:0] T_2119;
  wire [2:0] T_2120;
  wire [2:0] GEN_48;
  wire  T_2121;
  wire [2:0] T_2122;
  wire  T_2123;
  reg  T_2125;
  reg [31:0] GEN_107;
  wire  T_2127;
  wire  T_2128;
  wire [1:0] T_2130;
  wire  T_2131;
  wire  GEN_49;
  wire  T_2133;
  wire  T_2134;
  wire [1:0] T_2136;
  wire  T_2137;
  wire  GEN_50;
  wire  T_2139;
  wire  T_2143;
  wire  T_2145;
  wire  T_2146;
  wire [3:0] GEN_51;
  wire  T_2150;
  wire  T_2151;
  wire  T_2156;
  wire  T_2164;
  reg [2:0] T_2166;
  reg [31:0] GEN_108;
  wire  T_2168;
  wire [3:0] T_2170;
  wire [2:0] T_2171;
  wire [2:0] GEN_52;
  wire  T_2172;
  wire [2:0] T_2173;
  wire  T_2174;
  wire  T_2175;
  wire  T_2178;
  wire  T_2179;
  wire  T_2180;
  wire  T_2181;
  wire [2:0] T_2189_0;
  wire [3:0] GEN_412;
  wire  T_2191;
  wire  T_2193;
  wire  T_2195;
  reg [2:0] T_2197;
  reg [31:0] GEN_109;
  wire  T_2199;
  wire [3:0] T_2201;
  wire [2:0] T_2202;
  wire [2:0] GEN_53;
  wire  T_2203;
  wire [2:0] T_2204;
  wire  T_2205;
  reg  T_2207;
  reg [31:0] GEN_110;
  wire  T_2209;
  wire  T_2210;
  wire [1:0] T_2212;
  wire  T_2213;
  wire  GEN_54;
  wire  T_2215;
  wire  T_2216;
  wire [1:0] T_2218;
  wire  T_2219;
  wire  GEN_55;
  wire  T_2221;
  wire  T_2223;
  wire  T_2224;
  wire [25:0] GEN_56;
  wire [7:0] GEN_57;
  wire [3:0] GEN_58;
  wire  T_2231;
  wire  T_2233;
  wire  T_2234;
  wire  T_2236;
  wire  T_2237;
  wire  T_2239;
  wire  T_2240;
  wire  T_2241;
  wire  T_2243;
  wire  T_2244;
  wire  T_2247;
  wire  T_2248;
  wire  T_2250;
  wire  T_2251;
  wire [7:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire  T_2263;
  wire  T_2264;
  wire  T_2266;
  wire  T_2267;
  wire  T_2271;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2286;
  wire  T_2288;
  wire  T_2289;
  wire [2:0] GEN_59;
  wire  GEN_60;
  wire [1:0] GEN_61;
  wire  T_2303;
  wire [7:0] T_2307;
  wire [7:0] T_2308;
  wire [7:0] T_2310;
  wire [7:0] T_2311;
  wire [7:0] T_2312;
  wire [7:0] T_2314;
  wire [2:0] GEN_62;
  wire  GEN_63;
  wire [1:0] GEN_64;
  wire [7:0] GEN_65;
  wire  T_2316;
  wire [7:0] T_2333;
  wire [7:0] GEN_66;
  wire [2:0] GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [7:0] GEN_70;
  wire  T_2334;
  wire  T_2335;
  wire  T_2337;
  wire  T_2338;
  wire  T_2339;
  wire  T_2340;
  wire  T_2341;
  wire  T_2343;
  wire  T_2344;
  wire  T_2346;
  wire  T_2347;
  wire [2:0] T_2379_addr_beat;
  wire [25:0] T_2379_addr_block;
  wire [1:0] T_2379_client_xact_id;
  wire  T_2379_voluntary;
  wire [2:0] T_2379_r_type;
  wire [63:0] T_2379_data;
  wire  T_2379_client_id;
  wire [2:0] T_2440_addr_beat;
  wire [1:0] T_2440_client_xact_id;
  wire [2:0] T_2440_manager_xact_id;
  wire  T_2440_is_builtin_type;
  wire [3:0] T_2440_g_type;
  wire [63:0] T_2440_data;
  wire  T_2440_client_id;
  wire [7:0] GEN_0;
  wire [7:0] GEN_71;
  wire [7:0] GEN_72;
  wire [7:0] GEN_73;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire  T_2521;
  wire [7:0] GEN_1;
  wire  T_2522;
  wire [7:0] GEN_2;
  wire  T_2523;
  wire [7:0] GEN_3;
  wire  T_2524;
  wire [7:0] GEN_4;
  wire  T_2525;
  wire [7:0] GEN_5;
  wire  T_2526;
  wire [7:0] GEN_6;
  wire  T_2527;
  wire [7:0] GEN_7;
  wire  T_2528;
  wire [7:0] T_2532;
  wire [7:0] T_2536;
  wire [7:0] T_2540;
  wire [7:0] T_2544;
  wire [7:0] T_2548;
  wire [7:0] T_2552;
  wire [7:0] T_2556;
  wire [7:0] T_2560;
  wire [15:0] T_2561;
  wire [15:0] T_2562;
  wire [31:0] T_2563;
  wire [15:0] T_2564;
  wire [15:0] T_2565;
  wire [31:0] T_2566;
  wire [63:0] T_2567;
  wire [63:0] T_2568;
  wire [63:0] T_2569;
  wire [63:0] GEN_8;
  wire [63:0] GEN_127;
  wire [63:0] GEN_128;
  wire [63:0] GEN_129;
  wire [63:0] GEN_130;
  wire [63:0] GEN_131;
  wire [63:0] GEN_132;
  wire [63:0] GEN_133;
  wire [63:0] T_2570;
  wire [63:0] T_2571;
  wire [63:0] GEN_9;
  wire [63:0] GEN_134;
  wire [63:0] GEN_135;
  wire [63:0] GEN_136;
  wire [63:0] GEN_137;
  wire [63:0] GEN_138;
  wire [63:0] GEN_139;
  wire [63:0] GEN_140;
  wire [63:0] GEN_141;
  wire [7:0] GEN_10;
  wire [7:0] GEN_142;
  wire [7:0] GEN_143;
  wire [7:0] GEN_144;
  wire [7:0] GEN_145;
  wire [7:0] GEN_146;
  wire [7:0] GEN_147;
  wire [7:0] GEN_148;
  wire [7:0] GEN_149;
  wire [63:0] GEN_160;
  wire [63:0] GEN_161;
  wire [63:0] GEN_162;
  wire [63:0] GEN_163;
  wire [63:0] GEN_164;
  wire [63:0] GEN_165;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [7:0] GEN_169;
  wire [7:0] GEN_170;
  wire [7:0] GEN_171;
  wire [7:0] GEN_172;
  wire [7:0] GEN_173;
  wire [7:0] GEN_174;
  wire [7:0] GEN_175;
  wire [7:0] GEN_176;
  wire [1:0] T_2604_state;
  wire  T_2631;
  wire [7:0] T_2647;
  wire [7:0] T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2656;
  wire [7:0] T_2660;
  wire [7:0] T_2661;
  wire [7:0] T_2663;
  wire [7:0] T_2664;
  wire [7:0] T_2665;
  wire [7:0] T_2666;
  wire [7:0] GEN_177;
  wire  T_2677;
  wire  T_2679;
  wire  T_2680;
  wire  GEN_179;
  wire  T_2692;
  wire  T_2693;
  wire  GEN_180;
  wire  GEN_181;
  wire  GEN_182;
  wire  T_2702;
  wire  T_2710;
  reg [2:0] T_2712;
  reg [31:0] GEN_111;
  wire  T_2714;
  wire [3:0] T_2716;
  wire [2:0] T_2717;
  wire [2:0] GEN_183;
  wire  T_2718;
  wire [2:0] T_2719;
  wire  T_2720;
  wire  T_2723;
  wire  T_2724;
  wire  T_2725;
  wire [2:0] T_2733_0;
  wire [3:0] GEN_413;
  wire  T_2735;
  wire  T_2737;
  wire  T_2739;
  reg [2:0] T_2741;
  reg [31:0] GEN_112;
  wire  T_2743;
  wire [3:0] T_2745;
  wire [2:0] T_2746;
  wire [2:0] GEN_184;
  wire  T_2747;
  wire [2:0] T_2748;
  wire  T_2749;
  reg  T_2751;
  reg [31:0] GEN_113;
  wire  T_2753;
  wire  T_2754;
  wire [1:0] T_2756;
  wire  T_2757;
  wire  GEN_185;
  wire  T_2759;
  wire  T_2760;
  wire [1:0] T_2762;
  wire  T_2763;
  wire  GEN_186;
  wire  T_2765;
  wire [7:0] T_2774;
  wire  T_2775;
  wire  T_2776;
  wire  T_2777;
  wire  T_2791;
  wire [2:0] T_2792;
  wire [2:0] T_2828_addr_beat;
  wire [25:0] T_2828_addr_block;
  wire [2:0] T_2828_client_xact_id;
  wire  T_2828_voluntary;
  wire [2:0] T_2828_r_type;
  wire [63:0] T_2828_data;
  wire [63:0] GEN_11;
  wire [63:0] GEN_187;
  wire [63:0] GEN_188;
  wire [63:0] GEN_189;
  wire [63:0] GEN_190;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [63:0] GEN_193;
  wire  T_2857;
  wire  T_2860;
  wire [2:0] T_2871_0;
  wire  T_2873;
  wire  T_2874;
  wire  T_2875;
  reg [2:0] T_2877;
  reg [31:0] GEN_114;
  wire  T_2879;
  wire [3:0] T_2881;
  wire [2:0] T_2882;
  wire [2:0] GEN_195;
  wire  T_2883;
  wire [2:0] T_2884;
  wire  T_2885;
  wire  T_2891;
  wire  T_2892;
  wire [2:0] T_2900_0;
  wire [3:0] GEN_414;
  wire  T_2902;
  wire  T_2904;
  wire  T_2906;
  reg [2:0] T_2908;
  reg [31:0] GEN_115;
  wire  T_2910;
  wire [3:0] T_2912;
  wire [2:0] T_2913;
  wire [2:0] GEN_196;
  wire  T_2914;
  wire [2:0] T_2915;
  wire  T_2916;
  reg  T_2918;
  reg [31:0] GEN_116;
  wire  T_2920;
  wire  T_2921;
  wire [1:0] T_2923;
  wire  T_2924;
  wire  GEN_197;
  wire  T_2926;
  wire  T_2927;
  wire [1:0] T_2929;
  wire  T_2930;
  wire  GEN_198;
  wire  T_2932;
  wire  T_2933;
  wire [7:0] T_2937;
  wire  T_2938;
  wire  T_2940;
  wire [2:0] T_2949_0;
  wire [2:0] T_2949_1;
  wire [2:0] T_2949_2;
  wire  T_2967;
  wire  T_2968;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire [5:0] T_2984;
  wire [25:0] T_3015_addr_block;
  wire [2:0] T_3015_client_xact_id;
  wire [2:0] T_3015_addr_beat;
  wire  T_3015_is_builtin_type;
  wire [2:0] T_3015_a_type;
  wire [10:0] T_3015_union;
  wire [63:0] T_3015_data;
  wire [7:0] GEN_12;
  wire [7:0] GEN_199;
  wire [7:0] GEN_200;
  wire [7:0] GEN_201;
  wire [7:0] GEN_202;
  wire [7:0] GEN_203;
  wire [7:0] GEN_204;
  wire [7:0] GEN_205;
  wire [5:0] T_3080;
  wire [4:0] T_3081;
  wire [10:0] T_3082;
  wire [6:0] T_3084;
  wire [7:0] T_3085;
  wire [8:0] T_3087;
  wire [5:0] T_3099;
  wire [5:0] T_3101;
  wire [10:0] T_3103;
  wire [10:0] T_3105;
  wire [10:0] T_3107;
  wire [10:0] T_3109;
  wire [10:0] T_3111;
  wire [25:0] T_3140_addr_block;
  wire [2:0] T_3140_client_xact_id;
  wire [2:0] T_3140_addr_beat;
  wire  T_3140_is_builtin_type;
  wire [2:0] T_3140_a_type;
  wire [10:0] T_3140_union;
  wire [63:0] T_3140_data;
  wire [63:0] GEN_13;
  wire [63:0] GEN_206;
  wire [63:0] GEN_207;
  wire [63:0] GEN_208;
  wire [63:0] GEN_209;
  wire [63:0] GEN_210;
  wire [63:0] GEN_211;
  wire [63:0] GEN_212;
  wire [25:0] T_3168_addr_block;
  wire [2:0] T_3168_client_xact_id;
  wire [2:0] T_3168_addr_beat;
  wire  T_3168_is_builtin_type;
  wire [2:0] T_3168_a_type;
  wire [10:0] T_3168_union;
  wire [63:0] T_3168_data;
  wire  T_3197;
  wire [3:0] GEN_213;
  wire  GEN_214;
  wire [2:0] T_3207_0;
  wire [2:0] T_3207_1;
  wire [3:0] GEN_415;
  wire  T_3209;
  wire [3:0] GEN_416;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3214;
  wire [7:0] GEN_14;
  wire [7:0] GEN_215;
  wire [7:0] GEN_216;
  wire [7:0] GEN_217;
  wire [7:0] GEN_218;
  wire [7:0] GEN_219;
  wire [7:0] GEN_220;
  wire [7:0] GEN_221;
  wire  T_3215;
  wire [7:0] GEN_15;
  wire  T_3216;
  wire [7:0] GEN_16;
  wire  T_3217;
  wire [7:0] GEN_17;
  wire  T_3218;
  wire [7:0] GEN_18;
  wire  T_3219;
  wire [7:0] GEN_19;
  wire  T_3220;
  wire [7:0] GEN_20;
  wire  T_3221;
  wire [7:0] GEN_21;
  wire  T_3222;
  wire [7:0] T_3226;
  wire [7:0] T_3230;
  wire [7:0] T_3234;
  wire [7:0] T_3238;
  wire [7:0] T_3242;
  wire [7:0] T_3246;
  wire [7:0] T_3250;
  wire [7:0] T_3254;
  wire [15:0] T_3255;
  wire [15:0] T_3256;
  wire [31:0] T_3257;
  wire [15:0] T_3258;
  wire [15:0] T_3259;
  wire [31:0] T_3260;
  wire [63:0] T_3261;
  wire [63:0] T_3262;
  wire [63:0] T_3263;
  wire [63:0] GEN_22;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [63:0] GEN_273;
  wire [63:0] GEN_274;
  wire [63:0] GEN_275;
  wire [63:0] GEN_276;
  wire [63:0] GEN_277;
  wire [63:0] T_3264;
  wire [63:0] T_3265;
  wire [63:0] GEN_23;
  wire [63:0] GEN_278;
  wire [63:0] GEN_279;
  wire [63:0] GEN_280;
  wire [63:0] GEN_281;
  wire [63:0] GEN_282;
  wire [63:0] GEN_283;
  wire [63:0] GEN_284;
  wire [63:0] GEN_285;
  wire [7:0] GEN_24;
  wire [7:0] GEN_286;
  wire [7:0] GEN_287;
  wire [7:0] GEN_288;
  wire [7:0] GEN_289;
  wire [7:0] GEN_290;
  wire [7:0] GEN_291;
  wire [7:0] GEN_292;
  wire [7:0] GEN_293;
  wire [63:0] GEN_304;
  wire [63:0] GEN_305;
  wire [63:0] GEN_306;
  wire [63:0] GEN_307;
  wire [63:0] GEN_308;
  wire [63:0] GEN_309;
  wire [63:0] GEN_310;
  wire [63:0] GEN_311;
  wire [7:0] GEN_313;
  wire [7:0] GEN_314;
  wire [7:0] GEN_315;
  wire [7:0] GEN_316;
  wire [7:0] GEN_317;
  wire [7:0] GEN_318;
  wire [7:0] GEN_319;
  wire [7:0] GEN_320;
  wire  T_3268;
  wire  T_3269;
  wire  T_3281;
  wire  T_3283;
  wire [2:0] T_3291_0;
  wire [3:0] GEN_417;
  wire  T_3293;
  wire  T_3295;
  wire  T_3297;
  reg [2:0] T_3299;
  reg [31:0] GEN_117;
  wire  T_3301;
  wire [3:0] T_3303;
  wire [2:0] T_3304;
  wire [2:0] GEN_321;
  wire  T_3305;
  wire [2:0] T_3306;
  wire  T_3307;
  wire  T_3308;
  reg [2:0] T_3314;
  reg [31:0] GEN_118;
  reg  T_3324;
  reg [31:0] GEN_119;
  wire  T_3326;
  wire  T_3327;
  wire [1:0] T_3329;
  wire  T_3330;
  wire  GEN_323;
  wire  T_3332;
  wire  T_3333;
  wire [1:0] T_3335;
  wire  T_3336;
  wire  GEN_324;
  wire  T_3338;
  wire  T_3343;
  wire [7:0] T_3360;
  wire [2:0] T_3370_0;
  wire [2:0] T_3370_1;
  wire [3:0] GEN_418;
  wire  T_3372;
  wire [3:0] GEN_419;
  wire  T_3373;
  wire  T_3374;
  wire  T_3376;
  wire  T_3377;
  wire [7:0] T_3382;
  wire [7:0] T_3384;
  wire [7:0] T_3385;
  wire [7:0] T_3386;
  wire [7:0] GEN_327;
  wire  T_3389;
  wire  T_3390;
  wire  T_3393;
  wire  T_3395;
  wire  T_3412;
  wire [2:0] T_3413;
  wire  T_3414;
  wire [2:0] T_3415;
  wire  T_3416;
  wire [2:0] T_3417;
  wire  T_3418;
  wire [2:0] T_3419;
  wire  T_3420;
  wire [2:0] T_3421;
  wire  T_3422;
  wire [2:0] T_3423;
  wire  T_3424;
  wire [2:0] T_3425;
  wire [2:0] T_3426;
  wire [2:0] T_3455_addr_beat;
  wire [1:0] T_3455_client_xact_id;
  wire [2:0] T_3455_manager_xact_id;
  wire  T_3455_is_builtin_type;
  wire [3:0] T_3455_g_type;
  wire [63:0] T_3455_data;
  wire  T_3455_client_id;
  wire [63:0] GEN_25;
  wire [63:0] GEN_328;
  wire [63:0] GEN_329;
  wire [63:0] GEN_330;
  wire [63:0] GEN_331;
  wire [63:0] GEN_332;
  wire [63:0] GEN_333;
  wire [63:0] GEN_334;
  wire [2:0] T_3491_0;
  wire [3:0] GEN_420;
  wire  T_3493;
  wire  T_3495;
  wire  T_3497;
  reg [2:0] T_3499;
  reg [31:0] GEN_120;
  wire  T_3501;
  wire [3:0] T_3503;
  wire [2:0] T_3504;
  wire [2:0] GEN_335;
  wire  T_3505;
  wire [2:0] T_3506;
  wire  T_3507;
  wire  T_3512;
  wire  T_3514;
  wire [2:0] T_3522_0;
  wire [2:0] T_3522_1;
  wire [3:0] GEN_421;
  wire  T_3524;
  wire [3:0] GEN_422;
  wire  T_3525;
  wire  T_3526;
  wire  T_3528;
  wire [7:0] T_3529;
  wire  T_3530;
  wire  T_3532;
  wire  T_3533;
  wire  GEN_338;
  wire  GEN_339;
  wire [2:0] GEN_340;
  wire [1:0] GEN_341;
  wire [2:0] GEN_342;
  wire  GEN_343;
  wire [3:0] GEN_344;
  wire [63:0] GEN_345;
  wire  GEN_346;
  wire  GEN_349;
  wire  T_3540;
  wire [1:0] GEN_350;
  wire  T_3551;
  wire  T_3552;
  wire [2:0] T_3562_0;
  wire [2:0] T_3562_1;
  wire [2:0] T_3562_2;
  wire  T_3564;
  wire  T_3565;
  wire  T_3566;
  wire  T_3567;
  wire  T_3568;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3573;
  wire  T_3574;
  wire  T_3603;
  wire [7:0] T_3604;
  wire [7:0] T_3606;
  wire [7:0] T_3607;
  wire  T_3608;
  wire  T_3609;
  wire  T_3610;
  wire  T_3611;
  wire  T_3612;
  wire  T_3613;
  wire  T_3614;
  wire  T_3615;
  wire [7:0] T_3619;
  wire [7:0] T_3623;
  wire [7:0] T_3627;
  wire [7:0] T_3631;
  wire [7:0] T_3635;
  wire [7:0] T_3639;
  wire [7:0] T_3643;
  wire [7:0] T_3647;
  wire [15:0] T_3648;
  wire [15:0] T_3649;
  wire [31:0] T_3650;
  wire [15:0] T_3651;
  wire [15:0] T_3652;
  wire [31:0] T_3653;
  wire [63:0] T_3654;
  wire [63:0] T_3655;
  wire [63:0] GEN_26;
  wire [63:0] GEN_351;
  wire [63:0] GEN_352;
  wire [63:0] GEN_353;
  wire [63:0] GEN_354;
  wire [63:0] GEN_355;
  wire [63:0] GEN_356;
  wire [63:0] GEN_357;
  wire [63:0] T_3656;
  wire [63:0] T_3657;
  wire [63:0] T_3658;
  wire [63:0] GEN_27;
  wire [63:0] GEN_358;
  wire [63:0] GEN_359;
  wire [63:0] GEN_360;
  wire [63:0] GEN_361;
  wire [63:0] GEN_362;
  wire [63:0] GEN_363;
  wire [63:0] GEN_364;
  wire [63:0] GEN_365;
  wire [7:0] GEN_28;
  wire [7:0] GEN_366;
  wire [7:0] GEN_367;
  wire [7:0] GEN_368;
  wire [7:0] GEN_369;
  wire [7:0] GEN_370;
  wire [7:0] GEN_371;
  wire [7:0] GEN_372;
  wire [7:0] T_3695;
  wire [7:0] GEN_29;
  wire [7:0] GEN_373;
  wire [7:0] GEN_374;
  wire [7:0] GEN_375;
  wire [7:0] GEN_376;
  wire [7:0] GEN_377;
  wire [7:0] GEN_378;
  wire [7:0] GEN_379;
  wire [7:0] GEN_380;
  wire [63:0] GEN_383;
  wire [63:0] GEN_384;
  wire [63:0] GEN_385;
  wire [63:0] GEN_386;
  wire [63:0] GEN_387;
  wire [63:0] GEN_388;
  wire [63:0] GEN_389;
  wire [63:0] GEN_390;
  wire [7:0] GEN_393;
  wire [7:0] GEN_394;
  wire [7:0] GEN_395;
  wire [7:0] GEN_396;
  wire [7:0] GEN_397;
  wire [7:0] GEN_398;
  wire [7:0] GEN_399;
  wire [7:0] GEN_400;
  wire  T_3698;
  wire  T_3699;
  wire  T_3700;
  wire  T_3701;
  wire  T_3702;
  wire  T_3703;
  wire  T_3704;
  wire  T_3706;
  wire  T_3708;
  wire [3:0] GEN_401;
  wire [7:0] GEN_402;
  wire [7:0] GEN_403;
  wire [7:0] GEN_404;
  wire [7:0] GEN_405;
  wire [7:0] GEN_406;
  wire [7:0] GEN_407;
  wire [7:0] GEN_408;
  wire [7:0] GEN_409;
  wire  GEN_30;
  reg [31:0] GEN_121;
  wire  GEN_31;
  reg [31:0] GEN_122;
  Queue_10 ignt_q (
    .clk(ignt_q_clk),
    .reset(ignt_q_reset),
    .io_enq_ready(ignt_q_io_enq_ready),
    .io_enq_valid(ignt_q_io_enq_valid),
    .io_enq_bits_client_xact_id(ignt_q_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(ignt_q_io_enq_bits_addr_beat),
    .io_enq_bits_client_id(ignt_q_io_enq_bits_client_id),
    .io_enq_bits_is_builtin_type(ignt_q_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(ignt_q_io_enq_bits_a_type),
    .io_deq_ready(ignt_q_io_deq_ready),
    .io_deq_valid(ignt_q_io_deq_valid),
    .io_deq_bits_client_xact_id(ignt_q_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(ignt_q_io_deq_bits_addr_beat),
    .io_deq_bits_client_id(ignt_q_io_deq_bits_client_id),
    .io_deq_bits_is_builtin_type(ignt_q_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(ignt_q_io_deq_bits_a_type),
    .io_count(ignt_q_io_count)
  );
  assign io_inner_acquire_ready = T_1981;
  assign io_inner_grant_valid = GEN_349;
  assign io_inner_grant_bits_addr_beat = GEN_340;
  assign io_inner_grant_bits_client_xact_id = GEN_341;
  assign io_inner_grant_bits_manager_xact_id = GEN_342;
  assign io_inner_grant_bits_is_builtin_type = GEN_343;
  assign io_inner_grant_bits_g_type = GEN_344;
  assign io_inner_grant_bits_data = GEN_345;
  assign io_inner_grant_bits_client_id = GEN_346;
  assign io_inner_finish_ready = T_2337;
  assign io_inner_probe_valid = T_2083;
  assign io_inner_probe_bits_addr_block = T_2030_addr_block;
  assign io_inner_probe_bits_p_type = T_2030_p_type;
  assign io_inner_probe_bits_client_id = T_2030_client_id;
  assign io_inner_release_ready = T_2274;
  assign io_outer_acquire_valid = T_2968;
  assign io_outer_acquire_bits_addr_block = T_3168_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_3168_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_3168_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_3168_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_3168_a_type;
  assign io_outer_acquire_bits_union = T_3168_union;
  assign io_outer_acquire_bits_data = T_3168_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = T_2777;
  assign io_outer_release_bits_addr_beat = T_2828_addr_beat;
  assign io_outer_release_bits_addr_block = T_2828_addr_block;
  assign io_outer_release_bits_client_xact_id = T_2828_client_xact_id;
  assign io_outer_release_bits_voluntary = T_2828_voluntary;
  assign io_outer_release_bits_r_type = T_2828_r_type;
  assign io_outer_release_bits_data = T_2828_data;
  assign io_outer_grant_ready = GEN_214;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_30;
  assign io_outer_finish_bits_manager_id = GEN_31;
  assign io_alloc_iacq_matches = T_1749;
  assign io_alloc_iacq_can = T_1611;
  assign io_alloc_irel_matches = T_1752;
  assign io_alloc_irel_can = 1'h0;
  assign io_alloc_oprb_matches = T_1755;
  assign io_alloc_oprb_can = 1'h0;
  assign io_alloc_idle = T_1611;
  assign io_alloc_addr_block = xact_addr_block;
  assign all_pending_done = T_3706;
  assign xact_addr_beat = xact_iacq_addr_beat;
  assign xact_iacq_client_xact_id = T_1823_client_xact_id;
  assign xact_iacq_addr_beat = T_1823_addr_beat;
  assign xact_iacq_client_id = T_1823_client_id;
  assign xact_iacq_is_builtin_type = T_1823_is_builtin_type;
  assign xact_iacq_a_type = T_1823_a_type;
  assign vol_ignt_counter_pending = T_2221;
  assign vol_ignt_counter_up_idx = T_2173;
  assign vol_ignt_counter_up_done = T_2174;
  assign vol_ignt_counter_down_idx = T_2204;
  assign vol_ignt_counter_down_done = T_2205;
  assign scoreboard_6 = T_1850;
  assign ignt_data_idx = T_3506;
  assign ignt_data_done = T_3507;
  assign ifin_counter_pending = T_3338;
  assign ifin_counter_up_idx = T_3306;
  assign ifin_counter_up_done = T_3307;
  assign ifin_counter_down_idx = 3'h0;
  assign ifin_counter_down_done = T_3308;
  assign ognt_counter_pending = T_2932;
  assign ognt_counter_up_idx = T_2884;
  assign ognt_counter_up_done = T_2885;
  assign ognt_counter_down_idx = T_2915;
  assign ognt_counter_down_done = T_2916;
  assign vol_ognt_counter_pending = T_2765;
  assign vol_ognt_counter_up_idx = T_2719;
  assign vol_ognt_counter_up_done = T_2720;
  assign vol_ognt_counter_down_idx = T_2748;
  assign vol_ognt_counter_down_done = T_2749;
  assign T_170 = pending_orel_data != 8'h0;
  assign T_171 = pending_orel_send | T_170;
  assign scoreboard_3 = T_171 | vol_ognt_counter_pending;
  assign T_195_sharers = 1'h0;
  assign T_241_state = 2'h0;
  assign coh_inner_sharers = T_195_sharers;
  assign coh_outer_state = T_241_state;
  assign T_1611 = state == 4'h0;
  assign T_1612 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_1613 = T_1611 & T_1612;
  assign T_1614 = T_1613 & io_alloc_iacq_should;
  assign T_1623_0 = 3'h3;
  assign T_1625 = io_inner_acquire_bits_a_type == T_1623_0;
  assign T_1626 = io_inner_acquire_bits_is_builtin_type & T_1625;
  assign T_1627 = T_1614 & T_1626;
  assign T_1636_0 = 3'h3;
  assign T_1638 = io_inner_acquire_bits_a_type == T_1636_0;
  assign T_1639 = io_inner_acquire_bits_is_builtin_type & T_1638;
  assign T_1641 = T_1639 == 1'h0;
  assign T_1643 = io_inner_acquire_bits_addr_beat == 3'h0;
  assign T_1644 = T_1641 | T_1643;
  assign T_1646 = T_1644 == 1'h0;
  assign T_1647 = T_1627 & T_1646;
  assign T_1649 = T_1647 == 1'h0;
  assign T_1650 = T_1649 | reset;
  assign T_1652 = T_1650 == 1'h0;
  assign T_1653 = state != 4'h0;
  assign T_1654 = T_1653 & scoreboard_6;
  assign T_1656 = xact_iacq_a_type == 3'h5;
  assign T_1658 = xact_iacq_a_type == 3'h6;
  assign T_1659 = T_1656 | T_1658;
  assign T_1660 = xact_iacq_is_builtin_type & T_1659;
  assign T_1661 = T_1654 & T_1660;
  assign T_1663 = T_1661 == 1'h0;
  assign T_1664 = T_1663 | reset;
  assign T_1666 = T_1664 == 1'h0;
  assign T_1670 = xact_iacq_a_type == 3'h4;
  assign T_1671 = xact_iacq_is_builtin_type & T_1670;
  assign T_1672 = T_1654 & T_1671;
  assign T_1674 = T_1672 == 1'h0;
  assign T_1675 = T_1674 | reset;
  assign T_1677 = T_1675 == 1'h0;
  assign T_1691_0 = 64'h0;
  assign T_1691_1 = 64'h0;
  assign T_1691_2 = 64'h0;
  assign T_1691_3 = 64'h0;
  assign T_1691_4 = 64'h0;
  assign T_1691_5 = 64'h0;
  assign T_1691_6 = 64'h0;
  assign T_1691_7 = 64'h0;
  assign T_1709_0 = 8'h0;
  assign T_1709_1 = 8'h0;
  assign T_1709_2 = 8'h0;
  assign T_1709_3 = 8'h0;
  assign T_1709_4 = 8'h0;
  assign T_1709_5 = 8'h0;
  assign T_1709_6 = 8'h0;
  assign T_1709_7 = 8'h0;
  assign T_1714 = ~ wmask_buffer_0;
  assign T_1716 = T_1714 == 8'h0;
  assign T_1717 = ~ wmask_buffer_1;
  assign T_1719 = T_1717 == 8'h0;
  assign T_1720 = ~ wmask_buffer_2;
  assign T_1722 = T_1720 == 8'h0;
  assign T_1723 = ~ wmask_buffer_3;
  assign T_1725 = T_1723 == 8'h0;
  assign T_1726 = ~ wmask_buffer_4;
  assign T_1728 = T_1726 == 8'h0;
  assign T_1729 = ~ wmask_buffer_5;
  assign T_1731 = T_1729 == 8'h0;
  assign T_1732 = ~ wmask_buffer_6;
  assign T_1734 = T_1732 == 8'h0;
  assign T_1735 = ~ wmask_buffer_7;
  assign T_1737 = T_1735 == 8'h0;
  assign data_valid_0 = T_1716;
  assign data_valid_1 = T_1719;
  assign data_valid_2 = T_1722;
  assign data_valid_3 = T_1725;
  assign data_valid_4 = T_1728;
  assign data_valid_5 = T_1731;
  assign data_valid_6 = T_1734;
  assign data_valid_7 = T_1737;
  assign T_1748 = io_inner_acquire_bits_addr_block == xact_addr_block;
  assign T_1749 = T_1653 & T_1748;
  assign T_1751 = io_inner_release_bits_addr_block == xact_addr_block;
  assign T_1752 = T_1653 & T_1751;
  assign T_1754 = io_outer_probe_bits_addr_block == xact_addr_block;
  assign T_1755 = T_1653 & T_1754;
  assign T_1764 = xact_iacq_client_xact_id == io_inner_acquire_bits_client_xact_id;
  assign T_1765 = xact_iacq_client_id == io_inner_acquire_bits_client_id;
  assign T_1766 = T_1764 & T_1765;
  assign T_1767 = T_1766 & scoreboard_6;
  assign T_1768 = xact_iacq_addr_beat == io_inner_acquire_bits_addr_beat;
  assign T_1769 = T_1767 & T_1768;
  assign ignt_q_clk = clk;
  assign ignt_q_reset = reset;
  assign ignt_q_io_enq_valid = T_1822;
  assign ignt_q_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign ignt_q_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign ignt_q_io_enq_bits_client_id = io_inner_acquire_bits_client_id;
  assign ignt_q_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign ignt_q_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign ignt_q_io_deq_ready = GEN_339;
  assign T_1797 = T_1611 & io_alloc_iacq_should;
  assign T_1798 = T_1797 & io_inner_acquire_valid;
  assign T_1800 = T_1769 == 1'h0;
  assign T_1801 = T_1800 & scoreboard_6;
  assign T_1803 = T_1801 & T_1612;
  assign T_1812_0 = 3'h3;
  assign T_1814 = io_inner_acquire_bits_a_type == T_1812_0;
  assign T_1815 = io_inner_acquire_bits_is_builtin_type & T_1814;
  assign T_1817 = T_1815 == 1'h0;
  assign T_1820 = T_1817 | T_1643;
  assign T_1821 = T_1803 & T_1820;
  assign T_1822 = T_1798 | T_1821;
  assign T_1823_client_xact_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_xact_id : ignt_q_io_enq_bits_client_xact_id;
  assign T_1823_addr_beat = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_addr_beat : ignt_q_io_enq_bits_addr_beat;
  assign T_1823_client_id = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_client_id : ignt_q_io_enq_bits_client_id;
  assign T_1823_is_builtin_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_is_builtin_type : ignt_q_io_enq_bits_is_builtin_type;
  assign T_1823_a_type = ignt_q_io_deq_valid ? ignt_q_io_deq_bits_a_type : ignt_q_io_enq_bits_a_type;
  assign T_1850 = ignt_q_io_count > 2'h0;
  assign T_1852 = T_1653 | io_alloc_iacq_should;
  assign T_1862_0 = 3'h2;
  assign T_1862_1 = 3'h3;
  assign T_1862_2 = 3'h4;
  assign T_1864 = io_inner_acquire_bits_a_type == T_1862_0;
  assign T_1865 = io_inner_acquire_bits_a_type == T_1862_1;
  assign T_1866 = io_inner_acquire_bits_a_type == T_1862_2;
  assign T_1867 = T_1864 | T_1865;
  assign T_1868 = T_1867 | T_1866;
  assign T_1869 = io_inner_acquire_bits_is_builtin_type & T_1868;
  assign T_1870 = T_1612 & T_1869;
  assign T_1874 = T_1870 ? 8'hff : 8'h0;
  assign T_1875 = ~ T_1874;
  assign T_1877 = 8'h1 << io_inner_acquire_bits_addr_beat;
  assign T_1878 = ~ T_1877;
  assign T_1879 = T_1875 | T_1878;
  assign T_1880 = pending_put_data & T_1879;
  assign T_1890_0 = 3'h3;
  assign T_1892 = io_inner_acquire_bits_a_type == T_1890_0;
  assign T_1893 = io_inner_acquire_bits_is_builtin_type & T_1892;
  assign T_1894 = T_1612 & T_1893;
  assign T_1897 = T_1894 & T_1643;
  assign T_1906 = T_1897 ? 8'hfe : 8'h0;
  assign T_1907 = T_1880 | T_1906;
  assign GEN_34 = T_1852 ? T_1907 : pending_put_data;
  assign T_1915 = 4'h8 * 4'h0;
  assign T_1917 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1918 = io_inner_acquire_bits_is_builtin_type & T_1917;
  assign T_1920 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1921 = io_inner_acquire_bits_is_builtin_type & T_1920;
  assign T_1922 = T_1918 | T_1921;
  assign T_1923 = io_inner_acquire_bits_union[5:1];
  assign T_1924 = T_1922 ? 5'h1 : T_1923;
  assign T_1925 = io_inner_acquire_bits_union[10:8];
  assign T_1926 = io_inner_acquire_bits_union[7:6];
  assign T_1939_0 = 3'h2;
  assign T_1939_1 = 3'h3;
  assign T_1939_2 = 3'h4;
  assign T_1941 = io_inner_acquire_bits_a_type == T_1939_0;
  assign T_1942 = io_inner_acquire_bits_a_type == T_1939_1;
  assign T_1943 = io_inner_acquire_bits_a_type == T_1939_2;
  assign T_1944 = T_1941 | T_1942;
  assign T_1945 = T_1944 | T_1943;
  assign T_1946 = io_inner_acquire_bits_is_builtin_type & T_1945;
  assign T_1947 = T_1612 & T_1946;
  assign T_1951 = T_1947 ? 8'hff : 8'h0;
  assign T_1952 = ~ T_1951;
  assign T_1956 = T_1952 | T_1878;
  assign T_1958 = T_1921 ? T_1956 : 8'h0;
  assign GEN_35 = T_1798 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_36 = T_1798 ? 1'h0 : xact_allocate;
  assign GEN_37 = T_1798 ? T_1915 : xact_amo_shift_bytes;
  assign GEN_38 = T_1798 ? T_1924 : xact_op_code;
  assign GEN_39 = T_1798 ? T_1925 : xact_addr_byte;
  assign GEN_40 = T_1798 ? T_1926 : xact_op_size;
  assign GEN_44 = T_1798 ? T_1958 : GEN_34;
  assign GEN_45 = T_1798 ? 8'h0 : pending_ignt_data;
  assign GEN_46 = T_1798 ? 4'h5 : state;
  assign scoreboard_0 = pending_put_data != 8'h0;
  assign T_1976_0 = 3'h3;
  assign T_1978 = io_inner_acquire_bits_a_type == T_1976_0;
  assign T_1979 = io_inner_acquire_bits_is_builtin_type & T_1978;
  assign T_1980 = T_1767 & T_1979;
  assign T_1981 = T_1611 | T_1980;
  assign T_1982 = ~ pending_ignt_data;
  assign skip_outer_acquire = T_1982 == 8'h0;
  assign T_1991 = 3'h4 == xact_iacq_a_type;
  assign T_1992 = T_1991 ? 2'h0 : 2'h2;
  assign T_1993 = 3'h6 == xact_iacq_a_type;
  assign T_1994 = T_1993 ? 2'h0 : T_1992;
  assign T_1995 = 3'h5 == xact_iacq_a_type;
  assign T_1996 = T_1995 ? 2'h2 : T_1994;
  assign T_1997 = 3'h2 == xact_iacq_a_type;
  assign T_1998 = T_1997 ? 2'h0 : T_1996;
  assign T_1999 = 3'h0 == xact_iacq_a_type;
  assign T_2000 = T_1999 ? 2'h2 : T_1998;
  assign T_2001 = 3'h3 == xact_iacq_a_type;
  assign T_2002 = T_2001 ? 2'h0 : T_2000;
  assign T_2003 = 3'h1 == xact_iacq_a_type;
  assign T_2004 = T_2003 ? 2'h2 : T_2002;
  assign T_2005 = xact_iacq_is_builtin_type ? T_2004 : 2'h0;
  assign T_2030_addr_block = xact_addr_block;
  assign T_2030_p_type = T_2005;
  assign T_2030_client_id = 1'h0;
  assign T_2055 = skip_outer_acquire == 1'h0;
  assign T_2056 = T_2055 ? 4'h6 : 4'h7;
  assign T_2065_pending = T_2139;
  assign T_2065_up_idx = 3'h0;
  assign T_2065_up_done = T_2073;
  assign T_2065_down_idx = T_2122;
  assign T_2065_down_done = T_2123;
  assign T_2073 = io_inner_probe_ready & io_inner_probe_valid;
  assign T_2074 = ~ T_2073;
  assign T_2076 = 2'h1 << io_inner_probe_bits_client_id;
  assign T_2077 = ~ T_2076;
  assign GEN_410 = {{1'd0}, T_2074};
  assign T_2078 = GEN_410 | T_2077;
  assign GEN_411 = {{1'd0}, pending_iprbs};
  assign T_2079 = GEN_411 & T_2078;
  assign T_2080 = state == 4'h5;
  assign T_2083 = T_2080 & pending_iprbs;
  assign T_2100 = io_inner_release_ready & io_inner_release_valid;
  assign T_2103 = io_inner_release_bits_voluntary == 1'h0;
  assign T_2104 = T_1653 & T_2103;
  assign T_2105 = T_2100 & T_2104;
  assign T_2107 = io_inner_release_bits_r_type == 3'h0;
  assign T_2108 = io_inner_release_bits_r_type == 3'h1;
  assign T_2109 = io_inner_release_bits_r_type == 3'h2;
  assign T_2110 = T_2107 | T_2108;
  assign T_2111 = T_2110 | T_2109;
  assign T_2113 = T_2105 & T_2111;
  assign T_2117 = T_2115 == 3'h7;
  assign T_2119 = T_2115 + 3'h1;
  assign T_2120 = T_2119[2:0];
  assign GEN_48 = T_2113 ? T_2120 : T_2115;
  assign T_2121 = T_2113 & T_2117;
  assign T_2122 = T_2111 ? T_2115 : 3'h0;
  assign T_2123 = T_2111 ? T_2121 : T_2105;
  assign T_2127 = T_2123 == 1'h0;
  assign T_2128 = T_2073 & T_2127;
  assign T_2130 = T_2125 + 1'h1;
  assign T_2131 = T_2130[0:0];
  assign GEN_49 = T_2128 ? T_2131 : T_2125;
  assign T_2133 = T_2073 == 1'h0;
  assign T_2134 = T_2123 & T_2133;
  assign T_2136 = T_2125 - 1'h1;
  assign T_2137 = T_2136[0:0];
  assign GEN_50 = T_2134 ? T_2137 : GEN_49;
  assign T_2139 = T_2125 > 1'h0;
  assign T_2143 = pending_iprbs | T_2065_pending;
  assign T_2145 = T_2143 == 1'h0;
  assign T_2146 = T_2080 & T_2145;
  assign GEN_51 = T_2146 ? T_2056 : GEN_46;
  assign T_2150 = T_1611 ? io_alloc_irel_should : io_alloc_irel_matches;
  assign T_2151 = T_2150 & io_inner_release_bits_voluntary;
  assign T_2156 = T_2100 & T_2151;
  assign T_2164 = T_2156 & T_2111;
  assign T_2168 = T_2166 == 3'h7;
  assign T_2170 = T_2166 + 3'h1;
  assign T_2171 = T_2170[2:0];
  assign GEN_52 = T_2164 ? T_2171 : T_2166;
  assign T_2172 = T_2164 & T_2168;
  assign T_2173 = T_2111 ? T_2166 : 3'h0;
  assign T_2174 = T_2111 ? T_2172 : T_2156;
  assign T_2175 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_2178 = io_inner_grant_bits_g_type == 4'h0;
  assign T_2179 = io_inner_grant_bits_is_builtin_type & T_2178;
  assign T_2180 = T_1653 & T_2179;
  assign T_2181 = T_2175 & T_2180;
  assign T_2189_0 = 3'h5;
  assign GEN_412 = {{1'd0}, T_2189_0};
  assign T_2191 = io_inner_grant_bits_g_type == GEN_412;
  assign T_2193 = io_inner_grant_bits_is_builtin_type ? T_2191 : T_2178;
  assign T_2195 = T_2181 & T_2193;
  assign T_2199 = T_2197 == 3'h7;
  assign T_2201 = T_2197 + 3'h1;
  assign T_2202 = T_2201[2:0];
  assign GEN_53 = T_2195 ? T_2202 : T_2197;
  assign T_2203 = T_2195 & T_2199;
  assign T_2204 = T_2193 ? T_2197 : 3'h0;
  assign T_2205 = T_2193 ? T_2203 : T_2181;
  assign T_2209 = T_2205 == 1'h0;
  assign T_2210 = T_2174 & T_2209;
  assign T_2212 = T_2207 + 1'h1;
  assign T_2213 = T_2212[0:0];
  assign GEN_54 = T_2210 ? T_2213 : T_2207;
  assign T_2215 = T_2174 == 1'h0;
  assign T_2216 = T_2205 & T_2215;
  assign T_2218 = T_2207 - 1'h1;
  assign T_2219 = T_2218[0:0];
  assign GEN_55 = T_2216 ? T_2219 : GEN_54;
  assign T_2221 = T_2207 > 1'h0;
  assign T_2223 = T_1611 & io_alloc_irel_should;
  assign T_2224 = T_2223 & io_inner_release_valid;
  assign GEN_56 = T_2224 ? io_inner_release_bits_addr_block : GEN_35;
  assign GEN_57 = T_2224 ? 8'hff : pending_irel_data;
  assign GEN_58 = T_2224 ? 4'h7 : GEN_51;
  assign T_2231 = T_1751 & io_inner_release_bits_voluntary;
  assign T_2233 = state == 4'h8;
  assign T_2234 = T_1611 | T_2233;
  assign T_2236 = T_2234 == 1'h0;
  assign T_2237 = T_2231 & T_2236;
  assign T_2239 = all_pending_done == 1'h0;
  assign T_2240 = T_2237 & T_2239;
  assign T_2241 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_2243 = T_2241 == 1'h0;
  assign T_2244 = T_2240 & T_2243;
  assign T_2247 = T_2175 == 1'h0;
  assign T_2248 = T_2244 & T_2247;
  assign T_2250 = vol_ignt_counter_pending == 1'h0;
  assign T_2251 = T_2248 & T_2250;
  assign T_2252 = pending_orel_data >> io_inner_release_bits_addr_beat;
  assign T_2253 = T_2252[0];
  assign T_2254 = sending_orel & T_2253;
  assign T_2255 = io_outer_release_ready & io_outer_release_valid;
  assign T_2256 = io_inner_release_bits_addr_beat == io_outer_release_bits_addr_beat;
  assign T_2257 = T_2255 & T_2256;
  assign T_2263 = T_2254 | T_2257;
  assign T_2264 = T_2111 & T_2263;
  assign T_2266 = T_2264 == 1'h0;
  assign T_2267 = T_2251 & T_2266;
  assign T_2271 = T_1751 & T_2103;
  assign T_2273 = T_2271 & T_2080;
  assign T_2274 = T_2267 | T_2273;
  assign T_2275 = T_2274 & io_inner_release_valid;
  assign T_2276 = T_2224 | T_2275;
  assign T_2277 = T_2276 & io_inner_release_ready;
  assign T_2286 = T_2111 == 1'h0;
  assign T_2288 = io_inner_release_bits_addr_beat == 3'h0;
  assign T_2289 = T_2286 | T_2288;
  assign GEN_59 = io_inner_release_bits_voluntary ? io_inner_release_bits_r_type : xact_vol_ir_r_type;
  assign GEN_60 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_id : xact_vol_ir_src;
  assign GEN_61 = io_inner_release_bits_voluntary ? io_inner_release_bits_client_xact_id : xact_vol_ir_client_xact_id;
  assign T_2303 = T_2100 & T_2111;
  assign T_2307 = T_2303 ? 8'hff : 8'h0;
  assign T_2308 = ~ T_2307;
  assign T_2310 = 8'h1 << io_inner_release_bits_addr_beat;
  assign T_2311 = ~ T_2310;
  assign T_2312 = T_2308 | T_2311;
  assign T_2314 = T_2111 ? T_2312 : 8'h0;
  assign GEN_62 = T_2289 ? GEN_59 : xact_vol_ir_r_type;
  assign GEN_63 = T_2289 ? GEN_60 : xact_vol_ir_src;
  assign GEN_64 = T_2289 ? GEN_61 : xact_vol_ir_client_xact_id;
  assign GEN_65 = T_2289 ? T_2314 : GEN_57;
  assign T_2316 = T_2289 == 1'h0;
  assign T_2333 = pending_irel_data & T_2312;
  assign GEN_66 = T_2316 ? T_2333 : GEN_65;
  assign GEN_67 = T_2277 ? GEN_62 : xact_vol_ir_r_type;
  assign GEN_68 = T_2277 ? GEN_63 : xact_vol_ir_src;
  assign GEN_69 = T_2277 ? GEN_64 : xact_vol_ir_client_xact_id;
  assign GEN_70 = T_2277 ? GEN_66 : GEN_57;
  assign T_2334 = state == 4'h3;
  assign T_2335 = state == 4'h4;
  assign T_2337 = state == 4'h7;
  assign T_2338 = T_2334 | T_2335;
  assign T_2339 = T_2338 | T_2080;
  assign T_2340 = T_2339 | T_2337;
  assign T_2341 = T_2340 & vol_ignt_counter_pending;
  assign T_2343 = pending_irel_data != 8'h0;
  assign T_2344 = T_2343 | vol_ognt_counter_pending;
  assign T_2346 = T_2344 == 1'h0;
  assign T_2347 = T_2341 & T_2346;
  assign T_2379_addr_beat = 3'h0;
  assign T_2379_addr_block = xact_addr_block;
  assign T_2379_client_xact_id = xact_vol_ir_client_xact_id;
  assign T_2379_voluntary = 1'h1;
  assign T_2379_r_type = xact_vol_ir_r_type;
  assign T_2379_data = 64'h0;
  assign T_2379_client_id = xact_vol_ir_src;
  assign T_2440_addr_beat = 3'h0;
  assign T_2440_client_xact_id = T_2379_client_xact_id;
  assign T_2440_manager_xact_id = 3'h0;
  assign T_2440_is_builtin_type = 1'h1;
  assign T_2440_g_type = 4'h0;
  assign T_2440_data = 64'h0;
  assign T_2440_client_id = T_2379_client_id;
  assign GEN_0 = GEN_77;
  assign GEN_71 = 3'h1 == io_inner_release_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_72 = 3'h2 == io_inner_release_bits_addr_beat ? wmask_buffer_2 : GEN_71;
  assign GEN_73 = 3'h3 == io_inner_release_bits_addr_beat ? wmask_buffer_3 : GEN_72;
  assign GEN_74 = 3'h4 == io_inner_release_bits_addr_beat ? wmask_buffer_4 : GEN_73;
  assign GEN_75 = 3'h5 == io_inner_release_bits_addr_beat ? wmask_buffer_5 : GEN_74;
  assign GEN_76 = 3'h6 == io_inner_release_bits_addr_beat ? wmask_buffer_6 : GEN_75;
  assign GEN_77 = 3'h7 == io_inner_release_bits_addr_beat ? wmask_buffer_7 : GEN_76;
  assign T_2521 = GEN_0[0];
  assign GEN_1 = GEN_77;
  assign T_2522 = GEN_1[1];
  assign GEN_2 = GEN_77;
  assign T_2523 = GEN_2[2];
  assign GEN_3 = GEN_77;
  assign T_2524 = GEN_3[3];
  assign GEN_4 = GEN_77;
  assign T_2525 = GEN_4[4];
  assign GEN_5 = GEN_77;
  assign T_2526 = GEN_5[5];
  assign GEN_6 = GEN_77;
  assign T_2527 = GEN_6[6];
  assign GEN_7 = GEN_77;
  assign T_2528 = GEN_7[7];
  assign T_2532 = T_2521 ? 8'hff : 8'h0;
  assign T_2536 = T_2522 ? 8'hff : 8'h0;
  assign T_2540 = T_2523 ? 8'hff : 8'h0;
  assign T_2544 = T_2524 ? 8'hff : 8'h0;
  assign T_2548 = T_2525 ? 8'hff : 8'h0;
  assign T_2552 = T_2526 ? 8'hff : 8'h0;
  assign T_2556 = T_2527 ? 8'hff : 8'h0;
  assign T_2560 = T_2528 ? 8'hff : 8'h0;
  assign T_2561 = {T_2536,T_2532};
  assign T_2562 = {T_2544,T_2540};
  assign T_2563 = {T_2562,T_2561};
  assign T_2564 = {T_2552,T_2548};
  assign T_2565 = {T_2560,T_2556};
  assign T_2566 = {T_2565,T_2564};
  assign T_2567 = {T_2566,T_2563};
  assign T_2568 = ~ T_2567;
  assign T_2569 = T_2568 & io_inner_release_bits_data;
  assign GEN_8 = GEN_133;
  assign GEN_127 = 3'h1 == io_inner_release_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_128 = 3'h2 == io_inner_release_bits_addr_beat ? data_buffer_2 : GEN_127;
  assign GEN_129 = 3'h3 == io_inner_release_bits_addr_beat ? data_buffer_3 : GEN_128;
  assign GEN_130 = 3'h4 == io_inner_release_bits_addr_beat ? data_buffer_4 : GEN_129;
  assign GEN_131 = 3'h5 == io_inner_release_bits_addr_beat ? data_buffer_5 : GEN_130;
  assign GEN_132 = 3'h6 == io_inner_release_bits_addr_beat ? data_buffer_6 : GEN_131;
  assign GEN_133 = 3'h7 == io_inner_release_bits_addr_beat ? data_buffer_7 : GEN_132;
  assign T_2570 = T_2567 & GEN_8;
  assign T_2571 = T_2569 | T_2570;
  assign GEN_9 = T_2571;
  assign GEN_134 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_0;
  assign GEN_135 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_1;
  assign GEN_136 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_2;
  assign GEN_137 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_3;
  assign GEN_138 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_4;
  assign GEN_139 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_5;
  assign GEN_140 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_6;
  assign GEN_141 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_9 : data_buffer_7;
  assign GEN_10 = 8'hff;
  assign GEN_142 = 3'h0 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_0;
  assign GEN_143 = 3'h1 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_1;
  assign GEN_144 = 3'h2 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_2;
  assign GEN_145 = 3'h3 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_3;
  assign GEN_146 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_4;
  assign GEN_147 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_5;
  assign GEN_148 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_6;
  assign GEN_149 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_10 : wmask_buffer_7;
  assign GEN_160 = T_2303 ? GEN_134 : data_buffer_0;
  assign GEN_161 = T_2303 ? GEN_135 : data_buffer_1;
  assign GEN_162 = T_2303 ? GEN_136 : data_buffer_2;
  assign GEN_163 = T_2303 ? GEN_137 : data_buffer_3;
  assign GEN_164 = T_2303 ? GEN_138 : data_buffer_4;
  assign GEN_165 = T_2303 ? GEN_139 : data_buffer_5;
  assign GEN_166 = T_2303 ? GEN_140 : data_buffer_6;
  assign GEN_167 = T_2303 ? GEN_141 : data_buffer_7;
  assign GEN_169 = T_2303 ? GEN_142 : wmask_buffer_0;
  assign GEN_170 = T_2303 ? GEN_143 : wmask_buffer_1;
  assign GEN_171 = T_2303 ? GEN_144 : wmask_buffer_2;
  assign GEN_172 = T_2303 ? GEN_145 : wmask_buffer_3;
  assign GEN_173 = T_2303 ? GEN_146 : wmask_buffer_4;
  assign GEN_174 = T_2303 ? GEN_147 : wmask_buffer_5;
  assign GEN_175 = T_2303 ? GEN_148 : wmask_buffer_6;
  assign GEN_176 = T_2303 ? GEN_149 : wmask_buffer_7;
  assign T_2604_state = 2'h2;
  assign T_2631 = T_1653 | io_alloc_irel_should;
  assign T_2647 = T_2307 & T_2310;
  assign T_2648 = pending_orel_data | T_2647;
  assign T_2651 = io_outer_release_bits_r_type == 3'h0;
  assign T_2652 = io_outer_release_bits_r_type == 3'h1;
  assign T_2653 = io_outer_release_bits_r_type == 3'h2;
  assign T_2654 = T_2651 | T_2652;
  assign T_2655 = T_2654 | T_2653;
  assign T_2656 = T_2255 & T_2655;
  assign T_2660 = T_2656 ? 8'hff : 8'h0;
  assign T_2661 = ~ T_2660;
  assign T_2663 = 8'h1 << io_outer_release_bits_addr_beat;
  assign T_2664 = ~ T_2663;
  assign T_2665 = T_2661 | T_2664;
  assign T_2666 = T_2648 & T_2665;
  assign GEN_177 = T_2631 ? T_2666 : pending_orel_data;
  assign T_2677 = T_2655 == 1'h0;
  assign T_2679 = io_outer_release_bits_addr_beat == 3'h0;
  assign T_2680 = T_2677 | T_2679;
  assign GEN_179 = T_2680 ? 1'h1 : sending_orel;
  assign T_2692 = io_outer_release_bits_addr_beat == 3'h7;
  assign T_2693 = T_2677 | T_2692;
  assign GEN_180 = T_2693 ? 1'h0 : GEN_179;
  assign GEN_181 = T_2255 ? GEN_180 : sending_orel;
  assign GEN_182 = T_2255 ? 1'h0 : pending_orel_send;
  assign T_2702 = T_2255 & io_outer_release_bits_voluntary;
  assign T_2710 = T_2702 & T_2655;
  assign T_2714 = T_2712 == 3'h7;
  assign T_2716 = T_2712 + 3'h1;
  assign T_2717 = T_2716[2:0];
  assign GEN_183 = T_2710 ? T_2717 : T_2712;
  assign T_2718 = T_2710 & T_2714;
  assign T_2719 = T_2655 ? T_2712 : 3'h0;
  assign T_2720 = T_2655 ? T_2718 : T_2702;
  assign T_2723 = io_outer_grant_bits_g_type == 4'h0;
  assign T_2724 = io_outer_grant_bits_is_builtin_type & T_2723;
  assign T_2725 = T_2241 & T_2724;
  assign T_2733_0 = 3'h5;
  assign GEN_413 = {{1'd0}, T_2733_0};
  assign T_2735 = io_outer_grant_bits_g_type == GEN_413;
  assign T_2737 = io_outer_grant_bits_is_builtin_type ? T_2735 : T_2723;
  assign T_2739 = T_2725 & T_2737;
  assign T_2743 = T_2741 == 3'h7;
  assign T_2745 = T_2741 + 3'h1;
  assign T_2746 = T_2745[2:0];
  assign GEN_184 = T_2739 ? T_2746 : T_2741;
  assign T_2747 = T_2739 & T_2743;
  assign T_2748 = T_2737 ? T_2741 : 3'h0;
  assign T_2749 = T_2737 ? T_2747 : T_2725;
  assign T_2753 = T_2749 == 1'h0;
  assign T_2754 = T_2720 & T_2753;
  assign T_2756 = T_2751 + 1'h1;
  assign T_2757 = T_2756[0:0];
  assign GEN_185 = T_2754 ? T_2757 : T_2751;
  assign T_2759 = T_2720 == 1'h0;
  assign T_2760 = T_2749 & T_2759;
  assign T_2762 = T_2751 - 1'h1;
  assign T_2763 = T_2762[0:0];
  assign GEN_186 = T_2760 ? T_2763 : GEN_185;
  assign T_2765 = T_2751 > 1'h0;
  assign T_2774 = pending_orel_data >> vol_ognt_counter_up_idx;
  assign T_2775 = T_2774[0];
  assign T_2776 = T_2655 ? T_2775 : pending_orel_send;
  assign T_2777 = T_2337 & T_2776;
  assign T_2791 = T_2604_state == 2'h2;
  assign T_2792 = T_2791 ? 3'h0 : 3'h3;
  assign T_2828_addr_beat = vol_ognt_counter_up_idx;
  assign T_2828_addr_block = xact_addr_block;
  assign T_2828_client_xact_id = 3'h0;
  assign T_2828_voluntary = 1'h1;
  assign T_2828_r_type = T_2792;
  assign T_2828_data = GEN_11;
  assign GEN_11 = GEN_193;
  assign GEN_187 = 3'h1 == vol_ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_188 = 3'h2 == vol_ognt_counter_up_idx ? data_buffer_2 : GEN_187;
  assign GEN_189 = 3'h3 == vol_ognt_counter_up_idx ? data_buffer_3 : GEN_188;
  assign GEN_190 = 3'h4 == vol_ognt_counter_up_idx ? data_buffer_4 : GEN_189;
  assign GEN_191 = 3'h5 == vol_ognt_counter_up_idx ? data_buffer_5 : GEN_190;
  assign GEN_192 = 3'h6 == vol_ognt_counter_up_idx ? data_buffer_6 : GEN_191;
  assign GEN_193 = 3'h7 == vol_ognt_counter_up_idx ? data_buffer_7 : GEN_192;
  assign T_2857 = xact_iacq_is_builtin_type == 1'h0;
  assign T_2860 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2871_0 = 3'h3;
  assign T_2873 = io_outer_acquire_bits_a_type == T_2871_0;
  assign T_2874 = io_outer_acquire_bits_is_builtin_type & T_2873;
  assign T_2875 = T_2860 & T_2874;
  assign T_2879 = T_2877 == 3'h7;
  assign T_2881 = T_2877 + 3'h1;
  assign T_2882 = T_2881[2:0];
  assign GEN_195 = T_2875 ? T_2882 : T_2877;
  assign T_2883 = T_2875 & T_2879;
  assign T_2884 = T_2874 ? T_2877 : xact_addr_beat;
  assign T_2885 = T_2874 ? T_2883 : T_2860;
  assign T_2891 = T_2724 == 1'h0;
  assign T_2892 = T_2241 & T_2891;
  assign T_2900_0 = 3'h5;
  assign GEN_414 = {{1'd0}, T_2900_0};
  assign T_2902 = io_outer_grant_bits_g_type == GEN_414;
  assign T_2904 = io_outer_grant_bits_is_builtin_type ? T_2902 : T_2723;
  assign T_2906 = T_2892 & T_2904;
  assign T_2910 = T_2908 == 3'h7;
  assign T_2912 = T_2908 + 3'h1;
  assign T_2913 = T_2912[2:0];
  assign GEN_196 = T_2906 ? T_2913 : T_2908;
  assign T_2914 = T_2906 & T_2910;
  assign T_2915 = T_2904 ? T_2908 : xact_addr_beat;
  assign T_2916 = T_2904 ? T_2914 : T_2892;
  assign T_2920 = T_2916 == 1'h0;
  assign T_2921 = T_2885 & T_2920;
  assign T_2923 = T_2918 + 1'h1;
  assign T_2924 = T_2923[0:0];
  assign GEN_197 = T_2921 ? T_2924 : T_2918;
  assign T_2926 = T_2885 == 1'h0;
  assign T_2927 = T_2916 & T_2926;
  assign T_2929 = T_2918 - 1'h1;
  assign T_2930 = T_2929[0:0];
  assign GEN_198 = T_2927 ? T_2930 : GEN_197;
  assign T_2932 = T_2918 > 1'h0;
  assign T_2933 = state == 4'h6;
  assign T_2937 = pending_put_data >> ognt_counter_up_idx;
  assign T_2938 = T_2937[0];
  assign T_2940 = T_2938 == 1'h0;
  assign T_2949_0 = 3'h2;
  assign T_2949_1 = 3'h3;
  assign T_2949_2 = 3'h4;
  assign T_2967 = xact_allocate | T_2940;
  assign T_2968 = T_2933 & T_2967;
  assign T_2971 = xact_op_code == 5'h1;
  assign T_2972 = xact_op_code == 5'h7;
  assign T_2973 = T_2971 | T_2972;
  assign T_2974 = xact_op_code[3];
  assign T_2975 = xact_op_code == 5'h4;
  assign T_2976 = T_2974 | T_2975;
  assign T_2977 = T_2973 | T_2976;
  assign T_2978 = xact_op_code == 5'h3;
  assign T_2979 = T_2977 | T_2978;
  assign T_2980 = xact_op_code == 5'h6;
  assign T_2981 = T_2979 | T_2980;
  assign T_2984 = {xact_op_code,1'h1};
  assign T_3015_addr_block = xact_addr_block;
  assign T_3015_client_xact_id = 3'h0;
  assign T_3015_addr_beat = 3'h0;
  assign T_3015_is_builtin_type = 1'h0;
  assign T_3015_a_type = {{2'd0}, T_2981};
  assign T_3015_union = {{5'd0}, T_2984};
  assign T_3015_data = 64'h0;
  assign GEN_12 = GEN_205;
  assign GEN_199 = 3'h1 == ognt_counter_up_idx ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_200 = 3'h2 == ognt_counter_up_idx ? wmask_buffer_2 : GEN_199;
  assign GEN_201 = 3'h3 == ognt_counter_up_idx ? wmask_buffer_3 : GEN_200;
  assign GEN_202 = 3'h4 == ognt_counter_up_idx ? wmask_buffer_4 : GEN_201;
  assign GEN_203 = 3'h5 == ognt_counter_up_idx ? wmask_buffer_5 : GEN_202;
  assign GEN_204 = 3'h6 == ognt_counter_up_idx ? wmask_buffer_6 : GEN_203;
  assign GEN_205 = 3'h7 == ognt_counter_up_idx ? wmask_buffer_7 : GEN_204;
  assign T_3080 = {xact_op_code,1'h0};
  assign T_3081 = {xact_addr_byte,xact_op_size};
  assign T_3082 = {T_3081,T_3080};
  assign T_3084 = {xact_op_size,xact_op_code};
  assign T_3085 = {T_3084,1'h0};
  assign T_3087 = {GEN_12,1'h0};
  assign T_3099 = T_1993 ? 6'h2 : 6'h0;
  assign T_3101 = T_1995 ? 6'h0 : T_3099;
  assign T_3103 = T_1991 ? T_3082 : {{5'd0}, T_3101};
  assign T_3105 = T_2001 ? {{2'd0}, T_3087} : T_3103;
  assign T_3107 = T_1997 ? {{2'd0}, T_3087} : T_3105;
  assign T_3109 = T_2003 ? {{3'd0}, T_3085} : T_3107;
  assign T_3111 = T_1999 ? T_3082 : T_3109;
  assign T_3140_addr_block = xact_addr_block;
  assign T_3140_client_xact_id = 3'h0;
  assign T_3140_addr_beat = ognt_counter_up_idx;
  assign T_3140_is_builtin_type = 1'h1;
  assign T_3140_a_type = xact_iacq_a_type;
  assign T_3140_union = T_3111;
  assign T_3140_data = GEN_13;
  assign GEN_13 = GEN_212;
  assign GEN_206 = 3'h1 == ognt_counter_up_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_207 = 3'h2 == ognt_counter_up_idx ? data_buffer_2 : GEN_206;
  assign GEN_208 = 3'h3 == ognt_counter_up_idx ? data_buffer_3 : GEN_207;
  assign GEN_209 = 3'h4 == ognt_counter_up_idx ? data_buffer_4 : GEN_208;
  assign GEN_210 = 3'h5 == ognt_counter_up_idx ? data_buffer_5 : GEN_209;
  assign GEN_211 = 3'h6 == ognt_counter_up_idx ? data_buffer_6 : GEN_210;
  assign GEN_212 = 3'h7 == ognt_counter_up_idx ? data_buffer_7 : GEN_211;
  assign T_3168_addr_block = T_2857 ? T_3015_addr_block : T_3140_addr_block;
  assign T_3168_client_xact_id = T_2857 ? T_3015_client_xact_id : T_3140_client_xact_id;
  assign T_3168_addr_beat = T_2857 ? T_3015_addr_beat : T_3140_addr_beat;
  assign T_3168_is_builtin_type = T_2857 ? T_3015_is_builtin_type : T_3140_is_builtin_type;
  assign T_3168_a_type = T_2857 ? T_3015_a_type : T_3140_a_type;
  assign T_3168_union = T_2857 ? T_3015_union : T_3140_union;
  assign T_3168_data = T_2857 ? T_3015_data : T_3140_data;
  assign T_3197 = T_2933 & ognt_counter_up_done;
  assign GEN_213 = T_3197 ? 4'h7 : GEN_58;
  assign GEN_214 = ognt_counter_pending ? 1'h1 : vol_ognt_counter_pending;
  assign T_3207_0 = 3'h5;
  assign T_3207_1 = 3'h4;
  assign GEN_415 = {{1'd0}, T_3207_0};
  assign T_3209 = io_outer_grant_bits_g_type == GEN_415;
  assign GEN_416 = {{1'd0}, T_3207_1};
  assign T_3210 = io_outer_grant_bits_g_type == GEN_416;
  assign T_3211 = T_3209 | T_3210;
  assign T_3213 = io_outer_grant_bits_is_builtin_type ? T_3211 : T_2723;
  assign T_3214 = T_2241 & T_3213;
  assign GEN_14 = GEN_221;
  assign GEN_215 = 3'h1 == io_outer_grant_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_216 = 3'h2 == io_outer_grant_bits_addr_beat ? wmask_buffer_2 : GEN_215;
  assign GEN_217 = 3'h3 == io_outer_grant_bits_addr_beat ? wmask_buffer_3 : GEN_216;
  assign GEN_218 = 3'h4 == io_outer_grant_bits_addr_beat ? wmask_buffer_4 : GEN_217;
  assign GEN_219 = 3'h5 == io_outer_grant_bits_addr_beat ? wmask_buffer_5 : GEN_218;
  assign GEN_220 = 3'h6 == io_outer_grant_bits_addr_beat ? wmask_buffer_6 : GEN_219;
  assign GEN_221 = 3'h7 == io_outer_grant_bits_addr_beat ? wmask_buffer_7 : GEN_220;
  assign T_3215 = GEN_14[0];
  assign GEN_15 = GEN_221;
  assign T_3216 = GEN_15[1];
  assign GEN_16 = GEN_221;
  assign T_3217 = GEN_16[2];
  assign GEN_17 = GEN_221;
  assign T_3218 = GEN_17[3];
  assign GEN_18 = GEN_221;
  assign T_3219 = GEN_18[4];
  assign GEN_19 = GEN_221;
  assign T_3220 = GEN_19[5];
  assign GEN_20 = GEN_221;
  assign T_3221 = GEN_20[6];
  assign GEN_21 = GEN_221;
  assign T_3222 = GEN_21[7];
  assign T_3226 = T_3215 ? 8'hff : 8'h0;
  assign T_3230 = T_3216 ? 8'hff : 8'h0;
  assign T_3234 = T_3217 ? 8'hff : 8'h0;
  assign T_3238 = T_3218 ? 8'hff : 8'h0;
  assign T_3242 = T_3219 ? 8'hff : 8'h0;
  assign T_3246 = T_3220 ? 8'hff : 8'h0;
  assign T_3250 = T_3221 ? 8'hff : 8'h0;
  assign T_3254 = T_3222 ? 8'hff : 8'h0;
  assign T_3255 = {T_3230,T_3226};
  assign T_3256 = {T_3238,T_3234};
  assign T_3257 = {T_3256,T_3255};
  assign T_3258 = {T_3246,T_3242};
  assign T_3259 = {T_3254,T_3250};
  assign T_3260 = {T_3259,T_3258};
  assign T_3261 = {T_3260,T_3257};
  assign T_3262 = ~ T_3261;
  assign T_3263 = T_3262 & io_outer_grant_bits_data;
  assign GEN_22 = GEN_277;
  assign GEN_271 = 3'h1 == io_outer_grant_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_272 = 3'h2 == io_outer_grant_bits_addr_beat ? data_buffer_2 : GEN_271;
  assign GEN_273 = 3'h3 == io_outer_grant_bits_addr_beat ? data_buffer_3 : GEN_272;
  assign GEN_274 = 3'h4 == io_outer_grant_bits_addr_beat ? data_buffer_4 : GEN_273;
  assign GEN_275 = 3'h5 == io_outer_grant_bits_addr_beat ? data_buffer_5 : GEN_274;
  assign GEN_276 = 3'h6 == io_outer_grant_bits_addr_beat ? data_buffer_6 : GEN_275;
  assign GEN_277 = 3'h7 == io_outer_grant_bits_addr_beat ? data_buffer_7 : GEN_276;
  assign T_3264 = T_3261 & GEN_22;
  assign T_3265 = T_3263 | T_3264;
  assign GEN_23 = T_3265;
  assign GEN_278 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_160;
  assign GEN_279 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_161;
  assign GEN_280 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_162;
  assign GEN_281 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_163;
  assign GEN_282 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_164;
  assign GEN_283 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_165;
  assign GEN_284 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_166;
  assign GEN_285 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_23 : GEN_167;
  assign GEN_24 = 8'hff;
  assign GEN_286 = 3'h0 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_169;
  assign GEN_287 = 3'h1 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_170;
  assign GEN_288 = 3'h2 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_171;
  assign GEN_289 = 3'h3 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_172;
  assign GEN_290 = 3'h4 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_173;
  assign GEN_291 = 3'h5 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_174;
  assign GEN_292 = 3'h6 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_175;
  assign GEN_293 = 3'h7 == io_outer_grant_bits_addr_beat ? GEN_24 : GEN_176;
  assign GEN_304 = T_3214 ? GEN_278 : GEN_160;
  assign GEN_305 = T_3214 ? GEN_279 : GEN_161;
  assign GEN_306 = T_3214 ? GEN_280 : GEN_162;
  assign GEN_307 = T_3214 ? GEN_281 : GEN_163;
  assign GEN_308 = T_3214 ? GEN_282 : GEN_164;
  assign GEN_309 = T_3214 ? GEN_283 : GEN_165;
  assign GEN_310 = T_3214 ? GEN_284 : GEN_166;
  assign GEN_311 = T_3214 ? GEN_285 : GEN_167;
  assign GEN_313 = T_3214 ? GEN_286 : GEN_169;
  assign GEN_314 = T_3214 ? GEN_287 : GEN_170;
  assign GEN_315 = T_3214 ? GEN_288 : GEN_171;
  assign GEN_316 = T_3214 ? GEN_289 : GEN_172;
  assign GEN_317 = T_3214 ? GEN_290 : GEN_173;
  assign GEN_318 = T_3214 ? GEN_291 : GEN_174;
  assign GEN_319 = T_3214 ? GEN_292 : GEN_175;
  assign GEN_320 = T_3214 ? GEN_293 : GEN_176;
  assign T_3268 = scoreboard_3 | ognt_counter_pending;
  assign T_3269 = T_3268 | vol_ognt_counter_pending;
  assign T_3281 = T_2179 == 1'h0;
  assign T_3283 = T_2175 & T_3281;
  assign T_3291_0 = 3'h5;
  assign GEN_417 = {{1'd0}, T_3291_0};
  assign T_3293 = io_inner_grant_bits_g_type == GEN_417;
  assign T_3295 = io_inner_grant_bits_is_builtin_type ? T_3293 : T_2178;
  assign T_3297 = T_3283 & T_3295;
  assign T_3301 = T_3299 == 3'h7;
  assign T_3303 = T_3299 + 3'h1;
  assign T_3304 = T_3303[2:0];
  assign GEN_321 = T_3297 ? T_3304 : T_3299;
  assign T_3305 = T_3297 & T_3301;
  assign T_3306 = T_3295 ? T_3299 : 3'h0;
  assign T_3307 = T_3295 ? T_3305 : T_3283;
  assign T_3308 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_3326 = T_3308 == 1'h0;
  assign T_3327 = T_3307 & T_3326;
  assign T_3329 = T_3324 + 1'h1;
  assign T_3330 = T_3329[0:0];
  assign GEN_323 = T_3327 ? T_3330 : T_3324;
  assign T_3332 = T_3307 == 1'h0;
  assign T_3333 = T_3308 & T_3332;
  assign T_3335 = T_3324 - 1'h1;
  assign T_3336 = T_3335[0:0];
  assign GEN_324 = T_3333 ? T_3336 : GEN_323;
  assign T_3338 = T_3324 > 1'h0;
  assign T_3343 = T_1798 == 1'h0;
  assign T_3360 = pending_ignt_data | T_2647;
  assign T_3370_0 = 3'h5;
  assign T_3370_1 = 3'h4;
  assign GEN_418 = {{1'd0}, T_3370_0};
  assign T_3372 = io_outer_grant_bits_g_type == GEN_418;
  assign GEN_419 = {{1'd0}, T_3370_1};
  assign T_3373 = io_outer_grant_bits_g_type == GEN_419;
  assign T_3374 = T_3372 | T_3373;
  assign T_3376 = io_outer_grant_bits_is_builtin_type ? T_3374 : T_2723;
  assign T_3377 = T_2241 & T_3376;
  assign T_3382 = T_3377 ? 8'hff : 8'h0;
  assign T_3384 = 8'h1 << io_outer_grant_bits_addr_beat;
  assign T_3385 = T_3382 & T_3384;
  assign T_3386 = T_3360 | T_3385;
  assign GEN_327 = T_3343 ? T_3386 : GEN_45;
  assign T_3389 = state == 4'h1;
  assign T_3390 = T_1611 | T_3389;
  assign T_3393 = T_3390 | scoreboard_0;
  assign T_3395 = T_3393 == 1'h0;
  assign T_3412 = 3'h6 == ignt_q_io_deq_bits_a_type;
  assign T_3413 = T_3412 ? 3'h1 : 3'h3;
  assign T_3414 = 3'h5 == ignt_q_io_deq_bits_a_type;
  assign T_3415 = T_3414 ? 3'h1 : T_3413;
  assign T_3416 = 3'h4 == ignt_q_io_deq_bits_a_type;
  assign T_3417 = T_3416 ? 3'h4 : T_3415;
  assign T_3418 = 3'h3 == ignt_q_io_deq_bits_a_type;
  assign T_3419 = T_3418 ? 3'h3 : T_3417;
  assign T_3420 = 3'h2 == ignt_q_io_deq_bits_a_type;
  assign T_3421 = T_3420 ? 3'h3 : T_3419;
  assign T_3422 = 3'h1 == ignt_q_io_deq_bits_a_type;
  assign T_3423 = T_3422 ? 3'h5 : T_3421;
  assign T_3424 = 3'h0 == ignt_q_io_deq_bits_a_type;
  assign T_3425 = T_3424 ? 3'h4 : T_3423;
  assign T_3426 = ignt_q_io_deq_bits_is_builtin_type ? T_3425 : 3'h0;
  assign T_3455_addr_beat = ignt_q_io_deq_bits_addr_beat;
  assign T_3455_client_xact_id = ignt_q_io_deq_bits_client_xact_id;
  assign T_3455_manager_xact_id = 3'h4;
  assign T_3455_is_builtin_type = ignt_q_io_deq_bits_is_builtin_type;
  assign T_3455_g_type = {{1'd0}, T_3426};
  assign T_3455_data = GEN_25;
  assign T_3455_client_id = ignt_q_io_deq_bits_client_id;
  assign GEN_25 = GEN_334;
  assign GEN_328 = 3'h1 == ignt_data_idx ? data_buffer_1 : data_buffer_0;
  assign GEN_329 = 3'h2 == ignt_data_idx ? data_buffer_2 : GEN_328;
  assign GEN_330 = 3'h3 == ignt_data_idx ? data_buffer_3 : GEN_329;
  assign GEN_331 = 3'h4 == ignt_data_idx ? data_buffer_4 : GEN_330;
  assign GEN_332 = 3'h5 == ignt_data_idx ? data_buffer_5 : GEN_331;
  assign GEN_333 = 3'h6 == ignt_data_idx ? data_buffer_6 : GEN_332;
  assign GEN_334 = 3'h7 == ignt_data_idx ? data_buffer_7 : GEN_333;
  assign T_3491_0 = 3'h5;
  assign GEN_420 = {{1'd0}, T_3491_0};
  assign T_3493 = io_inner_grant_bits_g_type == GEN_420;
  assign T_3495 = io_inner_grant_bits_is_builtin_type ? T_3493 : T_2178;
  assign T_3497 = T_2175 & T_3495;
  assign T_3501 = T_3499 == 3'h7;
  assign T_3503 = T_3499 + 3'h1;
  assign T_3504 = T_3503[2:0];
  assign GEN_335 = T_3497 ? T_3504 : T_3499;
  assign T_3505 = T_3497 & T_3501;
  assign T_3506 = T_3495 ? T_3499 : ignt_q_io_deq_bits_addr_beat;
  assign T_3507 = T_3495 ? T_3505 : T_2175;
  assign T_3512 = T_2337 & scoreboard_6;
  assign T_3514 = T_3269 == 1'h0;
  assign T_3522_0 = 3'h5;
  assign T_3522_1 = 3'h4;
  assign GEN_421 = {{1'd0}, T_3522_0};
  assign T_3524 = io_inner_grant_bits_g_type == GEN_421;
  assign GEN_422 = {{1'd0}, T_3522_1};
  assign T_3525 = io_inner_grant_bits_g_type == GEN_422;
  assign T_3526 = T_3524 | T_3525;
  assign T_3528 = io_inner_grant_bits_is_builtin_type ? T_3526 : T_2178;
  assign T_3529 = pending_ignt_data >> ignt_data_idx;
  assign T_3530 = T_3529[0];
  assign T_3532 = T_3528 ? T_3530 : T_3395;
  assign T_3533 = T_3514 & T_3532;
  assign GEN_338 = T_3512 ? T_3533 : T_2347;
  assign GEN_339 = T_2250 ? ignt_data_done : 1'h0;
  assign GEN_340 = T_2250 ? ignt_data_idx : T_2440_addr_beat;
  assign GEN_341 = T_2250 ? T_3455_client_xact_id : T_2440_client_xact_id;
  assign GEN_342 = T_2250 ? T_3455_manager_xact_id : T_2440_manager_xact_id;
  assign GEN_343 = T_2250 ? T_3455_is_builtin_type : T_2440_is_builtin_type;
  assign GEN_344 = T_2250 ? T_3455_g_type : T_2440_g_type;
  assign GEN_345 = T_2250 ? T_3455_data : T_2440_data;
  assign GEN_346 = T_2250 ? T_3455_client_id : T_2440_client_id;
  assign GEN_349 = T_2250 ? GEN_338 : T_2347;
  assign T_3540 = ~ io_incoherent_0;
  assign GEN_350 = T_1798 ? {{1'd0}, T_3540} : T_2079;
  assign T_3551 = T_1767 & io_inner_acquire_valid;
  assign T_3552 = T_1798 | T_3551;
  assign T_3562_0 = 3'h2;
  assign T_3562_1 = 3'h3;
  assign T_3562_2 = 3'h4;
  assign T_3564 = io_inner_acquire_bits_a_type == T_3562_0;
  assign T_3565 = io_inner_acquire_bits_a_type == T_3562_1;
  assign T_3566 = io_inner_acquire_bits_a_type == T_3562_2;
  assign T_3567 = T_3564 | T_3565;
  assign T_3568 = T_3567 | T_3566;
  assign T_3569 = io_inner_acquire_bits_is_builtin_type & T_3568;
  assign T_3570 = T_1612 & T_3569;
  assign T_3571 = T_3570 & T_3552;
  assign T_3573 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_3574 = io_inner_acquire_bits_is_builtin_type & T_3573;
  assign T_3603 = T_1921 | T_1918;
  assign T_3604 = io_inner_acquire_bits_union[8:1];
  assign T_3606 = T_3603 ? T_3604 : 8'h0;
  assign T_3607 = T_3574 ? 8'hff : T_3606;
  assign T_3608 = T_3607[0];
  assign T_3609 = T_3607[1];
  assign T_3610 = T_3607[2];
  assign T_3611 = T_3607[3];
  assign T_3612 = T_3607[4];
  assign T_3613 = T_3607[5];
  assign T_3614 = T_3607[6];
  assign T_3615 = T_3607[7];
  assign T_3619 = T_3608 ? 8'hff : 8'h0;
  assign T_3623 = T_3609 ? 8'hff : 8'h0;
  assign T_3627 = T_3610 ? 8'hff : 8'h0;
  assign T_3631 = T_3611 ? 8'hff : 8'h0;
  assign T_3635 = T_3612 ? 8'hff : 8'h0;
  assign T_3639 = T_3613 ? 8'hff : 8'h0;
  assign T_3643 = T_3614 ? 8'hff : 8'h0;
  assign T_3647 = T_3615 ? 8'hff : 8'h0;
  assign T_3648 = {T_3623,T_3619};
  assign T_3649 = {T_3631,T_3627};
  assign T_3650 = {T_3649,T_3648};
  assign T_3651 = {T_3639,T_3635};
  assign T_3652 = {T_3647,T_3643};
  assign T_3653 = {T_3652,T_3651};
  assign T_3654 = {T_3653,T_3650};
  assign T_3655 = ~ T_3654;
  assign GEN_26 = GEN_357;
  assign GEN_351 = 3'h1 == io_inner_acquire_bits_addr_beat ? data_buffer_1 : data_buffer_0;
  assign GEN_352 = 3'h2 == io_inner_acquire_bits_addr_beat ? data_buffer_2 : GEN_351;
  assign GEN_353 = 3'h3 == io_inner_acquire_bits_addr_beat ? data_buffer_3 : GEN_352;
  assign GEN_354 = 3'h4 == io_inner_acquire_bits_addr_beat ? data_buffer_4 : GEN_353;
  assign GEN_355 = 3'h5 == io_inner_acquire_bits_addr_beat ? data_buffer_5 : GEN_354;
  assign GEN_356 = 3'h6 == io_inner_acquire_bits_addr_beat ? data_buffer_6 : GEN_355;
  assign GEN_357 = 3'h7 == io_inner_acquire_bits_addr_beat ? data_buffer_7 : GEN_356;
  assign T_3656 = T_3655 & GEN_26;
  assign T_3657 = T_3654 & io_inner_acquire_bits_data;
  assign T_3658 = T_3656 | T_3657;
  assign GEN_27 = T_3658;
  assign GEN_358 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_304;
  assign GEN_359 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_305;
  assign GEN_360 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_306;
  assign GEN_361 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_307;
  assign GEN_362 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_308;
  assign GEN_363 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_309;
  assign GEN_364 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_310;
  assign GEN_365 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_27 : GEN_311;
  assign GEN_28 = GEN_372;
  assign GEN_366 = 3'h1 == io_inner_acquire_bits_addr_beat ? wmask_buffer_1 : wmask_buffer_0;
  assign GEN_367 = 3'h2 == io_inner_acquire_bits_addr_beat ? wmask_buffer_2 : GEN_366;
  assign GEN_368 = 3'h3 == io_inner_acquire_bits_addr_beat ? wmask_buffer_3 : GEN_367;
  assign GEN_369 = 3'h4 == io_inner_acquire_bits_addr_beat ? wmask_buffer_4 : GEN_368;
  assign GEN_370 = 3'h5 == io_inner_acquire_bits_addr_beat ? wmask_buffer_5 : GEN_369;
  assign GEN_371 = 3'h6 == io_inner_acquire_bits_addr_beat ? wmask_buffer_6 : GEN_370;
  assign GEN_372 = 3'h7 == io_inner_acquire_bits_addr_beat ? wmask_buffer_7 : GEN_371;
  assign T_3695 = T_3607 | GEN_28;
  assign GEN_29 = T_3695;
  assign GEN_373 = 3'h0 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_313;
  assign GEN_374 = 3'h1 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_314;
  assign GEN_375 = 3'h2 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_315;
  assign GEN_376 = 3'h3 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_316;
  assign GEN_377 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_317;
  assign GEN_378 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_318;
  assign GEN_379 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_319;
  assign GEN_380 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_29 : GEN_320;
  assign GEN_383 = T_3571 ? GEN_358 : GEN_304;
  assign GEN_384 = T_3571 ? GEN_359 : GEN_305;
  assign GEN_385 = T_3571 ? GEN_360 : GEN_306;
  assign GEN_386 = T_3571 ? GEN_361 : GEN_307;
  assign GEN_387 = T_3571 ? GEN_362 : GEN_308;
  assign GEN_388 = T_3571 ? GEN_363 : GEN_309;
  assign GEN_389 = T_3571 ? GEN_364 : GEN_310;
  assign GEN_390 = T_3571 ? GEN_365 : GEN_311;
  assign GEN_393 = T_3571 ? GEN_373 : GEN_313;
  assign GEN_394 = T_3571 ? GEN_374 : GEN_314;
  assign GEN_395 = T_3571 ? GEN_375 : GEN_315;
  assign GEN_396 = T_3571 ? GEN_376 : GEN_316;
  assign GEN_397 = T_3571 ? GEN_377 : GEN_317;
  assign GEN_398 = T_3571 ? GEN_378 : GEN_318;
  assign GEN_399 = T_3571 ? GEN_379 : GEN_319;
  assign GEN_400 = T_3571 ? GEN_380 : GEN_320;
  assign T_3698 = scoreboard_0 | T_2343;
  assign T_3699 = T_3698 | vol_ignt_counter_pending;
  assign T_3700 = T_3699 | scoreboard_3;
  assign T_3701 = T_3700 | vol_ognt_counter_pending;
  assign T_3702 = T_3701 | ognt_counter_pending;
  assign T_3703 = T_3702 | scoreboard_6;
  assign T_3704 = T_3703 | ifin_counter_pending;
  assign T_3706 = T_3704 == 1'h0;
  assign T_3708 = T_2337 & all_pending_done;
  assign GEN_401 = T_3708 ? 4'h0 : GEN_213;
  assign GEN_402 = T_3708 ? 8'h0 : GEN_393;
  assign GEN_403 = T_3708 ? 8'h0 : GEN_394;
  assign GEN_404 = T_3708 ? 8'h0 : GEN_395;
  assign GEN_405 = T_3708 ? 8'h0 : GEN_396;
  assign GEN_406 = T_3708 ? 8'h0 : GEN_397;
  assign GEN_407 = T_3708 ? 8'h0 : GEN_398;
  assign GEN_408 = T_3708 ? 8'h0 : GEN_399;
  assign GEN_409 = T_3708 ? 8'h0 : GEN_400;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_30 = GEN_121[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_31 = GEN_122[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  state = GEN_32[3:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  xact_addr_block = GEN_33[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_41 = {1{$random}};
  xact_allocate = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_42 = {1{$random}};
  xact_amo_shift_bytes = GEN_42[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  xact_op_code = GEN_43[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_addr_byte = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_78 = {1{$random}};
  xact_op_size = GEN_78[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_79 = {1{$random}};
  xact_vol_ir_r_type = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_80 = {1{$random}};
  xact_vol_ir_src = GEN_80[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_81 = {1{$random}};
  xact_vol_ir_client_xact_id = GEN_81[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_82 = {1{$random}};
  pending_irel_data = GEN_82[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_83 = {1{$random}};
  pending_put_data = GEN_83[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_84 = {1{$random}};
  pending_ignt_data = GEN_84[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  pending_iprbs = GEN_85[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  pending_orel_send = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_87 = {1{$random}};
  pending_orel_data = GEN_87[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  sending_orel = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {2{$random}};
  data_buffer_0 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {2{$random}};
  data_buffer_1 = GEN_90[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_91 = {2{$random}};
  data_buffer_2 = GEN_91[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_92 = {2{$random}};
  data_buffer_3 = GEN_92[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_93 = {2{$random}};
  data_buffer_4 = GEN_93[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_94 = {2{$random}};
  data_buffer_5 = GEN_94[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_95 = {2{$random}};
  data_buffer_6 = GEN_95[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_96 = {2{$random}};
  data_buffer_7 = GEN_96[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_97 = {1{$random}};
  wmask_buffer_0 = GEN_97[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_98 = {1{$random}};
  wmask_buffer_1 = GEN_98[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_99 = {1{$random}};
  wmask_buffer_2 = GEN_99[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_100 = {1{$random}};
  wmask_buffer_3 = GEN_100[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_101 = {1{$random}};
  wmask_buffer_4 = GEN_101[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_102 = {1{$random}};
  wmask_buffer_5 = GEN_102[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_103 = {1{$random}};
  wmask_buffer_6 = GEN_103[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_104 = {1{$random}};
  wmask_buffer_7 = GEN_104[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_105 = {1{$random}};
  T_2091 = GEN_105[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_106 = {1{$random}};
  T_2115 = GEN_106[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_107 = {1{$random}};
  T_2125 = GEN_107[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_108 = {1{$random}};
  T_2166 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  T_2197 = GEN_109[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  T_2207 = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_111 = {1{$random}};
  T_2712 = GEN_111[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  T_2741 = GEN_112[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {1{$random}};
  T_2751 = GEN_113[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  T_2877 = GEN_114[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  T_2908 = GEN_115[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  T_2918 = GEN_116[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  T_3299 = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  T_3314 = GEN_118[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  T_3324 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  T_3499 = GEN_120[2:0];
  `endif
  GEN_121 = {1{$random}};
  GEN_122 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      if(T_3708) begin
        state <= 4'h0;
      end else begin
        if(T_3197) begin
          state <= 4'h7;
        end else begin
          if(T_2224) begin
            state <= 4'h7;
          end else begin
            if(T_2146) begin
              if(T_2055) begin
                state <= 4'h6;
              end else begin
                state <= 4'h7;
              end
            end else begin
              if(T_1798) begin
                state <= 4'h5;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_addr_block <= 26'h0;
    end else begin
      if(T_2224) begin
        xact_addr_block <= io_inner_release_bits_addr_block;
      end else begin
        if(T_1798) begin
          xact_addr_block <= io_inner_acquire_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_allocate <= 1'h0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_amo_shift_bytes <= T_1915;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        if(T_1922) begin
          xact_op_code <= 5'h1;
        end else begin
          xact_op_code <= T_1923;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_addr_byte <= T_1925;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1798) begin
        xact_op_size <= T_1926;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_r_type <= io_inner_release_bits_r_type;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_src <= io_inner_release_bits_client_id;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2277) begin
        if(T_2289) begin
          if(io_inner_release_bits_voluntary) begin
            xact_vol_ir_client_xact_id <= io_inner_release_bits_client_xact_id;
          end
        end
      end
    end
    if(reset) begin
      pending_irel_data <= 8'h0;
    end else begin
      if(T_2277) begin
        if(T_2316) begin
          pending_irel_data <= T_2333;
        end else begin
          if(T_2289) begin
            if(T_2111) begin
              pending_irel_data <= T_2312;
            end else begin
              pending_irel_data <= 8'h0;
            end
          end else begin
            if(T_2224) begin
              pending_irel_data <= 8'hff;
            end
          end
        end
      end else begin
        if(T_2224) begin
          pending_irel_data <= 8'hff;
        end
      end
    end
    if(reset) begin
      pending_put_data <= 8'h0;
    end else begin
      if(T_1798) begin
        if(T_1921) begin
          pending_put_data <= T_1956;
        end else begin
          pending_put_data <= 8'h0;
        end
      end else begin
        if(T_1852) begin
          pending_put_data <= T_1907;
        end
      end
    end
    if(reset) begin
      pending_ignt_data <= 8'h0;
    end else begin
      if(T_3343) begin
        pending_ignt_data <= T_3386;
      end else begin
        if(T_1798) begin
          pending_ignt_data <= 8'h0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      pending_iprbs <= GEN_350[0];
    end
    if(reset) begin
      pending_orel_send <= 1'h0;
    end else begin
      if(T_2255) begin
        pending_orel_send <= 1'h0;
      end
    end
    if(reset) begin
      pending_orel_data <= 8'h0;
    end else begin
      if(T_2631) begin
        pending_orel_data <= T_2666;
      end
    end
    if(reset) begin
      sending_orel <= 1'h0;
    end else begin
      if(T_2255) begin
        if(T_2693) begin
          sending_orel <= 1'h0;
        end else begin
          if(T_2680) begin
            sending_orel <= 1'h1;
          end
        end
      end
    end
    if(reset) begin
      data_buffer_0 <= T_1691_0;
    end else begin
      if(T_3571) begin
        if(3'h0 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_0 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              data_buffer_0 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  data_buffer_0 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h0 == io_outer_grant_bits_addr_beat) begin
            data_buffer_0 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                data_buffer_0 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h0 == io_inner_release_bits_addr_beat) begin
              data_buffer_0 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_1 <= T_1691_1;
    end else begin
      if(T_3571) begin
        if(3'h1 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_1 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              data_buffer_1 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  data_buffer_1 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h1 == io_outer_grant_bits_addr_beat) begin
            data_buffer_1 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                data_buffer_1 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h1 == io_inner_release_bits_addr_beat) begin
              data_buffer_1 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_2 <= T_1691_2;
    end else begin
      if(T_3571) begin
        if(3'h2 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_2 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              data_buffer_2 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  data_buffer_2 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h2 == io_outer_grant_bits_addr_beat) begin
            data_buffer_2 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                data_buffer_2 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h2 == io_inner_release_bits_addr_beat) begin
              data_buffer_2 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_3 <= T_1691_3;
    end else begin
      if(T_3571) begin
        if(3'h3 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_3 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              data_buffer_3 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  data_buffer_3 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h3 == io_outer_grant_bits_addr_beat) begin
            data_buffer_3 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                data_buffer_3 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h3 == io_inner_release_bits_addr_beat) begin
              data_buffer_3 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_4 <= T_1691_4;
    end else begin
      if(T_3571) begin
        if(3'h4 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_4 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              data_buffer_4 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  data_buffer_4 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h4 == io_outer_grant_bits_addr_beat) begin
            data_buffer_4 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                data_buffer_4 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h4 == io_inner_release_bits_addr_beat) begin
              data_buffer_4 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_5 <= T_1691_5;
    end else begin
      if(T_3571) begin
        if(3'h5 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_5 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              data_buffer_5 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  data_buffer_5 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h5 == io_outer_grant_bits_addr_beat) begin
            data_buffer_5 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                data_buffer_5 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h5 == io_inner_release_bits_addr_beat) begin
              data_buffer_5 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_6 <= T_1691_6;
    end else begin
      if(T_3571) begin
        if(3'h6 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_6 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              data_buffer_6 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  data_buffer_6 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h6 == io_outer_grant_bits_addr_beat) begin
            data_buffer_6 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                data_buffer_6 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h6 == io_inner_release_bits_addr_beat) begin
              data_buffer_6 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      data_buffer_7 <= T_1691_7;
    end else begin
      if(T_3571) begin
        if(3'h7 == io_inner_acquire_bits_addr_beat) begin
          data_buffer_7 <= GEN_27;
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              data_buffer_7 <= GEN_23;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  data_buffer_7 <= GEN_9;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end
      end else begin
        if(T_3214) begin
          if(3'h7 == io_outer_grant_bits_addr_beat) begin
            data_buffer_7 <= GEN_23;
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                data_buffer_7 <= GEN_9;
              end
            end
          end
        end else begin
          if(T_2303) begin
            if(3'h7 == io_inner_release_bits_addr_beat) begin
              data_buffer_7 <= GEN_9;
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_0 <= T_1709_0;
    end else begin
      if(T_3708) begin
        wmask_buffer_0 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h0 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_0 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h0 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h0 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_0 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h0 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_0 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h0 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_0 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h0 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_0 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_1 <= T_1709_1;
    end else begin
      if(T_3708) begin
        wmask_buffer_1 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h1 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_1 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h1 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h1 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_1 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h1 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_1 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h1 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_1 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h1 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_1 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_2 <= T_1709_2;
    end else begin
      if(T_3708) begin
        wmask_buffer_2 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h2 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_2 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h2 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h2 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_2 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h2 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_2 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h2 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_2 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h2 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_2 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_3 <= T_1709_3;
    end else begin
      if(T_3708) begin
        wmask_buffer_3 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h3 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_3 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h3 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h3 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_3 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h3 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_3 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h3 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_3 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h3 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_3 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_4 <= T_1709_4;
    end else begin
      if(T_3708) begin
        wmask_buffer_4 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h4 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_4 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h4 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h4 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_4 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h4 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_4 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h4 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_4 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h4 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_4 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_5 <= T_1709_5;
    end else begin
      if(T_3708) begin
        wmask_buffer_5 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h5 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_5 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h5 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h5 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_5 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h5 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_5 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h5 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_5 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h5 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_5 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_6 <= T_1709_6;
    end else begin
      if(T_3708) begin
        wmask_buffer_6 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h6 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_6 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h6 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h6 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_6 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h6 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_6 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h6 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_6 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h6 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_6 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      wmask_buffer_7 <= T_1709_7;
    end else begin
      if(T_3708) begin
        wmask_buffer_7 <= 8'h0;
      end else begin
        if(T_3571) begin
          if(3'h7 == io_inner_acquire_bits_addr_beat) begin
            wmask_buffer_7 <= GEN_29;
          end else begin
            if(T_3214) begin
              if(3'h7 == io_outer_grant_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_24;
              end else begin
                if(T_2303) begin
                  if(3'h7 == io_inner_release_bits_addr_beat) begin
                    wmask_buffer_7 <= GEN_10;
                  end
                end
              end
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end
        end else begin
          if(T_3214) begin
            if(3'h7 == io_outer_grant_bits_addr_beat) begin
              wmask_buffer_7 <= GEN_24;
            end else begin
              if(T_2303) begin
                if(3'h7 == io_inner_release_bits_addr_beat) begin
                  wmask_buffer_7 <= GEN_10;
                end
              end
            end
          end else begin
            if(T_2303) begin
              if(3'h7 == io_inner_release_bits_addr_beat) begin
                wmask_buffer_7 <= GEN_10;
              end
            end
          end
        end
      end
    end
    if(reset) begin
      T_2091 <= 3'h0;
    end
    if(reset) begin
      T_2115 <= 3'h0;
    end else begin
      if(T_2113) begin
        T_2115 <= T_2120;
      end
    end
    if(reset) begin
      T_2125 <= 1'h0;
    end else begin
      if(T_2134) begin
        T_2125 <= T_2137;
      end else begin
        if(T_2128) begin
          T_2125 <= T_2131;
        end
      end
    end
    if(reset) begin
      T_2166 <= 3'h0;
    end else begin
      if(T_2164) begin
        T_2166 <= T_2171;
      end
    end
    if(reset) begin
      T_2197 <= 3'h0;
    end else begin
      if(T_2195) begin
        T_2197 <= T_2202;
      end
    end
    if(reset) begin
      T_2207 <= 1'h0;
    end else begin
      if(T_2216) begin
        T_2207 <= T_2219;
      end else begin
        if(T_2210) begin
          T_2207 <= T_2213;
        end
      end
    end
    if(reset) begin
      T_2712 <= 3'h0;
    end else begin
      if(T_2710) begin
        T_2712 <= T_2717;
      end
    end
    if(reset) begin
      T_2741 <= 3'h0;
    end else begin
      if(T_2739) begin
        T_2741 <= T_2746;
      end
    end
    if(reset) begin
      T_2751 <= 1'h0;
    end else begin
      if(T_2760) begin
        T_2751 <= T_2763;
      end else begin
        if(T_2754) begin
          T_2751 <= T_2757;
        end
      end
    end
    if(reset) begin
      T_2877 <= 3'h0;
    end else begin
      if(T_2875) begin
        T_2877 <= T_2882;
      end
    end
    if(reset) begin
      T_2908 <= 3'h0;
    end else begin
      if(T_2906) begin
        T_2908 <= T_2913;
      end
    end
    if(reset) begin
      T_2918 <= 1'h0;
    end else begin
      if(T_2927) begin
        T_2918 <= T_2930;
      end else begin
        if(T_2921) begin
          T_2918 <= T_2924;
        end
      end
    end
    if(reset) begin
      T_3299 <= 3'h0;
    end else begin
      if(T_3297) begin
        T_3299 <= T_3304;
      end
    end
    if(reset) begin
      T_3314 <= 3'h0;
    end
    if(reset) begin
      T_3324 <= 1'h0;
    end else begin
      if(T_3333) begin
        T_3324 <= T_3336;
      end else begin
        if(T_3327) begin
          T_3324 <= T_3330;
        end
      end
    end
    if(reset) begin
      T_3499 <= 3'h0;
    end else begin
      if(T_3497) begin
        T_3499 <= T_3504;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1652) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at Broadcast.scala:98 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq.should &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1652) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1666) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support Prefetches.\n    at Broadcast.scala:102 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isPrefetch()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1666) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1677) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics.\n    at Broadcast.scala:105 assert(!(state =/= s_idle && pending_ignt && xact_iacq.isAtomic()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1677) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LockingRRArbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [10:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [10:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [2:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [10:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [2:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_addr_beat,
  input   io_in_3_bits_is_builtin_type,
  input  [2:0] io_in_3_bits_a_type,
  input  [10:0] io_in_3_bits_union,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [2:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_addr_beat,
  input   io_in_4_bits_is_builtin_type,
  input  [2:0] io_in_4_bits_a_type,
  input  [10:0] io_in_4_bits_union,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [10:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [2:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_is_builtin_type;
  wire [2:0] GEN_0_bits_a_type;
  wire [10:0] GEN_0_bits_union;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_10;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire [10:0] GEN_15;
  wire [63:0] GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [25:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [2:0] GEN_23;
  wire [10:0] GEN_24;
  wire [63:0] GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [25:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire  GEN_31;
  wire [2:0] GEN_32;
  wire [10:0] GEN_33;
  wire [63:0] GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [25:0] GEN_37;
  wire [2:0] GEN_38;
  wire [2:0] GEN_39;
  wire  GEN_40;
  wire [2:0] GEN_41;
  wire [10:0] GEN_42;
  wire [63:0] GEN_43;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [2:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_is_builtin_type;
  wire [2:0] GEN_1_bits_a_type;
  wire [10:0] GEN_1_bits_union;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [2:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_is_builtin_type;
  wire [2:0] GEN_2_bits_a_type;
  wire [10:0] GEN_2_bits_union;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [2:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_is_builtin_type;
  wire [2:0] GEN_3_bits_a_type;
  wire [10:0] GEN_3_bits_union;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [25:0] GEN_4_bits_addr_block;
  wire [2:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_is_builtin_type;
  wire [2:0] GEN_4_bits_a_type;
  wire [10:0] GEN_4_bits_union;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [25:0] GEN_5_bits_addr_block;
  wire [2:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_is_builtin_type;
  wire [2:0] GEN_5_bits_a_type;
  wire [10:0] GEN_5_bits_union;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [25:0] GEN_6_bits_addr_block;
  wire [2:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_is_builtin_type;
  wire [2:0] GEN_6_bits_a_type;
  wire [10:0] GEN_6_bits_union;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [25:0] GEN_7_bits_addr_block;
  wire [2:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_is_builtin_type;
  wire [2:0] GEN_7_bits_a_type;
  wire [10:0] GEN_7_bits_union;
  wire [63:0] GEN_7_bits_data;
  reg [2:0] T_1114;
  reg [31:0] GEN_0;
  reg [2:0] T_1116;
  reg [31:0] GEN_1;
  wire  T_1118;
  wire [2:0] T_1127_0;
  wire  T_1129;
  wire  T_1130;
  wire  T_1131;
  wire  T_1132;
  wire [3:0] T_1136;
  wire [2:0] T_1137;
  wire [2:0] GEN_296;
  wire [2:0] GEN_297;
  wire [2:0] GEN_298;
  reg [2:0] lastGrant;
  reg [31:0] GEN_2;
  wire [2:0] GEN_299;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  grantMask_4;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  validMask_4;
  wire  T_1146;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire  T_1156;
  wire  T_1158;
  wire  T_1160;
  wire  T_1162;
  wire  T_1164;
  wire  T_1166;
  wire  T_1168;
  wire  T_1170;
  wire  T_1174;
  wire  T_1175;
  wire  T_1176;
  wire  T_1177;
  wire  T_1178;
  wire  T_1179;
  wire  T_1180;
  wire  T_1182;
  wire  T_1183;
  wire  T_1184;
  wire  T_1186;
  wire  T_1187;
  wire  T_1188;
  wire  T_1190;
  wire  T_1191;
  wire  T_1192;
  wire  T_1194;
  wire  T_1195;
  wire  T_1196;
  wire  T_1198;
  wire  T_1199;
  wire  T_1200;
  wire [2:0] GEN_300;
  wire [2:0] GEN_301;
  wire [2:0] GEN_302;
  wire [2:0] GEN_303;
  wire [2:0] GEN_304;
  wire [2:0] GEN_305;
  wire [2:0] GEN_306;
  wire [2:0] GEN_307;
  assign io_in_0_ready = T_1184;
  assign io_in_1_ready = T_1188;
  assign io_in_2_ready = T_1192;
  assign io_in_3_ready = T_1196;
  assign io_in_4_ready = T_1200;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_addr_beat = GEN_3_bits_addr_beat;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_a_type = GEN_5_bits_a_type;
  assign io_out_bits_union = GEN_6_bits_union;
  assign io_out_bits_data = GEN_7_bits_data;
  assign io_chosen = GEN_298;
  assign choice = GEN_307;
  assign GEN_0_ready = GEN_35;
  assign GEN_0_valid = GEN_36;
  assign GEN_0_bits_addr_block = GEN_37;
  assign GEN_0_bits_client_xact_id = GEN_38;
  assign GEN_0_bits_addr_beat = GEN_39;
  assign GEN_0_bits_is_builtin_type = GEN_40;
  assign GEN_0_bits_a_type = GEN_41;
  assign GEN_0_bits_union = GEN_42;
  assign GEN_0_bits_data = GEN_43;
  assign GEN_8 = 3'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = 3'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 3'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 3'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 3'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = 3'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = 3'h1 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_15 = 3'h1 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_16 = 3'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_17 = 3'h2 == io_chosen ? io_in_2_ready : GEN_8;
  assign GEN_18 = 3'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_19 = 3'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_20 = 3'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_21 = 3'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_12;
  assign GEN_22 = 3'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_13;
  assign GEN_23 = 3'h2 == io_chosen ? io_in_2_bits_a_type : GEN_14;
  assign GEN_24 = 3'h2 == io_chosen ? io_in_2_bits_union : GEN_15;
  assign GEN_25 = 3'h2 == io_chosen ? io_in_2_bits_data : GEN_16;
  assign GEN_26 = 3'h3 == io_chosen ? io_in_3_ready : GEN_17;
  assign GEN_27 = 3'h3 == io_chosen ? io_in_3_valid : GEN_18;
  assign GEN_28 = 3'h3 == io_chosen ? io_in_3_bits_addr_block : GEN_19;
  assign GEN_29 = 3'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_20;
  assign GEN_30 = 3'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_21;
  assign GEN_31 = 3'h3 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_22;
  assign GEN_32 = 3'h3 == io_chosen ? io_in_3_bits_a_type : GEN_23;
  assign GEN_33 = 3'h3 == io_chosen ? io_in_3_bits_union : GEN_24;
  assign GEN_34 = 3'h3 == io_chosen ? io_in_3_bits_data : GEN_25;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_ready : GEN_26;
  assign GEN_36 = 3'h4 == io_chosen ? io_in_4_valid : GEN_27;
  assign GEN_37 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_28;
  assign GEN_38 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_29;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_30;
  assign GEN_40 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_31;
  assign GEN_41 = 3'h4 == io_chosen ? io_in_4_bits_a_type : GEN_32;
  assign GEN_42 = 3'h4 == io_chosen ? io_in_4_bits_union : GEN_33;
  assign GEN_43 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_34;
  assign GEN_1_ready = GEN_35;
  assign GEN_1_valid = GEN_36;
  assign GEN_1_bits_addr_block = GEN_37;
  assign GEN_1_bits_client_xact_id = GEN_38;
  assign GEN_1_bits_addr_beat = GEN_39;
  assign GEN_1_bits_is_builtin_type = GEN_40;
  assign GEN_1_bits_a_type = GEN_41;
  assign GEN_1_bits_union = GEN_42;
  assign GEN_1_bits_data = GEN_43;
  assign GEN_2_ready = GEN_35;
  assign GEN_2_valid = GEN_36;
  assign GEN_2_bits_addr_block = GEN_37;
  assign GEN_2_bits_client_xact_id = GEN_38;
  assign GEN_2_bits_addr_beat = GEN_39;
  assign GEN_2_bits_is_builtin_type = GEN_40;
  assign GEN_2_bits_a_type = GEN_41;
  assign GEN_2_bits_union = GEN_42;
  assign GEN_2_bits_data = GEN_43;
  assign GEN_3_ready = GEN_35;
  assign GEN_3_valid = GEN_36;
  assign GEN_3_bits_addr_block = GEN_37;
  assign GEN_3_bits_client_xact_id = GEN_38;
  assign GEN_3_bits_addr_beat = GEN_39;
  assign GEN_3_bits_is_builtin_type = GEN_40;
  assign GEN_3_bits_a_type = GEN_41;
  assign GEN_3_bits_union = GEN_42;
  assign GEN_3_bits_data = GEN_43;
  assign GEN_4_ready = GEN_35;
  assign GEN_4_valid = GEN_36;
  assign GEN_4_bits_addr_block = GEN_37;
  assign GEN_4_bits_client_xact_id = GEN_38;
  assign GEN_4_bits_addr_beat = GEN_39;
  assign GEN_4_bits_is_builtin_type = GEN_40;
  assign GEN_4_bits_a_type = GEN_41;
  assign GEN_4_bits_union = GEN_42;
  assign GEN_4_bits_data = GEN_43;
  assign GEN_5_ready = GEN_35;
  assign GEN_5_valid = GEN_36;
  assign GEN_5_bits_addr_block = GEN_37;
  assign GEN_5_bits_client_xact_id = GEN_38;
  assign GEN_5_bits_addr_beat = GEN_39;
  assign GEN_5_bits_is_builtin_type = GEN_40;
  assign GEN_5_bits_a_type = GEN_41;
  assign GEN_5_bits_union = GEN_42;
  assign GEN_5_bits_data = GEN_43;
  assign GEN_6_ready = GEN_35;
  assign GEN_6_valid = GEN_36;
  assign GEN_6_bits_addr_block = GEN_37;
  assign GEN_6_bits_client_xact_id = GEN_38;
  assign GEN_6_bits_addr_beat = GEN_39;
  assign GEN_6_bits_is_builtin_type = GEN_40;
  assign GEN_6_bits_a_type = GEN_41;
  assign GEN_6_bits_union = GEN_42;
  assign GEN_6_bits_data = GEN_43;
  assign GEN_7_ready = GEN_35;
  assign GEN_7_valid = GEN_36;
  assign GEN_7_bits_addr_block = GEN_37;
  assign GEN_7_bits_client_xact_id = GEN_38;
  assign GEN_7_bits_addr_beat = GEN_39;
  assign GEN_7_bits_is_builtin_type = GEN_40;
  assign GEN_7_bits_a_type = GEN_41;
  assign GEN_7_bits_union = GEN_42;
  assign GEN_7_bits_data = GEN_43;
  assign T_1118 = T_1114 != 3'h0;
  assign T_1127_0 = 3'h3;
  assign T_1129 = io_out_bits_a_type == T_1127_0;
  assign T_1130 = io_out_bits_is_builtin_type & T_1129;
  assign T_1131 = io_out_ready & io_out_valid;
  assign T_1132 = T_1131 & T_1130;
  assign T_1136 = T_1114 + 3'h1;
  assign T_1137 = T_1136[2:0];
  assign GEN_296 = T_1132 ? io_chosen : T_1116;
  assign GEN_297 = T_1132 ? T_1137 : T_1114;
  assign GEN_298 = T_1118 ? T_1116 : choice;
  assign GEN_299 = T_1131 ? io_chosen : lastGrant;
  assign grantMask_1 = 3'h1 > lastGrant;
  assign grantMask_2 = 3'h2 > lastGrant;
  assign grantMask_3 = 3'h3 > lastGrant;
  assign grantMask_4 = 3'h4 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign validMask_4 = io_in_4_valid & grantMask_4;
  assign T_1146 = validMask_1 | validMask_2;
  assign T_1147 = T_1146 | validMask_3;
  assign T_1148 = T_1147 | validMask_4;
  assign T_1149 = T_1148 | io_in_0_valid;
  assign T_1150 = T_1149 | io_in_1_valid;
  assign T_1151 = T_1150 | io_in_2_valid;
  assign T_1152 = T_1151 | io_in_3_valid;
  assign T_1156 = validMask_1 == 1'h0;
  assign T_1158 = T_1146 == 1'h0;
  assign T_1160 = T_1147 == 1'h0;
  assign T_1162 = T_1148 == 1'h0;
  assign T_1164 = T_1149 == 1'h0;
  assign T_1166 = T_1150 == 1'h0;
  assign T_1168 = T_1151 == 1'h0;
  assign T_1170 = T_1152 == 1'h0;
  assign T_1174 = grantMask_1 | T_1164;
  assign T_1175 = T_1156 & grantMask_2;
  assign T_1176 = T_1175 | T_1166;
  assign T_1177 = T_1158 & grantMask_3;
  assign T_1178 = T_1177 | T_1168;
  assign T_1179 = T_1160 & grantMask_4;
  assign T_1180 = T_1179 | T_1170;
  assign T_1182 = T_1116 == 3'h0;
  assign T_1183 = T_1118 ? T_1182 : T_1162;
  assign T_1184 = T_1183 & io_out_ready;
  assign T_1186 = T_1116 == 3'h1;
  assign T_1187 = T_1118 ? T_1186 : T_1174;
  assign T_1188 = T_1187 & io_out_ready;
  assign T_1190 = T_1116 == 3'h2;
  assign T_1191 = T_1118 ? T_1190 : T_1176;
  assign T_1192 = T_1191 & io_out_ready;
  assign T_1194 = T_1116 == 3'h3;
  assign T_1195 = T_1118 ? T_1194 : T_1178;
  assign T_1196 = T_1195 & io_out_ready;
  assign T_1198 = T_1116 == 3'h4;
  assign T_1199 = T_1118 ? T_1198 : T_1180;
  assign T_1200 = T_1199 & io_out_ready;
  assign GEN_300 = io_in_3_valid ? 3'h3 : 3'h4;
  assign GEN_301 = io_in_2_valid ? 3'h2 : GEN_300;
  assign GEN_302 = io_in_1_valid ? 3'h1 : GEN_301;
  assign GEN_303 = io_in_0_valid ? 3'h0 : GEN_302;
  assign GEN_304 = validMask_4 ? 3'h4 : GEN_303;
  assign GEN_305 = validMask_3 ? 3'h3 : GEN_304;
  assign GEN_306 = validMask_2 ? 3'h2 : GEN_305;
  assign GEN_307 = validMask_1 ? 3'h1 : GEN_306;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1114 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1116 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1114 <= 3'h0;
    end else begin
      if(T_1132) begin
        T_1114 <= T_1137;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1132) begin
        T_1116 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1131) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [25:0] io_in_2_bits_addr_block,
  input  [2:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_voluntary,
  input  [2:0] io_in_2_bits_r_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [25:0] io_in_3_bits_addr_block,
  input  [2:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_voluntary,
  input  [2:0] io_in_3_bits_r_type,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [25:0] io_in_4_bits_addr_block,
  input  [2:0] io_in_4_bits_client_xact_id,
  input   io_in_4_bits_voluntary,
  input  [2:0] io_in_4_bits_r_type,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [25:0] GEN_0_bits_addr_block;
  wire [2:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_voluntary;
  wire [2:0] GEN_0_bits_r_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [25:0] GEN_10;
  wire [2:0] GEN_11;
  wire  GEN_12;
  wire [2:0] GEN_13;
  wire [63:0] GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [25:0] GEN_18;
  wire [2:0] GEN_19;
  wire  GEN_20;
  wire [2:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_25;
  wire [25:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [2:0] GEN_29;
  wire [63:0] GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire [2:0] GEN_33;
  wire [25:0] GEN_34;
  wire [2:0] GEN_35;
  wire  GEN_36;
  wire [2:0] GEN_37;
  wire [63:0] GEN_38;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [25:0] GEN_1_bits_addr_block;
  wire [2:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_voluntary;
  wire [2:0] GEN_1_bits_r_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [25:0] GEN_2_bits_addr_block;
  wire [2:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_voluntary;
  wire [2:0] GEN_2_bits_r_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [25:0] GEN_3_bits_addr_block;
  wire [2:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_voluntary;
  wire [2:0] GEN_3_bits_r_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [25:0] GEN_4_bits_addr_block;
  wire [2:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_voluntary;
  wire [2:0] GEN_4_bits_r_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [25:0] GEN_5_bits_addr_block;
  wire [2:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_voluntary;
  wire [2:0] GEN_5_bits_r_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [25:0] GEN_6_bits_addr_block;
  wire [2:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_voluntary;
  wire [2:0] GEN_6_bits_r_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_1076;
  reg [31:0] GEN_0;
  reg [2:0] T_1078;
  reg [31:0] GEN_1;
  wire  T_1080;
  wire  T_1082;
  wire  T_1083;
  wire  T_1084;
  wire  T_1085;
  wire  T_1086;
  wire  T_1088;
  wire  T_1089;
  wire [3:0] T_1093;
  wire [2:0] T_1094;
  wire [2:0] GEN_231;
  wire [2:0] GEN_232;
  wire [2:0] GEN_233;
  reg [2:0] lastGrant;
  reg [31:0] GEN_2;
  wire [2:0] GEN_234;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  grantMask_4;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  validMask_4;
  wire  T_1103;
  wire  T_1104;
  wire  T_1105;
  wire  T_1106;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1113;
  wire  T_1115;
  wire  T_1117;
  wire  T_1119;
  wire  T_1121;
  wire  T_1123;
  wire  T_1125;
  wire  T_1127;
  wire  T_1131;
  wire  T_1132;
  wire  T_1133;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire  T_1137;
  wire  T_1139;
  wire  T_1140;
  wire  T_1141;
  wire  T_1143;
  wire  T_1144;
  wire  T_1145;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire [2:0] GEN_235;
  wire [2:0] GEN_236;
  wire [2:0] GEN_237;
  wire [2:0] GEN_238;
  wire [2:0] GEN_239;
  wire [2:0] GEN_240;
  wire [2:0] GEN_241;
  wire [2:0] GEN_242;
  assign io_in_0_ready = T_1141;
  assign io_in_1_ready = T_1145;
  assign io_in_2_ready = T_1149;
  assign io_in_3_ready = T_1153;
  assign io_in_4_ready = T_1157;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_addr_block = GEN_2_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_3_bits_client_xact_id;
  assign io_out_bits_voluntary = GEN_4_bits_voluntary;
  assign io_out_bits_r_type = GEN_5_bits_r_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_233;
  assign choice = GEN_242;
  assign GEN_0_ready = GEN_31;
  assign GEN_0_valid = GEN_32;
  assign GEN_0_bits_addr_beat = GEN_33;
  assign GEN_0_bits_addr_block = GEN_34;
  assign GEN_0_bits_client_xact_id = GEN_35;
  assign GEN_0_bits_voluntary = GEN_36;
  assign GEN_0_bits_r_type = GEN_37;
  assign GEN_0_bits_data = GEN_38;
  assign GEN_7 = 3'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = 3'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 3'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_10 = 3'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 3'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 3'h1 == io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_13 = 3'h1 == io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_14 = 3'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_15 = 3'h2 == io_chosen ? io_in_2_ready : GEN_7;
  assign GEN_16 = 3'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_17 = 3'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_9;
  assign GEN_18 = 3'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_19 = 3'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_20 = 3'h2 == io_chosen ? io_in_2_bits_voluntary : GEN_12;
  assign GEN_21 = 3'h2 == io_chosen ? io_in_2_bits_r_type : GEN_13;
  assign GEN_22 = 3'h2 == io_chosen ? io_in_2_bits_data : GEN_14;
  assign GEN_23 = 3'h3 == io_chosen ? io_in_3_ready : GEN_15;
  assign GEN_24 = 3'h3 == io_chosen ? io_in_3_valid : GEN_16;
  assign GEN_25 = 3'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_17;
  assign GEN_26 = 3'h3 == io_chosen ? io_in_3_bits_addr_block : GEN_18;
  assign GEN_27 = 3'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_19;
  assign GEN_28 = 3'h3 == io_chosen ? io_in_3_bits_voluntary : GEN_20;
  assign GEN_29 = 3'h3 == io_chosen ? io_in_3_bits_r_type : GEN_21;
  assign GEN_30 = 3'h3 == io_chosen ? io_in_3_bits_data : GEN_22;
  assign GEN_31 = 3'h4 == io_chosen ? io_in_4_ready : GEN_23;
  assign GEN_32 = 3'h4 == io_chosen ? io_in_4_valid : GEN_24;
  assign GEN_33 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_25;
  assign GEN_34 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_26;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_27;
  assign GEN_36 = 3'h4 == io_chosen ? io_in_4_bits_voluntary : GEN_28;
  assign GEN_37 = 3'h4 == io_chosen ? io_in_4_bits_r_type : GEN_29;
  assign GEN_38 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_30;
  assign GEN_1_ready = GEN_31;
  assign GEN_1_valid = GEN_32;
  assign GEN_1_bits_addr_beat = GEN_33;
  assign GEN_1_bits_addr_block = GEN_34;
  assign GEN_1_bits_client_xact_id = GEN_35;
  assign GEN_1_bits_voluntary = GEN_36;
  assign GEN_1_bits_r_type = GEN_37;
  assign GEN_1_bits_data = GEN_38;
  assign GEN_2_ready = GEN_31;
  assign GEN_2_valid = GEN_32;
  assign GEN_2_bits_addr_beat = GEN_33;
  assign GEN_2_bits_addr_block = GEN_34;
  assign GEN_2_bits_client_xact_id = GEN_35;
  assign GEN_2_bits_voluntary = GEN_36;
  assign GEN_2_bits_r_type = GEN_37;
  assign GEN_2_bits_data = GEN_38;
  assign GEN_3_ready = GEN_31;
  assign GEN_3_valid = GEN_32;
  assign GEN_3_bits_addr_beat = GEN_33;
  assign GEN_3_bits_addr_block = GEN_34;
  assign GEN_3_bits_client_xact_id = GEN_35;
  assign GEN_3_bits_voluntary = GEN_36;
  assign GEN_3_bits_r_type = GEN_37;
  assign GEN_3_bits_data = GEN_38;
  assign GEN_4_ready = GEN_31;
  assign GEN_4_valid = GEN_32;
  assign GEN_4_bits_addr_beat = GEN_33;
  assign GEN_4_bits_addr_block = GEN_34;
  assign GEN_4_bits_client_xact_id = GEN_35;
  assign GEN_4_bits_voluntary = GEN_36;
  assign GEN_4_bits_r_type = GEN_37;
  assign GEN_4_bits_data = GEN_38;
  assign GEN_5_ready = GEN_31;
  assign GEN_5_valid = GEN_32;
  assign GEN_5_bits_addr_beat = GEN_33;
  assign GEN_5_bits_addr_block = GEN_34;
  assign GEN_5_bits_client_xact_id = GEN_35;
  assign GEN_5_bits_voluntary = GEN_36;
  assign GEN_5_bits_r_type = GEN_37;
  assign GEN_5_bits_data = GEN_38;
  assign GEN_6_ready = GEN_31;
  assign GEN_6_valid = GEN_32;
  assign GEN_6_bits_addr_beat = GEN_33;
  assign GEN_6_bits_addr_block = GEN_34;
  assign GEN_6_bits_client_xact_id = GEN_35;
  assign GEN_6_bits_voluntary = GEN_36;
  assign GEN_6_bits_r_type = GEN_37;
  assign GEN_6_bits_data = GEN_38;
  assign T_1080 = T_1076 != 3'h0;
  assign T_1082 = io_out_bits_r_type == 3'h0;
  assign T_1083 = io_out_bits_r_type == 3'h1;
  assign T_1084 = io_out_bits_r_type == 3'h2;
  assign T_1085 = T_1082 | T_1083;
  assign T_1086 = T_1085 | T_1084;
  assign T_1088 = io_out_ready & io_out_valid;
  assign T_1089 = T_1088 & T_1086;
  assign T_1093 = T_1076 + 3'h1;
  assign T_1094 = T_1093[2:0];
  assign GEN_231 = T_1089 ? io_chosen : T_1078;
  assign GEN_232 = T_1089 ? T_1094 : T_1076;
  assign GEN_233 = T_1080 ? T_1078 : choice;
  assign GEN_234 = T_1088 ? io_chosen : lastGrant;
  assign grantMask_1 = 3'h1 > lastGrant;
  assign grantMask_2 = 3'h2 > lastGrant;
  assign grantMask_3 = 3'h3 > lastGrant;
  assign grantMask_4 = 3'h4 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign validMask_4 = io_in_4_valid & grantMask_4;
  assign T_1103 = validMask_1 | validMask_2;
  assign T_1104 = T_1103 | validMask_3;
  assign T_1105 = T_1104 | validMask_4;
  assign T_1106 = T_1105 | io_in_0_valid;
  assign T_1107 = T_1106 | io_in_1_valid;
  assign T_1108 = T_1107 | io_in_2_valid;
  assign T_1109 = T_1108 | io_in_3_valid;
  assign T_1113 = validMask_1 == 1'h0;
  assign T_1115 = T_1103 == 1'h0;
  assign T_1117 = T_1104 == 1'h0;
  assign T_1119 = T_1105 == 1'h0;
  assign T_1121 = T_1106 == 1'h0;
  assign T_1123 = T_1107 == 1'h0;
  assign T_1125 = T_1108 == 1'h0;
  assign T_1127 = T_1109 == 1'h0;
  assign T_1131 = grantMask_1 | T_1121;
  assign T_1132 = T_1113 & grantMask_2;
  assign T_1133 = T_1132 | T_1123;
  assign T_1134 = T_1115 & grantMask_3;
  assign T_1135 = T_1134 | T_1125;
  assign T_1136 = T_1117 & grantMask_4;
  assign T_1137 = T_1136 | T_1127;
  assign T_1139 = T_1078 == 3'h0;
  assign T_1140 = T_1080 ? T_1139 : T_1119;
  assign T_1141 = T_1140 & io_out_ready;
  assign T_1143 = T_1078 == 3'h1;
  assign T_1144 = T_1080 ? T_1143 : T_1131;
  assign T_1145 = T_1144 & io_out_ready;
  assign T_1147 = T_1078 == 3'h2;
  assign T_1148 = T_1080 ? T_1147 : T_1133;
  assign T_1149 = T_1148 & io_out_ready;
  assign T_1151 = T_1078 == 3'h3;
  assign T_1152 = T_1080 ? T_1151 : T_1135;
  assign T_1153 = T_1152 & io_out_ready;
  assign T_1155 = T_1078 == 3'h4;
  assign T_1156 = T_1080 ? T_1155 : T_1137;
  assign T_1157 = T_1156 & io_out_ready;
  assign GEN_235 = io_in_3_valid ? 3'h3 : 3'h4;
  assign GEN_236 = io_in_2_valid ? 3'h2 : GEN_235;
  assign GEN_237 = io_in_1_valid ? 3'h1 : GEN_236;
  assign GEN_238 = io_in_0_valid ? 3'h0 : GEN_237;
  assign GEN_239 = validMask_4 ? 3'h4 : GEN_238;
  assign GEN_240 = validMask_3 ? 3'h3 : GEN_239;
  assign GEN_241 = validMask_2 ? 3'h2 : GEN_240;
  assign GEN_242 = validMask_1 ? 3'h1 : GEN_241;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_1076 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1078 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1076 <= 3'h0;
    end else begin
      if(T_1089) begin
        T_1076 <= T_1094;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1089) begin
        T_1078 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1088) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_probe_ready,
  output  io_in_0_probe_valid,
  output [25:0] io_in_0_probe_bits_addr_block,
  output [1:0] io_in_0_probe_bits_p_type,
  output  io_in_0_release_ready,
  input   io_in_0_release_valid,
  input  [2:0] io_in_0_release_bits_addr_beat,
  input  [25:0] io_in_0_release_bits_addr_block,
  input  [2:0] io_in_0_release_bits_client_xact_id,
  input   io_in_0_release_bits_voluntary,
  input  [2:0] io_in_0_release_bits_r_type,
  input  [63:0] io_in_0_release_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  output  io_in_0_grant_bits_manager_id,
  output  io_in_0_finish_ready,
  input   io_in_0_finish_valid,
  input   io_in_0_finish_bits_manager_xact_id,
  input   io_in_0_finish_bits_manager_id,
  output  io_in_1_acquire_ready,
  input   io_in_1_acquire_valid,
  input  [25:0] io_in_1_acquire_bits_addr_block,
  input  [2:0] io_in_1_acquire_bits_client_xact_id,
  input  [2:0] io_in_1_acquire_bits_addr_beat,
  input   io_in_1_acquire_bits_is_builtin_type,
  input  [2:0] io_in_1_acquire_bits_a_type,
  input  [10:0] io_in_1_acquire_bits_union,
  input  [63:0] io_in_1_acquire_bits_data,
  input   io_in_1_probe_ready,
  output  io_in_1_probe_valid,
  output [25:0] io_in_1_probe_bits_addr_block,
  output [1:0] io_in_1_probe_bits_p_type,
  output  io_in_1_release_ready,
  input   io_in_1_release_valid,
  input  [2:0] io_in_1_release_bits_addr_beat,
  input  [25:0] io_in_1_release_bits_addr_block,
  input  [2:0] io_in_1_release_bits_client_xact_id,
  input   io_in_1_release_bits_voluntary,
  input  [2:0] io_in_1_release_bits_r_type,
  input  [63:0] io_in_1_release_bits_data,
  input   io_in_1_grant_ready,
  output  io_in_1_grant_valid,
  output [2:0] io_in_1_grant_bits_addr_beat,
  output [2:0] io_in_1_grant_bits_client_xact_id,
  output  io_in_1_grant_bits_manager_xact_id,
  output  io_in_1_grant_bits_is_builtin_type,
  output [3:0] io_in_1_grant_bits_g_type,
  output [63:0] io_in_1_grant_bits_data,
  output  io_in_1_grant_bits_manager_id,
  output  io_in_1_finish_ready,
  input   io_in_1_finish_valid,
  input   io_in_1_finish_bits_manager_xact_id,
  input   io_in_1_finish_bits_manager_id,
  output  io_in_2_acquire_ready,
  input   io_in_2_acquire_valid,
  input  [25:0] io_in_2_acquire_bits_addr_block,
  input  [2:0] io_in_2_acquire_bits_client_xact_id,
  input  [2:0] io_in_2_acquire_bits_addr_beat,
  input   io_in_2_acquire_bits_is_builtin_type,
  input  [2:0] io_in_2_acquire_bits_a_type,
  input  [10:0] io_in_2_acquire_bits_union,
  input  [63:0] io_in_2_acquire_bits_data,
  input   io_in_2_probe_ready,
  output  io_in_2_probe_valid,
  output [25:0] io_in_2_probe_bits_addr_block,
  output [1:0] io_in_2_probe_bits_p_type,
  output  io_in_2_release_ready,
  input   io_in_2_release_valid,
  input  [2:0] io_in_2_release_bits_addr_beat,
  input  [25:0] io_in_2_release_bits_addr_block,
  input  [2:0] io_in_2_release_bits_client_xact_id,
  input   io_in_2_release_bits_voluntary,
  input  [2:0] io_in_2_release_bits_r_type,
  input  [63:0] io_in_2_release_bits_data,
  input   io_in_2_grant_ready,
  output  io_in_2_grant_valid,
  output [2:0] io_in_2_grant_bits_addr_beat,
  output [2:0] io_in_2_grant_bits_client_xact_id,
  output  io_in_2_grant_bits_manager_xact_id,
  output  io_in_2_grant_bits_is_builtin_type,
  output [3:0] io_in_2_grant_bits_g_type,
  output [63:0] io_in_2_grant_bits_data,
  output  io_in_2_grant_bits_manager_id,
  output  io_in_2_finish_ready,
  input   io_in_2_finish_valid,
  input   io_in_2_finish_bits_manager_xact_id,
  input   io_in_2_finish_bits_manager_id,
  output  io_in_3_acquire_ready,
  input   io_in_3_acquire_valid,
  input  [25:0] io_in_3_acquire_bits_addr_block,
  input  [2:0] io_in_3_acquire_bits_client_xact_id,
  input  [2:0] io_in_3_acquire_bits_addr_beat,
  input   io_in_3_acquire_bits_is_builtin_type,
  input  [2:0] io_in_3_acquire_bits_a_type,
  input  [10:0] io_in_3_acquire_bits_union,
  input  [63:0] io_in_3_acquire_bits_data,
  input   io_in_3_probe_ready,
  output  io_in_3_probe_valid,
  output [25:0] io_in_3_probe_bits_addr_block,
  output [1:0] io_in_3_probe_bits_p_type,
  output  io_in_3_release_ready,
  input   io_in_3_release_valid,
  input  [2:0] io_in_3_release_bits_addr_beat,
  input  [25:0] io_in_3_release_bits_addr_block,
  input  [2:0] io_in_3_release_bits_client_xact_id,
  input   io_in_3_release_bits_voluntary,
  input  [2:0] io_in_3_release_bits_r_type,
  input  [63:0] io_in_3_release_bits_data,
  input   io_in_3_grant_ready,
  output  io_in_3_grant_valid,
  output [2:0] io_in_3_grant_bits_addr_beat,
  output [2:0] io_in_3_grant_bits_client_xact_id,
  output  io_in_3_grant_bits_manager_xact_id,
  output  io_in_3_grant_bits_is_builtin_type,
  output [3:0] io_in_3_grant_bits_g_type,
  output [63:0] io_in_3_grant_bits_data,
  output  io_in_3_grant_bits_manager_id,
  output  io_in_3_finish_ready,
  input   io_in_3_finish_valid,
  input   io_in_3_finish_bits_manager_xact_id,
  input   io_in_3_finish_bits_manager_id,
  output  io_in_4_acquire_ready,
  input   io_in_4_acquire_valid,
  input  [25:0] io_in_4_acquire_bits_addr_block,
  input  [2:0] io_in_4_acquire_bits_client_xact_id,
  input  [2:0] io_in_4_acquire_bits_addr_beat,
  input   io_in_4_acquire_bits_is_builtin_type,
  input  [2:0] io_in_4_acquire_bits_a_type,
  input  [10:0] io_in_4_acquire_bits_union,
  input  [63:0] io_in_4_acquire_bits_data,
  input   io_in_4_probe_ready,
  output  io_in_4_probe_valid,
  output [25:0] io_in_4_probe_bits_addr_block,
  output [1:0] io_in_4_probe_bits_p_type,
  output  io_in_4_release_ready,
  input   io_in_4_release_valid,
  input  [2:0] io_in_4_release_bits_addr_beat,
  input  [25:0] io_in_4_release_bits_addr_block,
  input  [2:0] io_in_4_release_bits_client_xact_id,
  input   io_in_4_release_bits_voluntary,
  input  [2:0] io_in_4_release_bits_r_type,
  input  [63:0] io_in_4_release_bits_data,
  input   io_in_4_grant_ready,
  output  io_in_4_grant_valid,
  output [2:0] io_in_4_grant_bits_addr_beat,
  output [2:0] io_in_4_grant_bits_client_xact_id,
  output  io_in_4_grant_bits_manager_xact_id,
  output  io_in_4_grant_bits_is_builtin_type,
  output [3:0] io_in_4_grant_bits_g_type,
  output [63:0] io_in_4_grant_bits_data,
  output  io_in_4_grant_bits_manager_id,
  output  io_in_4_finish_ready,
  input   io_in_4_finish_valid,
  input   io_in_4_finish_bits_manager_xact_id,
  input   io_in_4_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_probe_ready,
  input   io_out_probe_valid,
  input  [25:0] io_out_probe_bits_addr_block,
  input  [1:0] io_out_probe_bits_p_type,
  input   io_out_release_ready,
  output  io_out_release_valid,
  output [2:0] io_out_release_bits_addr_beat,
  output [25:0] io_out_release_bits_addr_block,
  output [2:0] io_out_release_bits_client_xact_id,
  output  io_out_release_bits_voluntary,
  output [2:0] io_out_release_bits_r_type,
  output [63:0] io_out_release_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data,
  input   io_out_grant_bits_manager_id,
  input   io_out_finish_ready,
  output  io_out_finish_valid,
  output  io_out_finish_bits_manager_xact_id,
  output  io_out_finish_bits_manager_id
);
  wire  LockingRRArbiter_5_1_clk;
  wire  LockingRRArbiter_5_1_reset;
  wire  LockingRRArbiter_5_1_io_in_0_ready;
  wire  LockingRRArbiter_5_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_0_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_0_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_0_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_0_bits_data;
  wire  LockingRRArbiter_5_1_io_in_1_ready;
  wire  LockingRRArbiter_5_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_1_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_1_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_1_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_1_bits_data;
  wire  LockingRRArbiter_5_1_io_in_2_ready;
  wire  LockingRRArbiter_5_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_2_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_2_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_2_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_2_bits_data;
  wire  LockingRRArbiter_5_1_io_in_3_ready;
  wire  LockingRRArbiter_5_1_io_in_3_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_3_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_3_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_3_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_3_bits_data;
  wire  LockingRRArbiter_5_1_io_in_4_ready;
  wire  LockingRRArbiter_5_1_io_in_4_valid;
  wire [25:0] LockingRRArbiter_5_1_io_in_4_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_in_4_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_in_4_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_in_4_bits_data;
  wire  LockingRRArbiter_5_1_io_out_ready;
  wire  LockingRRArbiter_5_1_io_out_valid;
  wire [25:0] LockingRRArbiter_5_1_io_out_bits_addr_block;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_addr_beat;
  wire  LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_5_1_io_out_bits_a_type;
  wire [10:0] LockingRRArbiter_5_1_io_out_bits_union;
  wire [63:0] LockingRRArbiter_5_1_io_out_bits_data;
  wire [2:0] LockingRRArbiter_5_1_io_chosen;
  wire [5:0] T_9040;
  wire [5:0] T_9042;
  wire [5:0] T_9044;
  wire [5:0] T_9046;
  wire [5:0] T_9048;
  wire  LockingRRArbiter_6_1_clk;
  wire  LockingRRArbiter_6_1_reset;
  wire  LockingRRArbiter_6_1_io_in_0_ready;
  wire  LockingRRArbiter_6_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_0_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_0_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_0_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_0_bits_data;
  wire  LockingRRArbiter_6_1_io_in_1_ready;
  wire  LockingRRArbiter_6_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_1_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_1_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_1_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_1_bits_data;
  wire  LockingRRArbiter_6_1_io_in_2_ready;
  wire  LockingRRArbiter_6_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_2_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_2_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_2_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_2_bits_data;
  wire  LockingRRArbiter_6_1_io_in_3_ready;
  wire  LockingRRArbiter_6_1_io_in_3_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_3_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_3_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_3_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_3_bits_data;
  wire  LockingRRArbiter_6_1_io_in_4_ready;
  wire  LockingRRArbiter_6_1_io_in_4_valid;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_in_4_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_in_4_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_in_4_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_in_4_bits_data;
  wire  LockingRRArbiter_6_1_io_out_ready;
  wire  LockingRRArbiter_6_1_io_out_valid;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_addr_beat;
  wire [25:0] LockingRRArbiter_6_1_io_out_bits_addr_block;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  wire  LockingRRArbiter_6_1_io_out_bits_voluntary;
  wire [2:0] LockingRRArbiter_6_1_io_out_bits_r_type;
  wire [63:0] LockingRRArbiter_6_1_io_out_bits_data;
  wire [2:0] LockingRRArbiter_6_1_io_chosen;
  wire [5:0] T_9050;
  wire [5:0] T_9052;
  wire [5:0] T_9054;
  wire [5:0] T_9056;
  wire [5:0] T_9058;
  wire  T_9059;
  wire  T_9060;
  wire  T_9061;
  wire  T_9062;
  wire  T_9067;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_9072;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_9077;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_9082;
  wire  GEN_6;
  wire  GEN_7;
  wire  T_9087;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  reg [31:0] GEN_18;
  wire  GEN_11;
  reg [31:0] GEN_19;
  wire  GEN_12;
  reg [31:0] GEN_20;
  wire  GEN_13;
  reg [31:0] GEN_21;
  wire  GEN_14;
  reg [31:0] GEN_22;
  wire  GEN_15;
  reg [31:0] GEN_23;
  wire  GEN_16;
  reg [31:0] GEN_24;
  wire  GEN_17;
  reg [31:0] GEN_25;
  LockingRRArbiter_5 LockingRRArbiter_5_1 (
    .clk(LockingRRArbiter_5_1_clk),
    .reset(LockingRRArbiter_5_1_reset),
    .io_in_0_ready(LockingRRArbiter_5_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_5_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_5_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_5_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(LockingRRArbiter_5_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(LockingRRArbiter_5_1_io_in_0_bits_a_type),
    .io_in_0_bits_union(LockingRRArbiter_5_1_io_in_0_bits_union),
    .io_in_0_bits_data(LockingRRArbiter_5_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_5_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_5_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_5_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_5_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(LockingRRArbiter_5_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(LockingRRArbiter_5_1_io_in_1_bits_a_type),
    .io_in_1_bits_union(LockingRRArbiter_5_1_io_in_1_bits_union),
    .io_in_1_bits_data(LockingRRArbiter_5_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_5_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_5_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_5_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_5_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(LockingRRArbiter_5_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(LockingRRArbiter_5_1_io_in_2_bits_a_type),
    .io_in_2_bits_union(LockingRRArbiter_5_1_io_in_2_bits_union),
    .io_in_2_bits_data(LockingRRArbiter_5_1_io_in_2_bits_data),
    .io_in_3_ready(LockingRRArbiter_5_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_5_1_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_5_1_io_in_3_bits_addr_block),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_5_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_addr_beat(LockingRRArbiter_5_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_a_type(LockingRRArbiter_5_1_io_in_3_bits_a_type),
    .io_in_3_bits_union(LockingRRArbiter_5_1_io_in_3_bits_union),
    .io_in_3_bits_data(LockingRRArbiter_5_1_io_in_3_bits_data),
    .io_in_4_ready(LockingRRArbiter_5_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_5_1_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_5_1_io_in_4_bits_addr_block),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_5_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_addr_beat(LockingRRArbiter_5_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_a_type(LockingRRArbiter_5_1_io_in_4_bits_a_type),
    .io_in_4_bits_union(LockingRRArbiter_5_1_io_in_4_bits_union),
    .io_in_4_bits_data(LockingRRArbiter_5_1_io_in_4_bits_data),
    .io_out_ready(LockingRRArbiter_5_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_5_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_5_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_5_1_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(LockingRRArbiter_5_1_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(LockingRRArbiter_5_1_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(LockingRRArbiter_5_1_io_out_bits_a_type),
    .io_out_bits_union(LockingRRArbiter_5_1_io_out_bits_union),
    .io_out_bits_data(LockingRRArbiter_5_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_5_1_io_chosen)
  );
  LockingRRArbiter_6 LockingRRArbiter_6_1 (
    .clk(LockingRRArbiter_6_1_clk),
    .reset(LockingRRArbiter_6_1_reset),
    .io_in_0_ready(LockingRRArbiter_6_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_6_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_6_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(LockingRRArbiter_6_1_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_6_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(LockingRRArbiter_6_1_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(LockingRRArbiter_6_1_io_in_0_bits_r_type),
    .io_in_0_bits_data(LockingRRArbiter_6_1_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_6_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_6_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_6_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(LockingRRArbiter_6_1_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_6_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(LockingRRArbiter_6_1_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(LockingRRArbiter_6_1_io_in_1_bits_r_type),
    .io_in_1_bits_data(LockingRRArbiter_6_1_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_6_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_6_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_6_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_addr_block(LockingRRArbiter_6_1_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_6_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_voluntary(LockingRRArbiter_6_1_io_in_2_bits_voluntary),
    .io_in_2_bits_r_type(LockingRRArbiter_6_1_io_in_2_bits_r_type),
    .io_in_2_bits_data(LockingRRArbiter_6_1_io_in_2_bits_data),
    .io_in_3_ready(LockingRRArbiter_6_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_6_1_io_in_3_valid),
    .io_in_3_bits_addr_beat(LockingRRArbiter_6_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_addr_block(LockingRRArbiter_6_1_io_in_3_bits_addr_block),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_6_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_voluntary(LockingRRArbiter_6_1_io_in_3_bits_voluntary),
    .io_in_3_bits_r_type(LockingRRArbiter_6_1_io_in_3_bits_r_type),
    .io_in_3_bits_data(LockingRRArbiter_6_1_io_in_3_bits_data),
    .io_in_4_ready(LockingRRArbiter_6_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_6_1_io_in_4_valid),
    .io_in_4_bits_addr_beat(LockingRRArbiter_6_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_addr_block(LockingRRArbiter_6_1_io_in_4_bits_addr_block),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_6_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_voluntary(LockingRRArbiter_6_1_io_in_4_bits_voluntary),
    .io_in_4_bits_r_type(LockingRRArbiter_6_1_io_in_4_bits_r_type),
    .io_in_4_bits_data(LockingRRArbiter_6_1_io_in_4_bits_data),
    .io_out_ready(LockingRRArbiter_6_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_6_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_6_1_io_out_bits_addr_beat),
    .io_out_bits_addr_block(LockingRRArbiter_6_1_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_6_1_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(LockingRRArbiter_6_1_io_out_bits_voluntary),
    .io_out_bits_r_type(LockingRRArbiter_6_1_io_out_bits_r_type),
    .io_out_bits_data(LockingRRArbiter_6_1_io_out_bits_data),
    .io_chosen(LockingRRArbiter_6_1_io_chosen)
  );
  assign io_in_0_acquire_ready = LockingRRArbiter_5_1_io_in_0_ready;
  assign io_in_0_probe_valid = io_out_probe_valid;
  assign io_in_0_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_0_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_0_release_ready = LockingRRArbiter_6_1_io_in_0_ready;
  assign io_in_0_grant_valid = GEN_0;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = 3'h0;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_0_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_0_finish_ready = GEN_10;
  assign io_in_1_acquire_ready = LockingRRArbiter_5_1_io_in_1_ready;
  assign io_in_1_probe_valid = io_out_probe_valid;
  assign io_in_1_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_1_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_1_release_ready = LockingRRArbiter_6_1_io_in_1_ready;
  assign io_in_1_grant_valid = GEN_2;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_bits_client_xact_id = 3'h0;
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_1_finish_ready = GEN_11;
  assign io_in_2_acquire_ready = LockingRRArbiter_5_1_io_in_2_ready;
  assign io_in_2_probe_valid = io_out_probe_valid;
  assign io_in_2_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_2_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_2_release_ready = LockingRRArbiter_6_1_io_in_2_ready;
  assign io_in_2_grant_valid = GEN_4;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_bits_client_xact_id = 3'h0;
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_2_finish_ready = GEN_12;
  assign io_in_3_acquire_ready = LockingRRArbiter_5_1_io_in_3_ready;
  assign io_in_3_probe_valid = io_out_probe_valid;
  assign io_in_3_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_3_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_3_release_ready = LockingRRArbiter_6_1_io_in_3_ready;
  assign io_in_3_grant_valid = GEN_6;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_bits_client_xact_id = 3'h0;
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_3_finish_ready = GEN_13;
  assign io_in_4_acquire_ready = LockingRRArbiter_5_1_io_in_4_ready;
  assign io_in_4_probe_valid = io_out_probe_valid;
  assign io_in_4_probe_bits_addr_block = io_out_probe_bits_addr_block;
  assign io_in_4_probe_bits_p_type = io_out_probe_bits_p_type;
  assign io_in_4_release_ready = LockingRRArbiter_6_1_io_in_4_ready;
  assign io_in_4_grant_valid = GEN_8;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_bits_client_xact_id = 3'h0;
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_grant_bits_manager_id = io_out_grant_bits_manager_id;
  assign io_in_4_finish_ready = GEN_14;
  assign io_out_acquire_valid = LockingRRArbiter_5_1_io_out_valid;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_5_1_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_5_1_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_5_1_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_5_1_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_5_1_io_out_bits_a_type;
  assign io_out_acquire_bits_union = LockingRRArbiter_5_1_io_out_bits_union;
  assign io_out_acquire_bits_data = LockingRRArbiter_5_1_io_out_bits_data;
  assign io_out_probe_ready = T_9062;
  assign io_out_release_valid = LockingRRArbiter_6_1_io_out_valid;
  assign io_out_release_bits_addr_beat = LockingRRArbiter_6_1_io_out_bits_addr_beat;
  assign io_out_release_bits_addr_block = LockingRRArbiter_6_1_io_out_bits_addr_block;
  assign io_out_release_bits_client_xact_id = LockingRRArbiter_6_1_io_out_bits_client_xact_id;
  assign io_out_release_bits_voluntary = LockingRRArbiter_6_1_io_out_bits_voluntary;
  assign io_out_release_bits_r_type = LockingRRArbiter_6_1_io_out_bits_r_type;
  assign io_out_release_bits_data = LockingRRArbiter_6_1_io_out_bits_data;
  assign io_out_grant_ready = GEN_9;
  assign io_out_finish_valid = GEN_15;
  assign io_out_finish_bits_manager_xact_id = GEN_16;
  assign io_out_finish_bits_manager_id = GEN_17;
  assign LockingRRArbiter_5_1_clk = clk;
  assign LockingRRArbiter_5_1_reset = reset;
  assign LockingRRArbiter_5_1_io_in_0_valid = io_in_0_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_0_bits_client_xact_id = T_9040[2:0];
  assign LockingRRArbiter_5_1_io_in_0_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_0_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_a_type = io_in_0_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_0_bits_union = io_in_0_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_0_bits_data = io_in_0_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_1_valid = io_in_1_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_block = io_in_1_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_1_bits_client_xact_id = T_9042[2:0];
  assign LockingRRArbiter_5_1_io_in_1_bits_addr_beat = io_in_1_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_1_bits_is_builtin_type = io_in_1_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_a_type = io_in_1_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_1_bits_union = io_in_1_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_1_bits_data = io_in_1_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_2_valid = io_in_2_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_block = io_in_2_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_2_bits_client_xact_id = T_9044[2:0];
  assign LockingRRArbiter_5_1_io_in_2_bits_addr_beat = io_in_2_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_2_bits_is_builtin_type = io_in_2_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_a_type = io_in_2_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_2_bits_union = io_in_2_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_2_bits_data = io_in_2_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_3_valid = io_in_3_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_3_bits_addr_block = io_in_3_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_3_bits_client_xact_id = T_9046[2:0];
  assign LockingRRArbiter_5_1_io_in_3_bits_addr_beat = io_in_3_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_3_bits_is_builtin_type = io_in_3_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_3_bits_a_type = io_in_3_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_3_bits_union = io_in_3_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_3_bits_data = io_in_3_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_in_4_valid = io_in_4_acquire_valid;
  assign LockingRRArbiter_5_1_io_in_4_bits_addr_block = io_in_4_acquire_bits_addr_block;
  assign LockingRRArbiter_5_1_io_in_4_bits_client_xact_id = T_9048[2:0];
  assign LockingRRArbiter_5_1_io_in_4_bits_addr_beat = io_in_4_acquire_bits_addr_beat;
  assign LockingRRArbiter_5_1_io_in_4_bits_is_builtin_type = io_in_4_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_5_1_io_in_4_bits_a_type = io_in_4_acquire_bits_a_type;
  assign LockingRRArbiter_5_1_io_in_4_bits_union = io_in_4_acquire_bits_union;
  assign LockingRRArbiter_5_1_io_in_4_bits_data = io_in_4_acquire_bits_data;
  assign LockingRRArbiter_5_1_io_out_ready = io_out_acquire_ready;
  assign T_9040 = {io_in_0_acquire_bits_client_xact_id,3'h0};
  assign T_9042 = {io_in_1_acquire_bits_client_xact_id,3'h1};
  assign T_9044 = {io_in_2_acquire_bits_client_xact_id,3'h2};
  assign T_9046 = {io_in_3_acquire_bits_client_xact_id,3'h3};
  assign T_9048 = {io_in_4_acquire_bits_client_xact_id,3'h4};
  assign LockingRRArbiter_6_1_clk = clk;
  assign LockingRRArbiter_6_1_reset = reset;
  assign LockingRRArbiter_6_1_io_in_0_valid = io_in_0_release_valid;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_beat = io_in_0_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_0_bits_addr_block = io_in_0_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_0_bits_client_xact_id = T_9050[2:0];
  assign LockingRRArbiter_6_1_io_in_0_bits_voluntary = io_in_0_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_0_bits_r_type = io_in_0_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_0_bits_data = io_in_0_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_1_valid = io_in_1_release_valid;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_beat = io_in_1_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_1_bits_addr_block = io_in_1_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_1_bits_client_xact_id = T_9052[2:0];
  assign LockingRRArbiter_6_1_io_in_1_bits_voluntary = io_in_1_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_1_bits_r_type = io_in_1_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_1_bits_data = io_in_1_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_2_valid = io_in_2_release_valid;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_beat = io_in_2_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_2_bits_addr_block = io_in_2_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_2_bits_client_xact_id = T_9054[2:0];
  assign LockingRRArbiter_6_1_io_in_2_bits_voluntary = io_in_2_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_2_bits_r_type = io_in_2_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_2_bits_data = io_in_2_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_3_valid = io_in_3_release_valid;
  assign LockingRRArbiter_6_1_io_in_3_bits_addr_beat = io_in_3_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_3_bits_addr_block = io_in_3_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_3_bits_client_xact_id = T_9056[2:0];
  assign LockingRRArbiter_6_1_io_in_3_bits_voluntary = io_in_3_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_3_bits_r_type = io_in_3_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_3_bits_data = io_in_3_release_bits_data;
  assign LockingRRArbiter_6_1_io_in_4_valid = io_in_4_release_valid;
  assign LockingRRArbiter_6_1_io_in_4_bits_addr_beat = io_in_4_release_bits_addr_beat;
  assign LockingRRArbiter_6_1_io_in_4_bits_addr_block = io_in_4_release_bits_addr_block;
  assign LockingRRArbiter_6_1_io_in_4_bits_client_xact_id = T_9058[2:0];
  assign LockingRRArbiter_6_1_io_in_4_bits_voluntary = io_in_4_release_bits_voluntary;
  assign LockingRRArbiter_6_1_io_in_4_bits_r_type = io_in_4_release_bits_r_type;
  assign LockingRRArbiter_6_1_io_in_4_bits_data = io_in_4_release_bits_data;
  assign LockingRRArbiter_6_1_io_out_ready = io_out_release_ready;
  assign T_9050 = {io_in_0_release_bits_client_xact_id,3'h0};
  assign T_9052 = {io_in_1_release_bits_client_xact_id,3'h1};
  assign T_9054 = {io_in_2_release_bits_client_xact_id,3'h2};
  assign T_9056 = {io_in_3_release_bits_client_xact_id,3'h3};
  assign T_9058 = {io_in_4_release_bits_client_xact_id,3'h4};
  assign T_9059 = io_in_0_probe_ready & io_in_1_probe_ready;
  assign T_9060 = T_9059 & io_in_2_probe_ready;
  assign T_9061 = T_9060 & io_in_3_probe_ready;
  assign T_9062 = T_9061 & io_in_4_probe_ready;
  assign T_9067 = io_out_grant_bits_client_xact_id == 3'h0;
  assign GEN_0 = T_9067 ? io_out_grant_valid : 1'h0;
  assign GEN_1 = T_9067 ? io_in_0_grant_ready : 1'h0;
  assign T_9072 = io_out_grant_bits_client_xact_id == 3'h1;
  assign GEN_2 = T_9072 ? io_out_grant_valid : 1'h0;
  assign GEN_3 = T_9072 ? io_in_1_grant_ready : GEN_1;
  assign T_9077 = io_out_grant_bits_client_xact_id == 3'h2;
  assign GEN_4 = T_9077 ? io_out_grant_valid : 1'h0;
  assign GEN_5 = T_9077 ? io_in_2_grant_ready : GEN_3;
  assign T_9082 = io_out_grant_bits_client_xact_id == 3'h3;
  assign GEN_6 = T_9082 ? io_out_grant_valid : 1'h0;
  assign GEN_7 = T_9082 ? io_in_3_grant_ready : GEN_5;
  assign T_9087 = io_out_grant_bits_client_xact_id == 3'h4;
  assign GEN_8 = T_9087 ? io_out_grant_valid : 1'h0;
  assign GEN_9 = T_9087 ? io_in_4_grant_ready : GEN_7;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_11 = GEN_19[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_12 = GEN_20[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_13 = GEN_21[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_14 = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_15 = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_16 = GEN_24[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_25[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_18 = {1{$random}};
  GEN_19 = {1{$random}};
  GEN_20 = {1{$random}};
  GEN_21 = {1{$random}};
  GEN_22 = {1{$random}};
  GEN_23 = {1{$random}};
  GEN_24 = {1{$random}};
  GEN_25 = {1{$random}};
  end
`endif
endmodule
module LockingRRArbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_p_type,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_p_type,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_p_type,
  input   io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [1:0] io_in_3_bits_p_type,
  input   io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [1:0] io_in_4_bits_p_type,
  input   io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_p_type,
  output  io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [1:0] GEN_0_bits_p_type;
  wire  GEN_0_bits_client_id;
  wire  GEN_4;
  wire  GEN_5;
  wire [25:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire [25:0] GEN_16;
  wire [1:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [25:0] GEN_21;
  wire [1:0] GEN_22;
  wire  GEN_23;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [1:0] GEN_1_bits_p_type;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [1:0] GEN_2_bits_p_type;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [1:0] GEN_3_bits_p_type;
  wire  GEN_3_bits_client_id;
  reg [2:0] T_962;
  reg [31:0] GEN_0;
  reg [2:0] T_964;
  reg [31:0] GEN_1;
  wire  T_966;
  wire  T_968;
  wire [2:0] GEN_86;
  reg [2:0] lastGrant;
  reg [31:0] GEN_2;
  wire [2:0] GEN_87;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  grantMask_4;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  validMask_4;
  wire  T_983;
  wire  T_984;
  wire  T_985;
  wire  T_986;
  wire  T_987;
  wire  T_988;
  wire  T_989;
  wire  T_993;
  wire  T_995;
  wire  T_997;
  wire  T_999;
  wire  T_1001;
  wire  T_1003;
  wire  T_1005;
  wire  T_1007;
  wire  T_1011;
  wire  T_1012;
  wire  T_1013;
  wire  T_1014;
  wire  T_1015;
  wire  T_1016;
  wire  T_1017;
  wire  T_1019;
  wire  T_1020;
  wire  T_1021;
  wire  T_1023;
  wire  T_1024;
  wire  T_1025;
  wire  T_1027;
  wire  T_1028;
  wire  T_1029;
  wire  T_1031;
  wire  T_1032;
  wire  T_1033;
  wire  T_1035;
  wire  T_1036;
  wire  T_1037;
  wire [2:0] GEN_88;
  wire [2:0] GEN_89;
  wire [2:0] GEN_90;
  wire [2:0] GEN_91;
  wire [2:0] GEN_92;
  wire [2:0] GEN_93;
  wire [2:0] GEN_94;
  wire [2:0] GEN_95;
  assign io_in_0_ready = T_1021;
  assign io_in_1_ready = T_1025;
  assign io_in_2_ready = T_1029;
  assign io_in_3_ready = T_1033;
  assign io_in_4_ready = T_1037;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_p_type = GEN_2_bits_p_type;
  assign io_out_bits_client_id = GEN_3_bits_client_id;
  assign io_chosen = GEN_86;
  assign choice = GEN_95;
  assign GEN_0_ready = GEN_19;
  assign GEN_0_valid = GEN_20;
  assign GEN_0_bits_addr_block = GEN_21;
  assign GEN_0_bits_p_type = GEN_22;
  assign GEN_0_bits_client_id = GEN_23;
  assign GEN_4 = 3'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_5 = 3'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 3'h1 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_7 = 3'h1 == io_chosen ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign GEN_8 = 3'h1 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_9 = 3'h2 == io_chosen ? io_in_2_ready : GEN_4;
  assign GEN_10 = 3'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_11 = 3'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_6;
  assign GEN_12 = 3'h2 == io_chosen ? io_in_2_bits_p_type : GEN_7;
  assign GEN_13 = 3'h2 == io_chosen ? io_in_2_bits_client_id : GEN_8;
  assign GEN_14 = 3'h3 == io_chosen ? io_in_3_ready : GEN_9;
  assign GEN_15 = 3'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_16 = 3'h3 == io_chosen ? io_in_3_bits_addr_block : GEN_11;
  assign GEN_17 = 3'h3 == io_chosen ? io_in_3_bits_p_type : GEN_12;
  assign GEN_18 = 3'h3 == io_chosen ? io_in_3_bits_client_id : GEN_13;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_ready : GEN_14;
  assign GEN_20 = 3'h4 == io_chosen ? io_in_4_valid : GEN_15;
  assign GEN_21 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_16;
  assign GEN_22 = 3'h4 == io_chosen ? io_in_4_bits_p_type : GEN_17;
  assign GEN_23 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_18;
  assign GEN_1_ready = GEN_19;
  assign GEN_1_valid = GEN_20;
  assign GEN_1_bits_addr_block = GEN_21;
  assign GEN_1_bits_p_type = GEN_22;
  assign GEN_1_bits_client_id = GEN_23;
  assign GEN_2_ready = GEN_19;
  assign GEN_2_valid = GEN_20;
  assign GEN_2_bits_addr_block = GEN_21;
  assign GEN_2_bits_p_type = GEN_22;
  assign GEN_2_bits_client_id = GEN_23;
  assign GEN_3_ready = GEN_19;
  assign GEN_3_valid = GEN_20;
  assign GEN_3_bits_addr_block = GEN_21;
  assign GEN_3_bits_p_type = GEN_22;
  assign GEN_3_bits_client_id = GEN_23;
  assign T_966 = T_962 != 3'h0;
  assign T_968 = io_out_ready & io_out_valid;
  assign GEN_86 = T_966 ? T_964 : choice;
  assign GEN_87 = T_968 ? io_chosen : lastGrant;
  assign grantMask_1 = 3'h1 > lastGrant;
  assign grantMask_2 = 3'h2 > lastGrant;
  assign grantMask_3 = 3'h3 > lastGrant;
  assign grantMask_4 = 3'h4 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign validMask_4 = io_in_4_valid & grantMask_4;
  assign T_983 = validMask_1 | validMask_2;
  assign T_984 = T_983 | validMask_3;
  assign T_985 = T_984 | validMask_4;
  assign T_986 = T_985 | io_in_0_valid;
  assign T_987 = T_986 | io_in_1_valid;
  assign T_988 = T_987 | io_in_2_valid;
  assign T_989 = T_988 | io_in_3_valid;
  assign T_993 = validMask_1 == 1'h0;
  assign T_995 = T_983 == 1'h0;
  assign T_997 = T_984 == 1'h0;
  assign T_999 = T_985 == 1'h0;
  assign T_1001 = T_986 == 1'h0;
  assign T_1003 = T_987 == 1'h0;
  assign T_1005 = T_988 == 1'h0;
  assign T_1007 = T_989 == 1'h0;
  assign T_1011 = grantMask_1 | T_1001;
  assign T_1012 = T_993 & grantMask_2;
  assign T_1013 = T_1012 | T_1003;
  assign T_1014 = T_995 & grantMask_3;
  assign T_1015 = T_1014 | T_1005;
  assign T_1016 = T_997 & grantMask_4;
  assign T_1017 = T_1016 | T_1007;
  assign T_1019 = T_964 == 3'h0;
  assign T_1020 = T_966 ? T_1019 : T_999;
  assign T_1021 = T_1020 & io_out_ready;
  assign T_1023 = T_964 == 3'h1;
  assign T_1024 = T_966 ? T_1023 : T_1011;
  assign T_1025 = T_1024 & io_out_ready;
  assign T_1027 = T_964 == 3'h2;
  assign T_1028 = T_966 ? T_1027 : T_1013;
  assign T_1029 = T_1028 & io_out_ready;
  assign T_1031 = T_964 == 3'h3;
  assign T_1032 = T_966 ? T_1031 : T_1015;
  assign T_1033 = T_1032 & io_out_ready;
  assign T_1035 = T_964 == 3'h4;
  assign T_1036 = T_966 ? T_1035 : T_1017;
  assign T_1037 = T_1036 & io_out_ready;
  assign GEN_88 = io_in_3_valid ? 3'h3 : 3'h4;
  assign GEN_89 = io_in_2_valid ? 3'h2 : GEN_88;
  assign GEN_90 = io_in_1_valid ? 3'h1 : GEN_89;
  assign GEN_91 = io_in_0_valid ? 3'h0 : GEN_90;
  assign GEN_92 = validMask_4 ? 3'h4 : GEN_91;
  assign GEN_93 = validMask_3 ? 3'h3 : GEN_92;
  assign GEN_94 = validMask_2 ? 3'h2 : GEN_93;
  assign GEN_95 = validMask_1 ? 3'h1 : GEN_94;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_962 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_964 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_962 <= 3'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(T_968) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module LockingRRArbiter_8(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  input   io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input   io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [1:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_manager_xact_id,
  input   io_in_4_bits_is_builtin_type,
  input  [3:0] io_in_4_bits_g_type,
  input  [63:0] io_in_4_bits_data,
  input   io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_0_bits_client_id;
  wire  GEN_8;
  wire  GEN_9;
  wire [2:0] GEN_10;
  wire [1:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [3:0] GEN_14;
  wire [63:0] GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [3:0] GEN_23;
  wire [63:0] GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [2:0] GEN_28;
  wire [1:0] GEN_29;
  wire [2:0] GEN_30;
  wire  GEN_31;
  wire [3:0] GEN_32;
  wire [63:0] GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [2:0] GEN_37;
  wire [1:0] GEN_38;
  wire [2:0] GEN_39;
  wire  GEN_40;
  wire [3:0] GEN_41;
  wire [63:0] GEN_42;
  wire  GEN_43;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_3_bits_client_id;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_4_bits_client_id;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_5_bits_client_id;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_6_bits_client_id;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [2:0] GEN_7_bits_addr_beat;
  wire [1:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_manager_xact_id;
  wire  GEN_7_bits_is_builtin_type;
  wire [3:0] GEN_7_bits_g_type;
  wire [63:0] GEN_7_bits_data;
  wire  GEN_7_bits_client_id;
  reg [2:0] T_1114;
  reg [31:0] GEN_1;
  reg [2:0] T_1116;
  reg [31:0] GEN_2;
  wire  T_1118;
  wire [2:0] T_1126_0;
  wire [3:0] GEN_0;
  wire  T_1128;
  wire  T_1129;
  wire  T_1130;
  wire  T_1132;
  wire  T_1133;
  wire [3:0] T_1137;
  wire [2:0] T_1138;
  wire [2:0] GEN_296;
  wire [2:0] GEN_297;
  wire [2:0] GEN_298;
  reg [2:0] lastGrant;
  reg [31:0] GEN_3;
  wire [2:0] GEN_299;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  grantMask_4;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  validMask_4;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire  T_1157;
  wire  T_1159;
  wire  T_1161;
  wire  T_1163;
  wire  T_1165;
  wire  T_1167;
  wire  T_1169;
  wire  T_1171;
  wire  T_1175;
  wire  T_1176;
  wire  T_1177;
  wire  T_1178;
  wire  T_1179;
  wire  T_1180;
  wire  T_1181;
  wire  T_1183;
  wire  T_1184;
  wire  T_1185;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1191;
  wire  T_1192;
  wire  T_1193;
  wire  T_1195;
  wire  T_1196;
  wire  T_1197;
  wire  T_1199;
  wire  T_1200;
  wire  T_1201;
  wire [2:0] GEN_300;
  wire [2:0] GEN_301;
  wire [2:0] GEN_302;
  wire [2:0] GEN_303;
  wire [2:0] GEN_304;
  wire [2:0] GEN_305;
  wire [2:0] GEN_306;
  wire [2:0] GEN_307;
  assign io_in_0_ready = T_1185;
  assign io_in_1_ready = T_1189;
  assign io_in_2_ready = T_1193;
  assign io_in_3_ready = T_1197;
  assign io_in_4_ready = T_1201;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_out_bits_client_id = GEN_7_bits_client_id;
  assign io_chosen = GEN_298;
  assign choice = GEN_307;
  assign GEN_0_ready = GEN_35;
  assign GEN_0_valid = GEN_36;
  assign GEN_0_bits_addr_beat = GEN_37;
  assign GEN_0_bits_client_xact_id = GEN_38;
  assign GEN_0_bits_manager_xact_id = GEN_39;
  assign GEN_0_bits_is_builtin_type = GEN_40;
  assign GEN_0_bits_g_type = GEN_41;
  assign GEN_0_bits_data = GEN_42;
  assign GEN_0_bits_client_id = GEN_43;
  assign GEN_8 = 3'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = 3'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 3'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_11 = 3'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = 3'h1 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_13 = 3'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = 3'h1 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_15 = 3'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_16 = 3'h1 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_17 = 3'h2 == io_chosen ? io_in_2_ready : GEN_8;
  assign GEN_18 = 3'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_19 = 3'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_10;
  assign GEN_20 = 3'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_11;
  assign GEN_21 = 3'h2 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_12;
  assign GEN_22 = 3'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_13;
  assign GEN_23 = 3'h2 == io_chosen ? io_in_2_bits_g_type : GEN_14;
  assign GEN_24 = 3'h2 == io_chosen ? io_in_2_bits_data : GEN_15;
  assign GEN_25 = 3'h2 == io_chosen ? io_in_2_bits_client_id : GEN_16;
  assign GEN_26 = 3'h3 == io_chosen ? io_in_3_ready : GEN_17;
  assign GEN_27 = 3'h3 == io_chosen ? io_in_3_valid : GEN_18;
  assign GEN_28 = 3'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_19;
  assign GEN_29 = 3'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_20;
  assign GEN_30 = 3'h3 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_21;
  assign GEN_31 = 3'h3 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_22;
  assign GEN_32 = 3'h3 == io_chosen ? io_in_3_bits_g_type : GEN_23;
  assign GEN_33 = 3'h3 == io_chosen ? io_in_3_bits_data : GEN_24;
  assign GEN_34 = 3'h3 == io_chosen ? io_in_3_bits_client_id : GEN_25;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_ready : GEN_26;
  assign GEN_36 = 3'h4 == io_chosen ? io_in_4_valid : GEN_27;
  assign GEN_37 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_28;
  assign GEN_38 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_29;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_manager_xact_id : GEN_30;
  assign GEN_40 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_31;
  assign GEN_41 = 3'h4 == io_chosen ? io_in_4_bits_g_type : GEN_32;
  assign GEN_42 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_33;
  assign GEN_43 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_34;
  assign GEN_1_ready = GEN_35;
  assign GEN_1_valid = GEN_36;
  assign GEN_1_bits_addr_beat = GEN_37;
  assign GEN_1_bits_client_xact_id = GEN_38;
  assign GEN_1_bits_manager_xact_id = GEN_39;
  assign GEN_1_bits_is_builtin_type = GEN_40;
  assign GEN_1_bits_g_type = GEN_41;
  assign GEN_1_bits_data = GEN_42;
  assign GEN_1_bits_client_id = GEN_43;
  assign GEN_2_ready = GEN_35;
  assign GEN_2_valid = GEN_36;
  assign GEN_2_bits_addr_beat = GEN_37;
  assign GEN_2_bits_client_xact_id = GEN_38;
  assign GEN_2_bits_manager_xact_id = GEN_39;
  assign GEN_2_bits_is_builtin_type = GEN_40;
  assign GEN_2_bits_g_type = GEN_41;
  assign GEN_2_bits_data = GEN_42;
  assign GEN_2_bits_client_id = GEN_43;
  assign GEN_3_ready = GEN_35;
  assign GEN_3_valid = GEN_36;
  assign GEN_3_bits_addr_beat = GEN_37;
  assign GEN_3_bits_client_xact_id = GEN_38;
  assign GEN_3_bits_manager_xact_id = GEN_39;
  assign GEN_3_bits_is_builtin_type = GEN_40;
  assign GEN_3_bits_g_type = GEN_41;
  assign GEN_3_bits_data = GEN_42;
  assign GEN_3_bits_client_id = GEN_43;
  assign GEN_4_ready = GEN_35;
  assign GEN_4_valid = GEN_36;
  assign GEN_4_bits_addr_beat = GEN_37;
  assign GEN_4_bits_client_xact_id = GEN_38;
  assign GEN_4_bits_manager_xact_id = GEN_39;
  assign GEN_4_bits_is_builtin_type = GEN_40;
  assign GEN_4_bits_g_type = GEN_41;
  assign GEN_4_bits_data = GEN_42;
  assign GEN_4_bits_client_id = GEN_43;
  assign GEN_5_ready = GEN_35;
  assign GEN_5_valid = GEN_36;
  assign GEN_5_bits_addr_beat = GEN_37;
  assign GEN_5_bits_client_xact_id = GEN_38;
  assign GEN_5_bits_manager_xact_id = GEN_39;
  assign GEN_5_bits_is_builtin_type = GEN_40;
  assign GEN_5_bits_g_type = GEN_41;
  assign GEN_5_bits_data = GEN_42;
  assign GEN_5_bits_client_id = GEN_43;
  assign GEN_6_ready = GEN_35;
  assign GEN_6_valid = GEN_36;
  assign GEN_6_bits_addr_beat = GEN_37;
  assign GEN_6_bits_client_xact_id = GEN_38;
  assign GEN_6_bits_manager_xact_id = GEN_39;
  assign GEN_6_bits_is_builtin_type = GEN_40;
  assign GEN_6_bits_g_type = GEN_41;
  assign GEN_6_bits_data = GEN_42;
  assign GEN_6_bits_client_id = GEN_43;
  assign GEN_7_ready = GEN_35;
  assign GEN_7_valid = GEN_36;
  assign GEN_7_bits_addr_beat = GEN_37;
  assign GEN_7_bits_client_xact_id = GEN_38;
  assign GEN_7_bits_manager_xact_id = GEN_39;
  assign GEN_7_bits_is_builtin_type = GEN_40;
  assign GEN_7_bits_g_type = GEN_41;
  assign GEN_7_bits_data = GEN_42;
  assign GEN_7_bits_client_id = GEN_43;
  assign T_1118 = T_1114 != 3'h0;
  assign T_1126_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1126_0};
  assign T_1128 = io_out_bits_g_type == GEN_0;
  assign T_1129 = io_out_bits_g_type == 4'h0;
  assign T_1130 = io_out_bits_is_builtin_type ? T_1128 : T_1129;
  assign T_1132 = io_out_ready & io_out_valid;
  assign T_1133 = T_1132 & T_1130;
  assign T_1137 = T_1114 + 3'h1;
  assign T_1138 = T_1137[2:0];
  assign GEN_296 = T_1133 ? io_chosen : T_1116;
  assign GEN_297 = T_1133 ? T_1138 : T_1114;
  assign GEN_298 = T_1118 ? T_1116 : choice;
  assign GEN_299 = T_1132 ? io_chosen : lastGrant;
  assign grantMask_1 = 3'h1 > lastGrant;
  assign grantMask_2 = 3'h2 > lastGrant;
  assign grantMask_3 = 3'h3 > lastGrant;
  assign grantMask_4 = 3'h4 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign validMask_4 = io_in_4_valid & grantMask_4;
  assign T_1147 = validMask_1 | validMask_2;
  assign T_1148 = T_1147 | validMask_3;
  assign T_1149 = T_1148 | validMask_4;
  assign T_1150 = T_1149 | io_in_0_valid;
  assign T_1151 = T_1150 | io_in_1_valid;
  assign T_1152 = T_1151 | io_in_2_valid;
  assign T_1153 = T_1152 | io_in_3_valid;
  assign T_1157 = validMask_1 == 1'h0;
  assign T_1159 = T_1147 == 1'h0;
  assign T_1161 = T_1148 == 1'h0;
  assign T_1163 = T_1149 == 1'h0;
  assign T_1165 = T_1150 == 1'h0;
  assign T_1167 = T_1151 == 1'h0;
  assign T_1169 = T_1152 == 1'h0;
  assign T_1171 = T_1153 == 1'h0;
  assign T_1175 = grantMask_1 | T_1165;
  assign T_1176 = T_1157 & grantMask_2;
  assign T_1177 = T_1176 | T_1167;
  assign T_1178 = T_1159 & grantMask_3;
  assign T_1179 = T_1178 | T_1169;
  assign T_1180 = T_1161 & grantMask_4;
  assign T_1181 = T_1180 | T_1171;
  assign T_1183 = T_1116 == 3'h0;
  assign T_1184 = T_1118 ? T_1183 : T_1163;
  assign T_1185 = T_1184 & io_out_ready;
  assign T_1187 = T_1116 == 3'h1;
  assign T_1188 = T_1118 ? T_1187 : T_1175;
  assign T_1189 = T_1188 & io_out_ready;
  assign T_1191 = T_1116 == 3'h2;
  assign T_1192 = T_1118 ? T_1191 : T_1177;
  assign T_1193 = T_1192 & io_out_ready;
  assign T_1195 = T_1116 == 3'h3;
  assign T_1196 = T_1118 ? T_1195 : T_1179;
  assign T_1197 = T_1196 & io_out_ready;
  assign T_1199 = T_1116 == 3'h4;
  assign T_1200 = T_1118 ? T_1199 : T_1181;
  assign T_1201 = T_1200 & io_out_ready;
  assign GEN_300 = io_in_3_valid ? 3'h3 : 3'h4;
  assign GEN_301 = io_in_2_valid ? 3'h2 : GEN_300;
  assign GEN_302 = io_in_1_valid ? 3'h1 : GEN_301;
  assign GEN_303 = io_in_0_valid ? 3'h0 : GEN_302;
  assign GEN_304 = validMask_4 ? 3'h4 : GEN_303;
  assign GEN_305 = validMask_3 ? 3'h3 : GEN_304;
  assign GEN_306 = validMask_2 ? 3'h2 : GEN_305;
  assign GEN_307 = validMask_1 ? 3'h1 : GEN_306;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_1114 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_1116 = GEN_2[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1114 <= 3'h0;
    end else begin
      if(T_1133) begin
        T_1114 <= T_1138;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1133) begin
        T_1116 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1132) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module L2BroadcastHub(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  wire  trackerList_0_clk;
  wire  trackerList_0_reset;
  wire  trackerList_0_io_inner_acquire_ready;
  wire  trackerList_0_io_inner_acquire_valid;
  wire [25:0] trackerList_0_io_inner_acquire_bits_addr_block;
  wire [1:0] trackerList_0_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_0_io_inner_acquire_bits_addr_beat;
  wire  trackerList_0_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_0_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_0_io_inner_acquire_bits_union;
  wire [63:0] trackerList_0_io_inner_acquire_bits_data;
  wire  trackerList_0_io_inner_acquire_bits_client_id;
  wire  trackerList_0_io_inner_grant_ready;
  wire  trackerList_0_io_inner_grant_valid;
  wire [2:0] trackerList_0_io_inner_grant_bits_addr_beat;
  wire [1:0] trackerList_0_io_inner_grant_bits_client_xact_id;
  wire [2:0] trackerList_0_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_0_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_0_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_0_io_inner_grant_bits_data;
  wire  trackerList_0_io_inner_grant_bits_client_id;
  wire  trackerList_0_io_inner_finish_ready;
  wire  trackerList_0_io_inner_finish_valid;
  wire [2:0] trackerList_0_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_0_io_inner_probe_ready;
  wire  trackerList_0_io_inner_probe_valid;
  wire [25:0] trackerList_0_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_0_io_inner_probe_bits_p_type;
  wire  trackerList_0_io_inner_probe_bits_client_id;
  wire  trackerList_0_io_inner_release_ready;
  wire  trackerList_0_io_inner_release_valid;
  wire [2:0] trackerList_0_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_0_io_inner_release_bits_addr_block;
  wire [1:0] trackerList_0_io_inner_release_bits_client_xact_id;
  wire  trackerList_0_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_0_io_inner_release_bits_r_type;
  wire [63:0] trackerList_0_io_inner_release_bits_data;
  wire  trackerList_0_io_inner_release_bits_client_id;
  wire  trackerList_0_io_incoherent_0;
  wire  trackerList_0_io_outer_acquire_ready;
  wire  trackerList_0_io_outer_acquire_valid;
  wire [25:0] trackerList_0_io_outer_acquire_bits_addr_block;
  wire [2:0] trackerList_0_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_0_io_outer_acquire_bits_addr_beat;
  wire  trackerList_0_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_0_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_0_io_outer_acquire_bits_union;
  wire [63:0] trackerList_0_io_outer_acquire_bits_data;
  wire  trackerList_0_io_outer_probe_ready;
  wire  trackerList_0_io_outer_probe_valid;
  wire [25:0] trackerList_0_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_0_io_outer_probe_bits_p_type;
  wire  trackerList_0_io_outer_release_ready;
  wire  trackerList_0_io_outer_release_valid;
  wire [2:0] trackerList_0_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_0_io_outer_release_bits_addr_block;
  wire [2:0] trackerList_0_io_outer_release_bits_client_xact_id;
  wire  trackerList_0_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_0_io_outer_release_bits_r_type;
  wire [63:0] trackerList_0_io_outer_release_bits_data;
  wire  trackerList_0_io_outer_grant_ready;
  wire  trackerList_0_io_outer_grant_valid;
  wire [2:0] trackerList_0_io_outer_grant_bits_addr_beat;
  wire [2:0] trackerList_0_io_outer_grant_bits_client_xact_id;
  wire  trackerList_0_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_0_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_0_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_0_io_outer_grant_bits_data;
  wire  trackerList_0_io_outer_grant_bits_manager_id;
  wire  trackerList_0_io_outer_finish_ready;
  wire  trackerList_0_io_outer_finish_valid;
  wire  trackerList_0_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_0_io_outer_finish_bits_manager_id;
  wire  trackerList_0_io_alloc_iacq_matches;
  wire  trackerList_0_io_alloc_iacq_can;
  wire  trackerList_0_io_alloc_iacq_should;
  wire  trackerList_0_io_alloc_irel_matches;
  wire  trackerList_0_io_alloc_irel_can;
  wire  trackerList_0_io_alloc_irel_should;
  wire  trackerList_0_io_alloc_oprb_matches;
  wire  trackerList_0_io_alloc_oprb_can;
  wire  trackerList_0_io_alloc_oprb_should;
  wire  trackerList_0_io_alloc_idle;
  wire [25:0] trackerList_0_io_alloc_addr_block;
  wire  trackerList_1_clk;
  wire  trackerList_1_reset;
  wire  trackerList_1_io_inner_acquire_ready;
  wire  trackerList_1_io_inner_acquire_valid;
  wire [25:0] trackerList_1_io_inner_acquire_bits_addr_block;
  wire [1:0] trackerList_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_1_io_inner_acquire_bits_addr_beat;
  wire  trackerList_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_1_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_1_io_inner_acquire_bits_union;
  wire [63:0] trackerList_1_io_inner_acquire_bits_data;
  wire  trackerList_1_io_inner_acquire_bits_client_id;
  wire  trackerList_1_io_inner_grant_ready;
  wire  trackerList_1_io_inner_grant_valid;
  wire [2:0] trackerList_1_io_inner_grant_bits_addr_beat;
  wire [1:0] trackerList_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] trackerList_1_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_1_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_1_io_inner_grant_bits_data;
  wire  trackerList_1_io_inner_grant_bits_client_id;
  wire  trackerList_1_io_inner_finish_ready;
  wire  trackerList_1_io_inner_finish_valid;
  wire [2:0] trackerList_1_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_1_io_inner_probe_ready;
  wire  trackerList_1_io_inner_probe_valid;
  wire [25:0] trackerList_1_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_1_io_inner_probe_bits_p_type;
  wire  trackerList_1_io_inner_probe_bits_client_id;
  wire  trackerList_1_io_inner_release_ready;
  wire  trackerList_1_io_inner_release_valid;
  wire [2:0] trackerList_1_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_1_io_inner_release_bits_addr_block;
  wire [1:0] trackerList_1_io_inner_release_bits_client_xact_id;
  wire  trackerList_1_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_1_io_inner_release_bits_r_type;
  wire [63:0] trackerList_1_io_inner_release_bits_data;
  wire  trackerList_1_io_inner_release_bits_client_id;
  wire  trackerList_1_io_incoherent_0;
  wire  trackerList_1_io_outer_acquire_ready;
  wire  trackerList_1_io_outer_acquire_valid;
  wire [25:0] trackerList_1_io_outer_acquire_bits_addr_block;
  wire [2:0] trackerList_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_1_io_outer_acquire_bits_addr_beat;
  wire  trackerList_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_1_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_1_io_outer_acquire_bits_union;
  wire [63:0] trackerList_1_io_outer_acquire_bits_data;
  wire  trackerList_1_io_outer_probe_ready;
  wire  trackerList_1_io_outer_probe_valid;
  wire [25:0] trackerList_1_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_1_io_outer_probe_bits_p_type;
  wire  trackerList_1_io_outer_release_ready;
  wire  trackerList_1_io_outer_release_valid;
  wire [2:0] trackerList_1_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_1_io_outer_release_bits_addr_block;
  wire [2:0] trackerList_1_io_outer_release_bits_client_xact_id;
  wire  trackerList_1_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_1_io_outer_release_bits_r_type;
  wire [63:0] trackerList_1_io_outer_release_bits_data;
  wire  trackerList_1_io_outer_grant_ready;
  wire  trackerList_1_io_outer_grant_valid;
  wire [2:0] trackerList_1_io_outer_grant_bits_addr_beat;
  wire [2:0] trackerList_1_io_outer_grant_bits_client_xact_id;
  wire  trackerList_1_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_1_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_1_io_outer_grant_bits_data;
  wire  trackerList_1_io_outer_grant_bits_manager_id;
  wire  trackerList_1_io_outer_finish_ready;
  wire  trackerList_1_io_outer_finish_valid;
  wire  trackerList_1_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_1_io_outer_finish_bits_manager_id;
  wire  trackerList_1_io_alloc_iacq_matches;
  wire  trackerList_1_io_alloc_iacq_can;
  wire  trackerList_1_io_alloc_iacq_should;
  wire  trackerList_1_io_alloc_irel_matches;
  wire  trackerList_1_io_alloc_irel_can;
  wire  trackerList_1_io_alloc_irel_should;
  wire  trackerList_1_io_alloc_oprb_matches;
  wire  trackerList_1_io_alloc_oprb_can;
  wire  trackerList_1_io_alloc_oprb_should;
  wire  trackerList_1_io_alloc_idle;
  wire [25:0] trackerList_1_io_alloc_addr_block;
  wire  trackerList_2_clk;
  wire  trackerList_2_reset;
  wire  trackerList_2_io_inner_acquire_ready;
  wire  trackerList_2_io_inner_acquire_valid;
  wire [25:0] trackerList_2_io_inner_acquire_bits_addr_block;
  wire [1:0] trackerList_2_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_2_io_inner_acquire_bits_addr_beat;
  wire  trackerList_2_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_2_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_2_io_inner_acquire_bits_union;
  wire [63:0] trackerList_2_io_inner_acquire_bits_data;
  wire  trackerList_2_io_inner_acquire_bits_client_id;
  wire  trackerList_2_io_inner_grant_ready;
  wire  trackerList_2_io_inner_grant_valid;
  wire [2:0] trackerList_2_io_inner_grant_bits_addr_beat;
  wire [1:0] trackerList_2_io_inner_grant_bits_client_xact_id;
  wire [2:0] trackerList_2_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_2_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_2_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_2_io_inner_grant_bits_data;
  wire  trackerList_2_io_inner_grant_bits_client_id;
  wire  trackerList_2_io_inner_finish_ready;
  wire  trackerList_2_io_inner_finish_valid;
  wire [2:0] trackerList_2_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_2_io_inner_probe_ready;
  wire  trackerList_2_io_inner_probe_valid;
  wire [25:0] trackerList_2_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_2_io_inner_probe_bits_p_type;
  wire  trackerList_2_io_inner_probe_bits_client_id;
  wire  trackerList_2_io_inner_release_ready;
  wire  trackerList_2_io_inner_release_valid;
  wire [2:0] trackerList_2_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_2_io_inner_release_bits_addr_block;
  wire [1:0] trackerList_2_io_inner_release_bits_client_xact_id;
  wire  trackerList_2_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_2_io_inner_release_bits_r_type;
  wire [63:0] trackerList_2_io_inner_release_bits_data;
  wire  trackerList_2_io_inner_release_bits_client_id;
  wire  trackerList_2_io_incoherent_0;
  wire  trackerList_2_io_outer_acquire_ready;
  wire  trackerList_2_io_outer_acquire_valid;
  wire [25:0] trackerList_2_io_outer_acquire_bits_addr_block;
  wire [2:0] trackerList_2_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_2_io_outer_acquire_bits_addr_beat;
  wire  trackerList_2_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_2_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_2_io_outer_acquire_bits_union;
  wire [63:0] trackerList_2_io_outer_acquire_bits_data;
  wire  trackerList_2_io_outer_probe_ready;
  wire  trackerList_2_io_outer_probe_valid;
  wire [25:0] trackerList_2_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_2_io_outer_probe_bits_p_type;
  wire  trackerList_2_io_outer_release_ready;
  wire  trackerList_2_io_outer_release_valid;
  wire [2:0] trackerList_2_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_2_io_outer_release_bits_addr_block;
  wire [2:0] trackerList_2_io_outer_release_bits_client_xact_id;
  wire  trackerList_2_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_2_io_outer_release_bits_r_type;
  wire [63:0] trackerList_2_io_outer_release_bits_data;
  wire  trackerList_2_io_outer_grant_ready;
  wire  trackerList_2_io_outer_grant_valid;
  wire [2:0] trackerList_2_io_outer_grant_bits_addr_beat;
  wire [2:0] trackerList_2_io_outer_grant_bits_client_xact_id;
  wire  trackerList_2_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_2_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_2_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_2_io_outer_grant_bits_data;
  wire  trackerList_2_io_outer_grant_bits_manager_id;
  wire  trackerList_2_io_outer_finish_ready;
  wire  trackerList_2_io_outer_finish_valid;
  wire  trackerList_2_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_2_io_outer_finish_bits_manager_id;
  wire  trackerList_2_io_alloc_iacq_matches;
  wire  trackerList_2_io_alloc_iacq_can;
  wire  trackerList_2_io_alloc_iacq_should;
  wire  trackerList_2_io_alloc_irel_matches;
  wire  trackerList_2_io_alloc_irel_can;
  wire  trackerList_2_io_alloc_irel_should;
  wire  trackerList_2_io_alloc_oprb_matches;
  wire  trackerList_2_io_alloc_oprb_can;
  wire  trackerList_2_io_alloc_oprb_should;
  wire  trackerList_2_io_alloc_idle;
  wire [25:0] trackerList_2_io_alloc_addr_block;
  wire  trackerList_3_clk;
  wire  trackerList_3_reset;
  wire  trackerList_3_io_inner_acquire_ready;
  wire  trackerList_3_io_inner_acquire_valid;
  wire [25:0] trackerList_3_io_inner_acquire_bits_addr_block;
  wire [1:0] trackerList_3_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_3_io_inner_acquire_bits_addr_beat;
  wire  trackerList_3_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_3_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_3_io_inner_acquire_bits_union;
  wire [63:0] trackerList_3_io_inner_acquire_bits_data;
  wire  trackerList_3_io_inner_acquire_bits_client_id;
  wire  trackerList_3_io_inner_grant_ready;
  wire  trackerList_3_io_inner_grant_valid;
  wire [2:0] trackerList_3_io_inner_grant_bits_addr_beat;
  wire [1:0] trackerList_3_io_inner_grant_bits_client_xact_id;
  wire [2:0] trackerList_3_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_3_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_3_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_3_io_inner_grant_bits_data;
  wire  trackerList_3_io_inner_grant_bits_client_id;
  wire  trackerList_3_io_inner_finish_ready;
  wire  trackerList_3_io_inner_finish_valid;
  wire [2:0] trackerList_3_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_3_io_inner_probe_ready;
  wire  trackerList_3_io_inner_probe_valid;
  wire [25:0] trackerList_3_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_3_io_inner_probe_bits_p_type;
  wire  trackerList_3_io_inner_probe_bits_client_id;
  wire  trackerList_3_io_inner_release_ready;
  wire  trackerList_3_io_inner_release_valid;
  wire [2:0] trackerList_3_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_3_io_inner_release_bits_addr_block;
  wire [1:0] trackerList_3_io_inner_release_bits_client_xact_id;
  wire  trackerList_3_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_3_io_inner_release_bits_r_type;
  wire [63:0] trackerList_3_io_inner_release_bits_data;
  wire  trackerList_3_io_inner_release_bits_client_id;
  wire  trackerList_3_io_incoherent_0;
  wire  trackerList_3_io_outer_acquire_ready;
  wire  trackerList_3_io_outer_acquire_valid;
  wire [25:0] trackerList_3_io_outer_acquire_bits_addr_block;
  wire [2:0] trackerList_3_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_3_io_outer_acquire_bits_addr_beat;
  wire  trackerList_3_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_3_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_3_io_outer_acquire_bits_union;
  wire [63:0] trackerList_3_io_outer_acquire_bits_data;
  wire  trackerList_3_io_outer_probe_ready;
  wire  trackerList_3_io_outer_probe_valid;
  wire [25:0] trackerList_3_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_3_io_outer_probe_bits_p_type;
  wire  trackerList_3_io_outer_release_ready;
  wire  trackerList_3_io_outer_release_valid;
  wire [2:0] trackerList_3_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_3_io_outer_release_bits_addr_block;
  wire [2:0] trackerList_3_io_outer_release_bits_client_xact_id;
  wire  trackerList_3_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_3_io_outer_release_bits_r_type;
  wire [63:0] trackerList_3_io_outer_release_bits_data;
  wire  trackerList_3_io_outer_grant_ready;
  wire  trackerList_3_io_outer_grant_valid;
  wire [2:0] trackerList_3_io_outer_grant_bits_addr_beat;
  wire [2:0] trackerList_3_io_outer_grant_bits_client_xact_id;
  wire  trackerList_3_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_3_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_3_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_3_io_outer_grant_bits_data;
  wire  trackerList_3_io_outer_grant_bits_manager_id;
  wire  trackerList_3_io_outer_finish_ready;
  wire  trackerList_3_io_outer_finish_valid;
  wire  trackerList_3_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_3_io_outer_finish_bits_manager_id;
  wire  trackerList_3_io_alloc_iacq_matches;
  wire  trackerList_3_io_alloc_iacq_can;
  wire  trackerList_3_io_alloc_iacq_should;
  wire  trackerList_3_io_alloc_irel_matches;
  wire  trackerList_3_io_alloc_irel_can;
  wire  trackerList_3_io_alloc_irel_should;
  wire  trackerList_3_io_alloc_oprb_matches;
  wire  trackerList_3_io_alloc_oprb_can;
  wire  trackerList_3_io_alloc_oprb_should;
  wire  trackerList_3_io_alloc_idle;
  wire [25:0] trackerList_3_io_alloc_addr_block;
  wire  trackerList_4_clk;
  wire  trackerList_4_reset;
  wire  trackerList_4_io_inner_acquire_ready;
  wire  trackerList_4_io_inner_acquire_valid;
  wire [25:0] trackerList_4_io_inner_acquire_bits_addr_block;
  wire [1:0] trackerList_4_io_inner_acquire_bits_client_xact_id;
  wire [2:0] trackerList_4_io_inner_acquire_bits_addr_beat;
  wire  trackerList_4_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_4_io_inner_acquire_bits_a_type;
  wire [10:0] trackerList_4_io_inner_acquire_bits_union;
  wire [63:0] trackerList_4_io_inner_acquire_bits_data;
  wire  trackerList_4_io_inner_acquire_bits_client_id;
  wire  trackerList_4_io_inner_grant_ready;
  wire  trackerList_4_io_inner_grant_valid;
  wire [2:0] trackerList_4_io_inner_grant_bits_addr_beat;
  wire [1:0] trackerList_4_io_inner_grant_bits_client_xact_id;
  wire [2:0] trackerList_4_io_inner_grant_bits_manager_xact_id;
  wire  trackerList_4_io_inner_grant_bits_is_builtin_type;
  wire [3:0] trackerList_4_io_inner_grant_bits_g_type;
  wire [63:0] trackerList_4_io_inner_grant_bits_data;
  wire  trackerList_4_io_inner_grant_bits_client_id;
  wire  trackerList_4_io_inner_finish_ready;
  wire  trackerList_4_io_inner_finish_valid;
  wire [2:0] trackerList_4_io_inner_finish_bits_manager_xact_id;
  wire  trackerList_4_io_inner_probe_ready;
  wire  trackerList_4_io_inner_probe_valid;
  wire [25:0] trackerList_4_io_inner_probe_bits_addr_block;
  wire [1:0] trackerList_4_io_inner_probe_bits_p_type;
  wire  trackerList_4_io_inner_probe_bits_client_id;
  wire  trackerList_4_io_inner_release_ready;
  wire  trackerList_4_io_inner_release_valid;
  wire [2:0] trackerList_4_io_inner_release_bits_addr_beat;
  wire [25:0] trackerList_4_io_inner_release_bits_addr_block;
  wire [1:0] trackerList_4_io_inner_release_bits_client_xact_id;
  wire  trackerList_4_io_inner_release_bits_voluntary;
  wire [2:0] trackerList_4_io_inner_release_bits_r_type;
  wire [63:0] trackerList_4_io_inner_release_bits_data;
  wire  trackerList_4_io_inner_release_bits_client_id;
  wire  trackerList_4_io_incoherent_0;
  wire  trackerList_4_io_outer_acquire_ready;
  wire  trackerList_4_io_outer_acquire_valid;
  wire [25:0] trackerList_4_io_outer_acquire_bits_addr_block;
  wire [2:0] trackerList_4_io_outer_acquire_bits_client_xact_id;
  wire [2:0] trackerList_4_io_outer_acquire_bits_addr_beat;
  wire  trackerList_4_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] trackerList_4_io_outer_acquire_bits_a_type;
  wire [10:0] trackerList_4_io_outer_acquire_bits_union;
  wire [63:0] trackerList_4_io_outer_acquire_bits_data;
  wire  trackerList_4_io_outer_probe_ready;
  wire  trackerList_4_io_outer_probe_valid;
  wire [25:0] trackerList_4_io_outer_probe_bits_addr_block;
  wire [1:0] trackerList_4_io_outer_probe_bits_p_type;
  wire  trackerList_4_io_outer_release_ready;
  wire  trackerList_4_io_outer_release_valid;
  wire [2:0] trackerList_4_io_outer_release_bits_addr_beat;
  wire [25:0] trackerList_4_io_outer_release_bits_addr_block;
  wire [2:0] trackerList_4_io_outer_release_bits_client_xact_id;
  wire  trackerList_4_io_outer_release_bits_voluntary;
  wire [2:0] trackerList_4_io_outer_release_bits_r_type;
  wire [63:0] trackerList_4_io_outer_release_bits_data;
  wire  trackerList_4_io_outer_grant_ready;
  wire  trackerList_4_io_outer_grant_valid;
  wire [2:0] trackerList_4_io_outer_grant_bits_addr_beat;
  wire [2:0] trackerList_4_io_outer_grant_bits_client_xact_id;
  wire  trackerList_4_io_outer_grant_bits_manager_xact_id;
  wire  trackerList_4_io_outer_grant_bits_is_builtin_type;
  wire [3:0] trackerList_4_io_outer_grant_bits_g_type;
  wire [63:0] trackerList_4_io_outer_grant_bits_data;
  wire  trackerList_4_io_outer_grant_bits_manager_id;
  wire  trackerList_4_io_outer_finish_ready;
  wire  trackerList_4_io_outer_finish_valid;
  wire  trackerList_4_io_outer_finish_bits_manager_xact_id;
  wire  trackerList_4_io_outer_finish_bits_manager_id;
  wire  trackerList_4_io_alloc_iacq_matches;
  wire  trackerList_4_io_alloc_iacq_can;
  wire  trackerList_4_io_alloc_iacq_should;
  wire  trackerList_4_io_alloc_irel_matches;
  wire  trackerList_4_io_alloc_irel_can;
  wire  trackerList_4_io_alloc_irel_should;
  wire  trackerList_4_io_alloc_oprb_matches;
  wire  trackerList_4_io_alloc_oprb_can;
  wire  trackerList_4_io_alloc_oprb_should;
  wire  trackerList_4_io_alloc_idle;
  wire [25:0] trackerList_4_io_alloc_addr_block;
  wire  outer_arb_clk;
  wire  outer_arb_reset;
  wire  outer_arb_io_in_0_acquire_ready;
  wire  outer_arb_io_in_0_acquire_valid;
  wire [25:0] outer_arb_io_in_0_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_0_acquire_bits_addr_beat;
  wire  outer_arb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_0_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_0_acquire_bits_union;
  wire [63:0] outer_arb_io_in_0_acquire_bits_data;
  wire  outer_arb_io_in_0_probe_ready;
  wire  outer_arb_io_in_0_probe_valid;
  wire [25:0] outer_arb_io_in_0_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_0_probe_bits_p_type;
  wire  outer_arb_io_in_0_release_ready;
  wire  outer_arb_io_in_0_release_valid;
  wire [2:0] outer_arb_io_in_0_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_0_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_0_release_bits_client_xact_id;
  wire  outer_arb_io_in_0_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_0_release_bits_r_type;
  wire [63:0] outer_arb_io_in_0_release_bits_data;
  wire  outer_arb_io_in_0_grant_ready;
  wire  outer_arb_io_in_0_grant_valid;
  wire [2:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire  outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_0_grant_bits_data;
  wire  outer_arb_io_in_0_grant_bits_manager_id;
  wire  outer_arb_io_in_0_finish_ready;
  wire  outer_arb_io_in_0_finish_valid;
  wire  outer_arb_io_in_0_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_0_finish_bits_manager_id;
  wire  outer_arb_io_in_1_acquire_ready;
  wire  outer_arb_io_in_1_acquire_valid;
  wire [25:0] outer_arb_io_in_1_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_1_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_1_acquire_bits_addr_beat;
  wire  outer_arb_io_in_1_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_1_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_1_acquire_bits_union;
  wire [63:0] outer_arb_io_in_1_acquire_bits_data;
  wire  outer_arb_io_in_1_probe_ready;
  wire  outer_arb_io_in_1_probe_valid;
  wire [25:0] outer_arb_io_in_1_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_1_probe_bits_p_type;
  wire  outer_arb_io_in_1_release_ready;
  wire  outer_arb_io_in_1_release_valid;
  wire [2:0] outer_arb_io_in_1_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_1_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_1_release_bits_client_xact_id;
  wire  outer_arb_io_in_1_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_1_release_bits_r_type;
  wire [63:0] outer_arb_io_in_1_release_bits_data;
  wire  outer_arb_io_in_1_grant_ready;
  wire  outer_arb_io_in_1_grant_valid;
  wire [2:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire  outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_1_grant_bits_data;
  wire  outer_arb_io_in_1_grant_bits_manager_id;
  wire  outer_arb_io_in_1_finish_ready;
  wire  outer_arb_io_in_1_finish_valid;
  wire  outer_arb_io_in_1_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_1_finish_bits_manager_id;
  wire  outer_arb_io_in_2_acquire_ready;
  wire  outer_arb_io_in_2_acquire_valid;
  wire [25:0] outer_arb_io_in_2_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_2_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_2_acquire_bits_addr_beat;
  wire  outer_arb_io_in_2_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_2_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_2_acquire_bits_union;
  wire [63:0] outer_arb_io_in_2_acquire_bits_data;
  wire  outer_arb_io_in_2_probe_ready;
  wire  outer_arb_io_in_2_probe_valid;
  wire [25:0] outer_arb_io_in_2_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_2_probe_bits_p_type;
  wire  outer_arb_io_in_2_release_ready;
  wire  outer_arb_io_in_2_release_valid;
  wire [2:0] outer_arb_io_in_2_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_2_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_2_release_bits_client_xact_id;
  wire  outer_arb_io_in_2_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_2_release_bits_r_type;
  wire [63:0] outer_arb_io_in_2_release_bits_data;
  wire  outer_arb_io_in_2_grant_ready;
  wire  outer_arb_io_in_2_grant_valid;
  wire [2:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire  outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_2_grant_bits_data;
  wire  outer_arb_io_in_2_grant_bits_manager_id;
  wire  outer_arb_io_in_2_finish_ready;
  wire  outer_arb_io_in_2_finish_valid;
  wire  outer_arb_io_in_2_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_2_finish_bits_manager_id;
  wire  outer_arb_io_in_3_acquire_ready;
  wire  outer_arb_io_in_3_acquire_valid;
  wire [25:0] outer_arb_io_in_3_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_3_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_3_acquire_bits_addr_beat;
  wire  outer_arb_io_in_3_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_3_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_3_acquire_bits_union;
  wire [63:0] outer_arb_io_in_3_acquire_bits_data;
  wire  outer_arb_io_in_3_probe_ready;
  wire  outer_arb_io_in_3_probe_valid;
  wire [25:0] outer_arb_io_in_3_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_3_probe_bits_p_type;
  wire  outer_arb_io_in_3_release_ready;
  wire  outer_arb_io_in_3_release_valid;
  wire [2:0] outer_arb_io_in_3_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_3_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_3_release_bits_client_xact_id;
  wire  outer_arb_io_in_3_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_3_release_bits_r_type;
  wire [63:0] outer_arb_io_in_3_release_bits_data;
  wire  outer_arb_io_in_3_grant_ready;
  wire  outer_arb_io_in_3_grant_valid;
  wire [2:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire  outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_3_grant_bits_data;
  wire  outer_arb_io_in_3_grant_bits_manager_id;
  wire  outer_arb_io_in_3_finish_ready;
  wire  outer_arb_io_in_3_finish_valid;
  wire  outer_arb_io_in_3_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_3_finish_bits_manager_id;
  wire  outer_arb_io_in_4_acquire_ready;
  wire  outer_arb_io_in_4_acquire_valid;
  wire [25:0] outer_arb_io_in_4_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_4_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_4_acquire_bits_addr_beat;
  wire  outer_arb_io_in_4_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_4_acquire_bits_a_type;
  wire [10:0] outer_arb_io_in_4_acquire_bits_union;
  wire [63:0] outer_arb_io_in_4_acquire_bits_data;
  wire  outer_arb_io_in_4_probe_ready;
  wire  outer_arb_io_in_4_probe_valid;
  wire [25:0] outer_arb_io_in_4_probe_bits_addr_block;
  wire [1:0] outer_arb_io_in_4_probe_bits_p_type;
  wire  outer_arb_io_in_4_release_ready;
  wire  outer_arb_io_in_4_release_valid;
  wire [2:0] outer_arb_io_in_4_release_bits_addr_beat;
  wire [25:0] outer_arb_io_in_4_release_bits_addr_block;
  wire [2:0] outer_arb_io_in_4_release_bits_client_xact_id;
  wire  outer_arb_io_in_4_release_bits_voluntary;
  wire [2:0] outer_arb_io_in_4_release_bits_r_type;
  wire [63:0] outer_arb_io_in_4_release_bits_data;
  wire  outer_arb_io_in_4_grant_ready;
  wire  outer_arb_io_in_4_grant_valid;
  wire [2:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire  outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire [63:0] outer_arb_io_in_4_grant_bits_data;
  wire  outer_arb_io_in_4_grant_bits_manager_id;
  wire  outer_arb_io_in_4_finish_ready;
  wire  outer_arb_io_in_4_finish_valid;
  wire  outer_arb_io_in_4_finish_bits_manager_xact_id;
  wire  outer_arb_io_in_4_finish_bits_manager_id;
  wire  outer_arb_io_out_acquire_ready;
  wire  outer_arb_io_out_acquire_valid;
  wire [25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire  outer_arb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_out_acquire_bits_a_type;
  wire [10:0] outer_arb_io_out_acquire_bits_union;
  wire [63:0] outer_arb_io_out_acquire_bits_data;
  wire  outer_arb_io_out_probe_ready;
  wire  outer_arb_io_out_probe_valid;
  wire [25:0] outer_arb_io_out_probe_bits_addr_block;
  wire [1:0] outer_arb_io_out_probe_bits_p_type;
  wire  outer_arb_io_out_release_ready;
  wire  outer_arb_io_out_release_valid;
  wire [2:0] outer_arb_io_out_release_bits_addr_beat;
  wire [25:0] outer_arb_io_out_release_bits_addr_block;
  wire [2:0] outer_arb_io_out_release_bits_client_xact_id;
  wire  outer_arb_io_out_release_bits_voluntary;
  wire [2:0] outer_arb_io_out_release_bits_r_type;
  wire [63:0] outer_arb_io_out_release_bits_data;
  wire  outer_arb_io_out_grant_ready;
  wire  outer_arb_io_out_grant_valid;
  wire [2:0] outer_arb_io_out_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_out_grant_bits_client_xact_id;
  wire  outer_arb_io_out_grant_bits_manager_xact_id;
  wire  outer_arb_io_out_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_out_grant_bits_g_type;
  wire [63:0] outer_arb_io_out_grant_bits_data;
  wire  outer_arb_io_out_grant_bits_manager_id;
  wire  outer_arb_io_out_finish_ready;
  wire  outer_arb_io_out_finish_valid;
  wire  outer_arb_io_out_finish_bits_manager_xact_id;
  wire  outer_arb_io_out_finish_bits_manager_id;
  wire  T_1215;
  wire  T_1216;
  wire  irel_vs_iacq_conflict;
  wire  T_1218;
  wire [1:0] T_1219;
  wire [1:0] T_1220;
  wire [2:0] T_1221;
  wire [4:0] T_1222;
  wire [1:0] T_1223;
  wire [1:0] T_1224;
  wire [2:0] T_1225;
  wire [4:0] T_1226;
  wire  T_1227;
  wire  T_1228;
  wire  T_1229;
  wire  T_1230;
  wire  T_1231;
  wire [4:0] T_1239;
  wire [4:0] T_1240;
  wire [4:0] T_1241;
  wire [4:0] T_1242;
  wire [4:0] T_1243;
  wire [1:0] T_1244;
  wire [1:0] T_1245;
  wire [2:0] T_1246;
  wire [4:0] T_1247;
  wire  T_1249;
  wire  T_1251;
  wire [4:0] T_1253;
  wire [4:0] T_1254;
  wire  T_1256;
  wire  T_1257;
  wire  T_1260;
  wire  T_1261;
  wire  T_1262;
  wire  T_1263;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire  T_1271;
  wire  T_1272;
  wire  T_1273;
  wire  T_1276;
  wire  T_1277;
  wire  T_1278;
  wire  T_1281;
  wire  T_1282;
  wire  T_1283;
  wire [1:0] T_1284;
  wire [1:0] T_1285;
  wire [2:0] T_1286;
  wire [4:0] T_1287;
  wire [1:0] T_1288;
  wire [1:0] T_1289;
  wire [2:0] T_1290;
  wire [4:0] T_1291;
  wire  T_1292;
  wire  T_1293;
  wire  T_1294;
  wire  T_1295;
  wire  T_1296;
  wire [4:0] T_1304;
  wire [4:0] T_1305;
  wire [4:0] T_1306;
  wire [4:0] T_1307;
  wire [4:0] T_1308;
  wire [1:0] T_1309;
  wire [1:0] T_1310;
  wire [2:0] T_1311;
  wire [4:0] T_1312;
  wire  T_1314;
  wire  T_1316;
  wire [4:0] T_1319;
  wire [4:0] T_1320;
  wire  T_1322;
  wire  T_1327;
  wire  T_1328;
  wire  T_1332;
  wire  T_1333;
  wire  T_1337;
  wire  T_1338;
  wire  T_1342;
  wire  T_1343;
  wire  T_1347;
  wire  T_1348;
  wire  LockingRRArbiter_7_1_clk;
  wire  LockingRRArbiter_7_1_reset;
  wire  LockingRRArbiter_7_1_io_in_0_ready;
  wire  LockingRRArbiter_7_1_io_in_0_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_0_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_1_ready;
  wire  LockingRRArbiter_7_1_io_in_1_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_1_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_2_ready;
  wire  LockingRRArbiter_7_1_io_in_2_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_2_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_3_ready;
  wire  LockingRRArbiter_7_1_io_in_3_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_3_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_3_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_3_bits_client_id;
  wire  LockingRRArbiter_7_1_io_in_4_ready;
  wire  LockingRRArbiter_7_1_io_in_4_valid;
  wire [25:0] LockingRRArbiter_7_1_io_in_4_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_in_4_bits_p_type;
  wire  LockingRRArbiter_7_1_io_in_4_bits_client_id;
  wire  LockingRRArbiter_7_1_io_out_ready;
  wire  LockingRRArbiter_7_1_io_out_valid;
  wire [25:0] LockingRRArbiter_7_1_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_7_1_io_out_bits_p_type;
  wire  LockingRRArbiter_7_1_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_7_1_io_chosen;
  wire  LockingRRArbiter_8_1_clk;
  wire  LockingRRArbiter_8_1_reset;
  wire  LockingRRArbiter_8_1_io_in_0_ready;
  wire  LockingRRArbiter_8_1_io_in_0_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_0_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_0_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_0_bits_data;
  wire  LockingRRArbiter_8_1_io_in_0_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_1_ready;
  wire  LockingRRArbiter_8_1_io_in_1_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_1_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_1_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_1_bits_data;
  wire  LockingRRArbiter_8_1_io_in_1_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_2_ready;
  wire  LockingRRArbiter_8_1_io_in_2_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_2_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_2_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_2_bits_data;
  wire  LockingRRArbiter_8_1_io_in_2_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_3_ready;
  wire  LockingRRArbiter_8_1_io_in_3_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_3_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_3_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_3_bits_data;
  wire  LockingRRArbiter_8_1_io_in_3_bits_client_id;
  wire  LockingRRArbiter_8_1_io_in_4_ready;
  wire  LockingRRArbiter_8_1_io_in_4_valid;
  wire [2:0] LockingRRArbiter_8_1_io_in_4_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_in_4_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_in_4_bits_data;
  wire  LockingRRArbiter_8_1_io_in_4_bits_client_id;
  wire  LockingRRArbiter_8_1_io_out_ready;
  wire  LockingRRArbiter_8_1_io_out_valid;
  wire [2:0] LockingRRArbiter_8_1_io_out_bits_addr_beat;
  wire [1:0] LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  wire  LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_8_1_io_out_bits_g_type;
  wire [63:0] LockingRRArbiter_8_1_io_out_bits_data;
  wire  LockingRRArbiter_8_1_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_8_1_io_chosen;
  wire  T_1351;
  wire  T_1352;
  wire  T_1354;
  wire  T_1355;
  wire  T_1357;
  wire  T_1358;
  wire  T_1360;
  wire  T_1361;
  wire  T_1363;
  wire  T_1364;
  wire [2:0] T_1366;
  wire  T_1368;
  wire [2:0] T_1370;
  wire  T_1372;
  wire  T_1376;
  wire  T_1377;
  wire  T_1382;
  wire  T_1383;
  wire  T_1384;
  wire  T_1388;
  wire  T_1389;
  wire  T_1391;
  wire  GEN_0;
  reg [31:0] GEN_5;
  wire  GEN_1;
  reg [31:0] GEN_6;
  wire  GEN_2;
  reg [31:0] GEN_7;
  wire  GEN_3;
  reg [31:0] GEN_8;
  wire  GEN_4;
  reg [31:0] GEN_9;
  BufferedBroadcastVoluntaryReleaseTracker trackerList_0 (
    .clk(trackerList_0_clk),
    .reset(trackerList_0_reset),
    .io_inner_acquire_ready(trackerList_0_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_0_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_0_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_0_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_0_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_0_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_0_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_0_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_0_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_0_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_0_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_0_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_0_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_0_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_0_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_0_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_0_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_0_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_0_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_0_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_0_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_0_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_0_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_0_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_0_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_0_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_0_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_0_io_inner_release_ready),
    .io_inner_release_valid(trackerList_0_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_0_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_0_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_0_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_0_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_0_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_0_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_0_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_0_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_0_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_0_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_0_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_0_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_0_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_0_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_0_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_0_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_0_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_0_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_0_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_0_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_0_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_0_io_outer_release_ready),
    .io_outer_release_valid(trackerList_0_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_0_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_0_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_0_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_0_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_0_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_0_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_0_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_0_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_0_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_0_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_0_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_0_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_0_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_0_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_0_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_0_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_0_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_0_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_0_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_0_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_0_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_0_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_0_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_0_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_0_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_0_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_0_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_0_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_0_io_alloc_idle),
    .io_alloc_addr_block(trackerList_0_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker trackerList_1 (
    .clk(trackerList_1_clk),
    .reset(trackerList_1_reset),
    .io_inner_acquire_ready(trackerList_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_1_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_1_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_1_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_1_io_inner_release_ready),
    .io_inner_release_valid(trackerList_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_1_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_1_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_1_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_1_io_outer_release_ready),
    .io_outer_release_valid(trackerList_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_1_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_1_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_1_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_1_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_1_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_1_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_1_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_1_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_1_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_1_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_1_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_1_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_1_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_1_io_alloc_idle),
    .io_alloc_addr_block(trackerList_1_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker_1 trackerList_2 (
    .clk(trackerList_2_clk),
    .reset(trackerList_2_reset),
    .io_inner_acquire_ready(trackerList_2_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_2_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_2_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_2_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_2_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_2_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_2_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_2_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_2_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_2_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_2_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_2_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_2_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_2_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_2_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_2_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_2_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_2_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_2_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_2_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_2_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_2_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_2_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_2_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_2_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_2_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_2_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_2_io_inner_release_ready),
    .io_inner_release_valid(trackerList_2_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_2_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_2_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_2_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_2_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_2_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_2_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_2_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_2_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_2_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_2_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_2_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_2_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_2_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_2_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_2_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_2_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_2_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_2_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_2_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_2_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_2_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_2_io_outer_release_ready),
    .io_outer_release_valid(trackerList_2_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_2_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_2_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_2_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_2_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_2_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_2_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_2_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_2_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_2_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_2_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_2_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_2_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_2_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_2_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_2_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_2_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_2_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_2_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_2_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_2_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_2_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_2_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_2_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_2_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_2_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_2_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_2_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_2_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_2_io_alloc_idle),
    .io_alloc_addr_block(trackerList_2_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker_2 trackerList_3 (
    .clk(trackerList_3_clk),
    .reset(trackerList_3_reset),
    .io_inner_acquire_ready(trackerList_3_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_3_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_3_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_3_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_3_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_3_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_3_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_3_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_3_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_3_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_3_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_3_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_3_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_3_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_3_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_3_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_3_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_3_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_3_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_3_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_3_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_3_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_3_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_3_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_3_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_3_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_3_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_3_io_inner_release_ready),
    .io_inner_release_valid(trackerList_3_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_3_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_3_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_3_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_3_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_3_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_3_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_3_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_3_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_3_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_3_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_3_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_3_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_3_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_3_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_3_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_3_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_3_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_3_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_3_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_3_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_3_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_3_io_outer_release_ready),
    .io_outer_release_valid(trackerList_3_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_3_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_3_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_3_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_3_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_3_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_3_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_3_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_3_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_3_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_3_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_3_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_3_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_3_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_3_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_3_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_3_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_3_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_3_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_3_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_3_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_3_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_3_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_3_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_3_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_3_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_3_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_3_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_3_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_3_io_alloc_idle),
    .io_alloc_addr_block(trackerList_3_io_alloc_addr_block)
  );
  BufferedBroadcastAcquireTracker_3 trackerList_4 (
    .clk(trackerList_4_clk),
    .reset(trackerList_4_reset),
    .io_inner_acquire_ready(trackerList_4_io_inner_acquire_ready),
    .io_inner_acquire_valid(trackerList_4_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(trackerList_4_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(trackerList_4_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(trackerList_4_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(trackerList_4_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(trackerList_4_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(trackerList_4_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(trackerList_4_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(trackerList_4_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(trackerList_4_io_inner_grant_ready),
    .io_inner_grant_valid(trackerList_4_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(trackerList_4_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(trackerList_4_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(trackerList_4_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(trackerList_4_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(trackerList_4_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(trackerList_4_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(trackerList_4_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(trackerList_4_io_inner_finish_ready),
    .io_inner_finish_valid(trackerList_4_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(trackerList_4_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(trackerList_4_io_inner_probe_ready),
    .io_inner_probe_valid(trackerList_4_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(trackerList_4_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(trackerList_4_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(trackerList_4_io_inner_probe_bits_client_id),
    .io_inner_release_ready(trackerList_4_io_inner_release_ready),
    .io_inner_release_valid(trackerList_4_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(trackerList_4_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(trackerList_4_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(trackerList_4_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(trackerList_4_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(trackerList_4_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(trackerList_4_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(trackerList_4_io_inner_release_bits_client_id),
    .io_incoherent_0(trackerList_4_io_incoherent_0),
    .io_outer_acquire_ready(trackerList_4_io_outer_acquire_ready),
    .io_outer_acquire_valid(trackerList_4_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(trackerList_4_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(trackerList_4_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(trackerList_4_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(trackerList_4_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(trackerList_4_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(trackerList_4_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(trackerList_4_io_outer_acquire_bits_data),
    .io_outer_probe_ready(trackerList_4_io_outer_probe_ready),
    .io_outer_probe_valid(trackerList_4_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(trackerList_4_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(trackerList_4_io_outer_probe_bits_p_type),
    .io_outer_release_ready(trackerList_4_io_outer_release_ready),
    .io_outer_release_valid(trackerList_4_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(trackerList_4_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(trackerList_4_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(trackerList_4_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(trackerList_4_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(trackerList_4_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(trackerList_4_io_outer_release_bits_data),
    .io_outer_grant_ready(trackerList_4_io_outer_grant_ready),
    .io_outer_grant_valid(trackerList_4_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(trackerList_4_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(trackerList_4_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(trackerList_4_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(trackerList_4_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(trackerList_4_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(trackerList_4_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(trackerList_4_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(trackerList_4_io_outer_finish_ready),
    .io_outer_finish_valid(trackerList_4_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(trackerList_4_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(trackerList_4_io_outer_finish_bits_manager_id),
    .io_alloc_iacq_matches(trackerList_4_io_alloc_iacq_matches),
    .io_alloc_iacq_can(trackerList_4_io_alloc_iacq_can),
    .io_alloc_iacq_should(trackerList_4_io_alloc_iacq_should),
    .io_alloc_irel_matches(trackerList_4_io_alloc_irel_matches),
    .io_alloc_irel_can(trackerList_4_io_alloc_irel_can),
    .io_alloc_irel_should(trackerList_4_io_alloc_irel_should),
    .io_alloc_oprb_matches(trackerList_4_io_alloc_oprb_matches),
    .io_alloc_oprb_can(trackerList_4_io_alloc_oprb_can),
    .io_alloc_oprb_should(trackerList_4_io_alloc_oprb_should),
    .io_alloc_idle(trackerList_4_io_alloc_idle),
    .io_alloc_addr_block(trackerList_4_io_alloc_addr_block)
  );
  ClientTileLinkIOArbiter outer_arb (
    .clk(outer_arb_clk),
    .reset(outer_arb_reset),
    .io_in_0_acquire_ready(outer_arb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(outer_arb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(outer_arb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(outer_arb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(outer_arb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(outer_arb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(outer_arb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(outer_arb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(outer_arb_io_in_0_acquire_bits_data),
    .io_in_0_probe_ready(outer_arb_io_in_0_probe_ready),
    .io_in_0_probe_valid(outer_arb_io_in_0_probe_valid),
    .io_in_0_probe_bits_addr_block(outer_arb_io_in_0_probe_bits_addr_block),
    .io_in_0_probe_bits_p_type(outer_arb_io_in_0_probe_bits_p_type),
    .io_in_0_release_ready(outer_arb_io_in_0_release_ready),
    .io_in_0_release_valid(outer_arb_io_in_0_release_valid),
    .io_in_0_release_bits_addr_beat(outer_arb_io_in_0_release_bits_addr_beat),
    .io_in_0_release_bits_addr_block(outer_arb_io_in_0_release_bits_addr_block),
    .io_in_0_release_bits_client_xact_id(outer_arb_io_in_0_release_bits_client_xact_id),
    .io_in_0_release_bits_voluntary(outer_arb_io_in_0_release_bits_voluntary),
    .io_in_0_release_bits_r_type(outer_arb_io_in_0_release_bits_r_type),
    .io_in_0_release_bits_data(outer_arb_io_in_0_release_bits_data),
    .io_in_0_grant_ready(outer_arb_io_in_0_grant_ready),
    .io_in_0_grant_valid(outer_arb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(outer_arb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(outer_arb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(outer_arb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(outer_arb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(outer_arb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(outer_arb_io_in_0_grant_bits_data),
    .io_in_0_grant_bits_manager_id(outer_arb_io_in_0_grant_bits_manager_id),
    .io_in_0_finish_ready(outer_arb_io_in_0_finish_ready),
    .io_in_0_finish_valid(outer_arb_io_in_0_finish_valid),
    .io_in_0_finish_bits_manager_xact_id(outer_arb_io_in_0_finish_bits_manager_xact_id),
    .io_in_0_finish_bits_manager_id(outer_arb_io_in_0_finish_bits_manager_id),
    .io_in_1_acquire_ready(outer_arb_io_in_1_acquire_ready),
    .io_in_1_acquire_valid(outer_arb_io_in_1_acquire_valid),
    .io_in_1_acquire_bits_addr_block(outer_arb_io_in_1_acquire_bits_addr_block),
    .io_in_1_acquire_bits_client_xact_id(outer_arb_io_in_1_acquire_bits_client_xact_id),
    .io_in_1_acquire_bits_addr_beat(outer_arb_io_in_1_acquire_bits_addr_beat),
    .io_in_1_acquire_bits_is_builtin_type(outer_arb_io_in_1_acquire_bits_is_builtin_type),
    .io_in_1_acquire_bits_a_type(outer_arb_io_in_1_acquire_bits_a_type),
    .io_in_1_acquire_bits_union(outer_arb_io_in_1_acquire_bits_union),
    .io_in_1_acquire_bits_data(outer_arb_io_in_1_acquire_bits_data),
    .io_in_1_probe_ready(outer_arb_io_in_1_probe_ready),
    .io_in_1_probe_valid(outer_arb_io_in_1_probe_valid),
    .io_in_1_probe_bits_addr_block(outer_arb_io_in_1_probe_bits_addr_block),
    .io_in_1_probe_bits_p_type(outer_arb_io_in_1_probe_bits_p_type),
    .io_in_1_release_ready(outer_arb_io_in_1_release_ready),
    .io_in_1_release_valid(outer_arb_io_in_1_release_valid),
    .io_in_1_release_bits_addr_beat(outer_arb_io_in_1_release_bits_addr_beat),
    .io_in_1_release_bits_addr_block(outer_arb_io_in_1_release_bits_addr_block),
    .io_in_1_release_bits_client_xact_id(outer_arb_io_in_1_release_bits_client_xact_id),
    .io_in_1_release_bits_voluntary(outer_arb_io_in_1_release_bits_voluntary),
    .io_in_1_release_bits_r_type(outer_arb_io_in_1_release_bits_r_type),
    .io_in_1_release_bits_data(outer_arb_io_in_1_release_bits_data),
    .io_in_1_grant_ready(outer_arb_io_in_1_grant_ready),
    .io_in_1_grant_valid(outer_arb_io_in_1_grant_valid),
    .io_in_1_grant_bits_addr_beat(outer_arb_io_in_1_grant_bits_addr_beat),
    .io_in_1_grant_bits_client_xact_id(outer_arb_io_in_1_grant_bits_client_xact_id),
    .io_in_1_grant_bits_manager_xact_id(outer_arb_io_in_1_grant_bits_manager_xact_id),
    .io_in_1_grant_bits_is_builtin_type(outer_arb_io_in_1_grant_bits_is_builtin_type),
    .io_in_1_grant_bits_g_type(outer_arb_io_in_1_grant_bits_g_type),
    .io_in_1_grant_bits_data(outer_arb_io_in_1_grant_bits_data),
    .io_in_1_grant_bits_manager_id(outer_arb_io_in_1_grant_bits_manager_id),
    .io_in_1_finish_ready(outer_arb_io_in_1_finish_ready),
    .io_in_1_finish_valid(outer_arb_io_in_1_finish_valid),
    .io_in_1_finish_bits_manager_xact_id(outer_arb_io_in_1_finish_bits_manager_xact_id),
    .io_in_1_finish_bits_manager_id(outer_arb_io_in_1_finish_bits_manager_id),
    .io_in_2_acquire_ready(outer_arb_io_in_2_acquire_ready),
    .io_in_2_acquire_valid(outer_arb_io_in_2_acquire_valid),
    .io_in_2_acquire_bits_addr_block(outer_arb_io_in_2_acquire_bits_addr_block),
    .io_in_2_acquire_bits_client_xact_id(outer_arb_io_in_2_acquire_bits_client_xact_id),
    .io_in_2_acquire_bits_addr_beat(outer_arb_io_in_2_acquire_bits_addr_beat),
    .io_in_2_acquire_bits_is_builtin_type(outer_arb_io_in_2_acquire_bits_is_builtin_type),
    .io_in_2_acquire_bits_a_type(outer_arb_io_in_2_acquire_bits_a_type),
    .io_in_2_acquire_bits_union(outer_arb_io_in_2_acquire_bits_union),
    .io_in_2_acquire_bits_data(outer_arb_io_in_2_acquire_bits_data),
    .io_in_2_probe_ready(outer_arb_io_in_2_probe_ready),
    .io_in_2_probe_valid(outer_arb_io_in_2_probe_valid),
    .io_in_2_probe_bits_addr_block(outer_arb_io_in_2_probe_bits_addr_block),
    .io_in_2_probe_bits_p_type(outer_arb_io_in_2_probe_bits_p_type),
    .io_in_2_release_ready(outer_arb_io_in_2_release_ready),
    .io_in_2_release_valid(outer_arb_io_in_2_release_valid),
    .io_in_2_release_bits_addr_beat(outer_arb_io_in_2_release_bits_addr_beat),
    .io_in_2_release_bits_addr_block(outer_arb_io_in_2_release_bits_addr_block),
    .io_in_2_release_bits_client_xact_id(outer_arb_io_in_2_release_bits_client_xact_id),
    .io_in_2_release_bits_voluntary(outer_arb_io_in_2_release_bits_voluntary),
    .io_in_2_release_bits_r_type(outer_arb_io_in_2_release_bits_r_type),
    .io_in_2_release_bits_data(outer_arb_io_in_2_release_bits_data),
    .io_in_2_grant_ready(outer_arb_io_in_2_grant_ready),
    .io_in_2_grant_valid(outer_arb_io_in_2_grant_valid),
    .io_in_2_grant_bits_addr_beat(outer_arb_io_in_2_grant_bits_addr_beat),
    .io_in_2_grant_bits_client_xact_id(outer_arb_io_in_2_grant_bits_client_xact_id),
    .io_in_2_grant_bits_manager_xact_id(outer_arb_io_in_2_grant_bits_manager_xact_id),
    .io_in_2_grant_bits_is_builtin_type(outer_arb_io_in_2_grant_bits_is_builtin_type),
    .io_in_2_grant_bits_g_type(outer_arb_io_in_2_grant_bits_g_type),
    .io_in_2_grant_bits_data(outer_arb_io_in_2_grant_bits_data),
    .io_in_2_grant_bits_manager_id(outer_arb_io_in_2_grant_bits_manager_id),
    .io_in_2_finish_ready(outer_arb_io_in_2_finish_ready),
    .io_in_2_finish_valid(outer_arb_io_in_2_finish_valid),
    .io_in_2_finish_bits_manager_xact_id(outer_arb_io_in_2_finish_bits_manager_xact_id),
    .io_in_2_finish_bits_manager_id(outer_arb_io_in_2_finish_bits_manager_id),
    .io_in_3_acquire_ready(outer_arb_io_in_3_acquire_ready),
    .io_in_3_acquire_valid(outer_arb_io_in_3_acquire_valid),
    .io_in_3_acquire_bits_addr_block(outer_arb_io_in_3_acquire_bits_addr_block),
    .io_in_3_acquire_bits_client_xact_id(outer_arb_io_in_3_acquire_bits_client_xact_id),
    .io_in_3_acquire_bits_addr_beat(outer_arb_io_in_3_acquire_bits_addr_beat),
    .io_in_3_acquire_bits_is_builtin_type(outer_arb_io_in_3_acquire_bits_is_builtin_type),
    .io_in_3_acquire_bits_a_type(outer_arb_io_in_3_acquire_bits_a_type),
    .io_in_3_acquire_bits_union(outer_arb_io_in_3_acquire_bits_union),
    .io_in_3_acquire_bits_data(outer_arb_io_in_3_acquire_bits_data),
    .io_in_3_probe_ready(outer_arb_io_in_3_probe_ready),
    .io_in_3_probe_valid(outer_arb_io_in_3_probe_valid),
    .io_in_3_probe_bits_addr_block(outer_arb_io_in_3_probe_bits_addr_block),
    .io_in_3_probe_bits_p_type(outer_arb_io_in_3_probe_bits_p_type),
    .io_in_3_release_ready(outer_arb_io_in_3_release_ready),
    .io_in_3_release_valid(outer_arb_io_in_3_release_valid),
    .io_in_3_release_bits_addr_beat(outer_arb_io_in_3_release_bits_addr_beat),
    .io_in_3_release_bits_addr_block(outer_arb_io_in_3_release_bits_addr_block),
    .io_in_3_release_bits_client_xact_id(outer_arb_io_in_3_release_bits_client_xact_id),
    .io_in_3_release_bits_voluntary(outer_arb_io_in_3_release_bits_voluntary),
    .io_in_3_release_bits_r_type(outer_arb_io_in_3_release_bits_r_type),
    .io_in_3_release_bits_data(outer_arb_io_in_3_release_bits_data),
    .io_in_3_grant_ready(outer_arb_io_in_3_grant_ready),
    .io_in_3_grant_valid(outer_arb_io_in_3_grant_valid),
    .io_in_3_grant_bits_addr_beat(outer_arb_io_in_3_grant_bits_addr_beat),
    .io_in_3_grant_bits_client_xact_id(outer_arb_io_in_3_grant_bits_client_xact_id),
    .io_in_3_grant_bits_manager_xact_id(outer_arb_io_in_3_grant_bits_manager_xact_id),
    .io_in_3_grant_bits_is_builtin_type(outer_arb_io_in_3_grant_bits_is_builtin_type),
    .io_in_3_grant_bits_g_type(outer_arb_io_in_3_grant_bits_g_type),
    .io_in_3_grant_bits_data(outer_arb_io_in_3_grant_bits_data),
    .io_in_3_grant_bits_manager_id(outer_arb_io_in_3_grant_bits_manager_id),
    .io_in_3_finish_ready(outer_arb_io_in_3_finish_ready),
    .io_in_3_finish_valid(outer_arb_io_in_3_finish_valid),
    .io_in_3_finish_bits_manager_xact_id(outer_arb_io_in_3_finish_bits_manager_xact_id),
    .io_in_3_finish_bits_manager_id(outer_arb_io_in_3_finish_bits_manager_id),
    .io_in_4_acquire_ready(outer_arb_io_in_4_acquire_ready),
    .io_in_4_acquire_valid(outer_arb_io_in_4_acquire_valid),
    .io_in_4_acquire_bits_addr_block(outer_arb_io_in_4_acquire_bits_addr_block),
    .io_in_4_acquire_bits_client_xact_id(outer_arb_io_in_4_acquire_bits_client_xact_id),
    .io_in_4_acquire_bits_addr_beat(outer_arb_io_in_4_acquire_bits_addr_beat),
    .io_in_4_acquire_bits_is_builtin_type(outer_arb_io_in_4_acquire_bits_is_builtin_type),
    .io_in_4_acquire_bits_a_type(outer_arb_io_in_4_acquire_bits_a_type),
    .io_in_4_acquire_bits_union(outer_arb_io_in_4_acquire_bits_union),
    .io_in_4_acquire_bits_data(outer_arb_io_in_4_acquire_bits_data),
    .io_in_4_probe_ready(outer_arb_io_in_4_probe_ready),
    .io_in_4_probe_valid(outer_arb_io_in_4_probe_valid),
    .io_in_4_probe_bits_addr_block(outer_arb_io_in_4_probe_bits_addr_block),
    .io_in_4_probe_bits_p_type(outer_arb_io_in_4_probe_bits_p_type),
    .io_in_4_release_ready(outer_arb_io_in_4_release_ready),
    .io_in_4_release_valid(outer_arb_io_in_4_release_valid),
    .io_in_4_release_bits_addr_beat(outer_arb_io_in_4_release_bits_addr_beat),
    .io_in_4_release_bits_addr_block(outer_arb_io_in_4_release_bits_addr_block),
    .io_in_4_release_bits_client_xact_id(outer_arb_io_in_4_release_bits_client_xact_id),
    .io_in_4_release_bits_voluntary(outer_arb_io_in_4_release_bits_voluntary),
    .io_in_4_release_bits_r_type(outer_arb_io_in_4_release_bits_r_type),
    .io_in_4_release_bits_data(outer_arb_io_in_4_release_bits_data),
    .io_in_4_grant_ready(outer_arb_io_in_4_grant_ready),
    .io_in_4_grant_valid(outer_arb_io_in_4_grant_valid),
    .io_in_4_grant_bits_addr_beat(outer_arb_io_in_4_grant_bits_addr_beat),
    .io_in_4_grant_bits_client_xact_id(outer_arb_io_in_4_grant_bits_client_xact_id),
    .io_in_4_grant_bits_manager_xact_id(outer_arb_io_in_4_grant_bits_manager_xact_id),
    .io_in_4_grant_bits_is_builtin_type(outer_arb_io_in_4_grant_bits_is_builtin_type),
    .io_in_4_grant_bits_g_type(outer_arb_io_in_4_grant_bits_g_type),
    .io_in_4_grant_bits_data(outer_arb_io_in_4_grant_bits_data),
    .io_in_4_grant_bits_manager_id(outer_arb_io_in_4_grant_bits_manager_id),
    .io_in_4_finish_ready(outer_arb_io_in_4_finish_ready),
    .io_in_4_finish_valid(outer_arb_io_in_4_finish_valid),
    .io_in_4_finish_bits_manager_xact_id(outer_arb_io_in_4_finish_bits_manager_xact_id),
    .io_in_4_finish_bits_manager_id(outer_arb_io_in_4_finish_bits_manager_id),
    .io_out_acquire_ready(outer_arb_io_out_acquire_ready),
    .io_out_acquire_valid(outer_arb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(outer_arb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(outer_arb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(outer_arb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(outer_arb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(outer_arb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(outer_arb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(outer_arb_io_out_acquire_bits_data),
    .io_out_probe_ready(outer_arb_io_out_probe_ready),
    .io_out_probe_valid(outer_arb_io_out_probe_valid),
    .io_out_probe_bits_addr_block(outer_arb_io_out_probe_bits_addr_block),
    .io_out_probe_bits_p_type(outer_arb_io_out_probe_bits_p_type),
    .io_out_release_ready(outer_arb_io_out_release_ready),
    .io_out_release_valid(outer_arb_io_out_release_valid),
    .io_out_release_bits_addr_beat(outer_arb_io_out_release_bits_addr_beat),
    .io_out_release_bits_addr_block(outer_arb_io_out_release_bits_addr_block),
    .io_out_release_bits_client_xact_id(outer_arb_io_out_release_bits_client_xact_id),
    .io_out_release_bits_voluntary(outer_arb_io_out_release_bits_voluntary),
    .io_out_release_bits_r_type(outer_arb_io_out_release_bits_r_type),
    .io_out_release_bits_data(outer_arb_io_out_release_bits_data),
    .io_out_grant_ready(outer_arb_io_out_grant_ready),
    .io_out_grant_valid(outer_arb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(outer_arb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(outer_arb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(outer_arb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(outer_arb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(outer_arb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(outer_arb_io_out_grant_bits_data),
    .io_out_grant_bits_manager_id(outer_arb_io_out_grant_bits_manager_id),
    .io_out_finish_ready(outer_arb_io_out_finish_ready),
    .io_out_finish_valid(outer_arb_io_out_finish_valid),
    .io_out_finish_bits_manager_xact_id(outer_arb_io_out_finish_bits_manager_xact_id),
    .io_out_finish_bits_manager_id(outer_arb_io_out_finish_bits_manager_id)
  );
  LockingRRArbiter_7 LockingRRArbiter_7_1 (
    .clk(LockingRRArbiter_7_1_clk),
    .reset(LockingRRArbiter_7_1_reset),
    .io_in_0_ready(LockingRRArbiter_7_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_7_1_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_7_1_io_in_0_bits_addr_block),
    .io_in_0_bits_p_type(LockingRRArbiter_7_1_io_in_0_bits_p_type),
    .io_in_0_bits_client_id(LockingRRArbiter_7_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_7_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_7_1_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_7_1_io_in_1_bits_addr_block),
    .io_in_1_bits_p_type(LockingRRArbiter_7_1_io_in_1_bits_p_type),
    .io_in_1_bits_client_id(LockingRRArbiter_7_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_7_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_7_1_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_7_1_io_in_2_bits_addr_block),
    .io_in_2_bits_p_type(LockingRRArbiter_7_1_io_in_2_bits_p_type),
    .io_in_2_bits_client_id(LockingRRArbiter_7_1_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_7_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_7_1_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_7_1_io_in_3_bits_addr_block),
    .io_in_3_bits_p_type(LockingRRArbiter_7_1_io_in_3_bits_p_type),
    .io_in_3_bits_client_id(LockingRRArbiter_7_1_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_7_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_7_1_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_7_1_io_in_4_bits_addr_block),
    .io_in_4_bits_p_type(LockingRRArbiter_7_1_io_in_4_bits_p_type),
    .io_in_4_bits_client_id(LockingRRArbiter_7_1_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_7_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_7_1_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_7_1_io_out_bits_addr_block),
    .io_out_bits_p_type(LockingRRArbiter_7_1_io_out_bits_p_type),
    .io_out_bits_client_id(LockingRRArbiter_7_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_7_1_io_chosen)
  );
  LockingRRArbiter_8 LockingRRArbiter_8_1 (
    .clk(LockingRRArbiter_8_1_clk),
    .reset(LockingRRArbiter_8_1_reset),
    .io_in_0_ready(LockingRRArbiter_8_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_8_1_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_8_1_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_8_1_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(LockingRRArbiter_8_1_io_in_0_bits_g_type),
    .io_in_0_bits_data(LockingRRArbiter_8_1_io_in_0_bits_data),
    .io_in_0_bits_client_id(LockingRRArbiter_8_1_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_8_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_8_1_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_8_1_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_8_1_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(LockingRRArbiter_8_1_io_in_1_bits_g_type),
    .io_in_1_bits_data(LockingRRArbiter_8_1_io_in_1_bits_data),
    .io_in_1_bits_client_id(LockingRRArbiter_8_1_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_8_1_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_8_1_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_8_1_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_8_1_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(LockingRRArbiter_8_1_io_in_2_bits_g_type),
    .io_in_2_bits_data(LockingRRArbiter_8_1_io_in_2_bits_data),
    .io_in_2_bits_client_id(LockingRRArbiter_8_1_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_8_1_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_8_1_io_in_3_valid),
    .io_in_3_bits_addr_beat(LockingRRArbiter_8_1_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_8_1_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(LockingRRArbiter_8_1_io_in_3_bits_g_type),
    .io_in_3_bits_data(LockingRRArbiter_8_1_io_in_3_bits_data),
    .io_in_3_bits_client_id(LockingRRArbiter_8_1_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_8_1_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_8_1_io_in_4_valid),
    .io_in_4_bits_addr_beat(LockingRRArbiter_8_1_io_in_4_bits_addr_beat),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_8_1_io_in_4_bits_client_xact_id),
    .io_in_4_bits_manager_xact_id(LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_g_type(LockingRRArbiter_8_1_io_in_4_bits_g_type),
    .io_in_4_bits_data(LockingRRArbiter_8_1_io_in_4_bits_data),
    .io_in_4_bits_client_id(LockingRRArbiter_8_1_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_8_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_8_1_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_8_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(LockingRRArbiter_8_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(LockingRRArbiter_8_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(LockingRRArbiter_8_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(LockingRRArbiter_8_1_io_out_bits_g_type),
    .io_out_bits_data(LockingRRArbiter_8_1_io_out_bits_data),
    .io_out_bits_client_id(LockingRRArbiter_8_1_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_8_1_io_chosen)
  );
  assign io_inner_acquire_ready = T_1257;
  assign io_inner_grant_valid = LockingRRArbiter_8_1_io_out_valid;
  assign io_inner_grant_bits_addr_beat = LockingRRArbiter_8_1_io_out_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_8_1_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_8_1_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_8_1_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_8_1_io_out_bits_g_type;
  assign io_inner_grant_bits_data = LockingRRArbiter_8_1_io_out_bits_data;
  assign io_inner_grant_bits_client_id = LockingRRArbiter_8_1_io_out_bits_client_id;
  assign io_inner_finish_ready = T_1384;
  assign io_inner_probe_valid = LockingRRArbiter_7_1_io_out_valid;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_7_1_io_out_bits_addr_block;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_7_1_io_out_bits_p_type;
  assign io_inner_probe_bits_client_id = LockingRRArbiter_7_1_io_out_bits_client_id;
  assign io_inner_release_ready = T_1322;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_data = outer_arb_io_out_acquire_bits_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = outer_arb_io_out_release_valid;
  assign io_outer_release_bits_addr_beat = outer_arb_io_out_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = outer_arb_io_out_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = outer_arb_io_out_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = outer_arb_io_out_release_bits_voluntary;
  assign io_outer_release_bits_r_type = outer_arb_io_out_release_bits_r_type;
  assign io_outer_release_bits_data = outer_arb_io_out_release_bits_data;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = outer_arb_io_out_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = outer_arb_io_out_finish_bits_manager_id;
  assign trackerList_0_clk = clk;
  assign trackerList_0_reset = reset;
  assign trackerList_0_io_inner_acquire_valid = T_1260;
  assign trackerList_0_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_0_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_0_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_0_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_0_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_0_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_0_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_0_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_0_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_0_ready;
  assign trackerList_0_io_inner_finish_valid = T_1352;
  assign trackerList_0_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_0_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_0_ready;
  assign trackerList_0_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_0_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_0_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_0_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_0_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_0_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_0_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_0_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_0_io_incoherent_0 = io_incoherent_0;
  assign trackerList_0_io_outer_acquire_ready = outer_arb_io_in_0_acquire_ready;
  assign trackerList_0_io_outer_probe_valid = outer_arb_io_in_0_probe_valid;
  assign trackerList_0_io_outer_probe_bits_addr_block = outer_arb_io_in_0_probe_bits_addr_block;
  assign trackerList_0_io_outer_probe_bits_p_type = outer_arb_io_in_0_probe_bits_p_type;
  assign trackerList_0_io_outer_release_ready = outer_arb_io_in_0_release_ready;
  assign trackerList_0_io_outer_grant_valid = outer_arb_io_in_0_grant_valid;
  assign trackerList_0_io_outer_grant_bits_addr_beat = outer_arb_io_in_0_grant_bits_addr_beat;
  assign trackerList_0_io_outer_grant_bits_client_xact_id = outer_arb_io_in_0_grant_bits_client_xact_id;
  assign trackerList_0_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_0_grant_bits_manager_xact_id;
  assign trackerList_0_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_0_grant_bits_is_builtin_type;
  assign trackerList_0_io_outer_grant_bits_g_type = outer_arb_io_in_0_grant_bits_g_type;
  assign trackerList_0_io_outer_grant_bits_data = outer_arb_io_in_0_grant_bits_data;
  assign trackerList_0_io_outer_grant_bits_manager_id = outer_arb_io_in_0_grant_bits_manager_id;
  assign trackerList_0_io_outer_finish_ready = outer_arb_io_in_0_finish_ready;
  assign trackerList_0_io_alloc_iacq_should = T_1263;
  assign trackerList_0_io_alloc_irel_should = T_1328;
  assign trackerList_0_io_alloc_oprb_should = GEN_0;
  assign trackerList_1_clk = clk;
  assign trackerList_1_reset = reset;
  assign trackerList_1_io_inner_acquire_valid = T_1260;
  assign trackerList_1_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_1_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_1_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_1_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_1_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_1_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_1_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_1_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_1_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_1_ready;
  assign trackerList_1_io_inner_finish_valid = T_1355;
  assign trackerList_1_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_1_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_1_ready;
  assign trackerList_1_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_1_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_1_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_1_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_1_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_1_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_1_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_1_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_1_io_incoherent_0 = io_incoherent_0;
  assign trackerList_1_io_outer_acquire_ready = outer_arb_io_in_1_acquire_ready;
  assign trackerList_1_io_outer_probe_valid = outer_arb_io_in_1_probe_valid;
  assign trackerList_1_io_outer_probe_bits_addr_block = outer_arb_io_in_1_probe_bits_addr_block;
  assign trackerList_1_io_outer_probe_bits_p_type = outer_arb_io_in_1_probe_bits_p_type;
  assign trackerList_1_io_outer_release_ready = outer_arb_io_in_1_release_ready;
  assign trackerList_1_io_outer_grant_valid = outer_arb_io_in_1_grant_valid;
  assign trackerList_1_io_outer_grant_bits_addr_beat = outer_arb_io_in_1_grant_bits_addr_beat;
  assign trackerList_1_io_outer_grant_bits_client_xact_id = outer_arb_io_in_1_grant_bits_client_xact_id;
  assign trackerList_1_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_1_grant_bits_manager_xact_id;
  assign trackerList_1_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_1_grant_bits_is_builtin_type;
  assign trackerList_1_io_outer_grant_bits_g_type = outer_arb_io_in_1_grant_bits_g_type;
  assign trackerList_1_io_outer_grant_bits_data = outer_arb_io_in_1_grant_bits_data;
  assign trackerList_1_io_outer_grant_bits_manager_id = outer_arb_io_in_1_grant_bits_manager_id;
  assign trackerList_1_io_outer_finish_ready = outer_arb_io_in_1_finish_ready;
  assign trackerList_1_io_alloc_iacq_should = T_1268;
  assign trackerList_1_io_alloc_irel_should = T_1333;
  assign trackerList_1_io_alloc_oprb_should = GEN_1;
  assign trackerList_2_clk = clk;
  assign trackerList_2_reset = reset;
  assign trackerList_2_io_inner_acquire_valid = T_1260;
  assign trackerList_2_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_2_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_2_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_2_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_2_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_2_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_2_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_2_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_2_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_2_ready;
  assign trackerList_2_io_inner_finish_valid = T_1358;
  assign trackerList_2_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_2_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_2_ready;
  assign trackerList_2_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_2_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_2_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_2_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_2_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_2_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_2_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_2_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_2_io_incoherent_0 = io_incoherent_0;
  assign trackerList_2_io_outer_acquire_ready = outer_arb_io_in_2_acquire_ready;
  assign trackerList_2_io_outer_probe_valid = outer_arb_io_in_2_probe_valid;
  assign trackerList_2_io_outer_probe_bits_addr_block = outer_arb_io_in_2_probe_bits_addr_block;
  assign trackerList_2_io_outer_probe_bits_p_type = outer_arb_io_in_2_probe_bits_p_type;
  assign trackerList_2_io_outer_release_ready = outer_arb_io_in_2_release_ready;
  assign trackerList_2_io_outer_grant_valid = outer_arb_io_in_2_grant_valid;
  assign trackerList_2_io_outer_grant_bits_addr_beat = outer_arb_io_in_2_grant_bits_addr_beat;
  assign trackerList_2_io_outer_grant_bits_client_xact_id = outer_arb_io_in_2_grant_bits_client_xact_id;
  assign trackerList_2_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_2_grant_bits_manager_xact_id;
  assign trackerList_2_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_2_grant_bits_is_builtin_type;
  assign trackerList_2_io_outer_grant_bits_g_type = outer_arb_io_in_2_grant_bits_g_type;
  assign trackerList_2_io_outer_grant_bits_data = outer_arb_io_in_2_grant_bits_data;
  assign trackerList_2_io_outer_grant_bits_manager_id = outer_arb_io_in_2_grant_bits_manager_id;
  assign trackerList_2_io_outer_finish_ready = outer_arb_io_in_2_finish_ready;
  assign trackerList_2_io_alloc_iacq_should = T_1273;
  assign trackerList_2_io_alloc_irel_should = T_1338;
  assign trackerList_2_io_alloc_oprb_should = GEN_2;
  assign trackerList_3_clk = clk;
  assign trackerList_3_reset = reset;
  assign trackerList_3_io_inner_acquire_valid = T_1260;
  assign trackerList_3_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_3_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_3_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_3_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_3_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_3_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_3_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_3_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_3_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_3_ready;
  assign trackerList_3_io_inner_finish_valid = T_1361;
  assign trackerList_3_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_3_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_3_ready;
  assign trackerList_3_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_3_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_3_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_3_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_3_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_3_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_3_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_3_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_3_io_incoherent_0 = io_incoherent_0;
  assign trackerList_3_io_outer_acquire_ready = outer_arb_io_in_3_acquire_ready;
  assign trackerList_3_io_outer_probe_valid = outer_arb_io_in_3_probe_valid;
  assign trackerList_3_io_outer_probe_bits_addr_block = outer_arb_io_in_3_probe_bits_addr_block;
  assign trackerList_3_io_outer_probe_bits_p_type = outer_arb_io_in_3_probe_bits_p_type;
  assign trackerList_3_io_outer_release_ready = outer_arb_io_in_3_release_ready;
  assign trackerList_3_io_outer_grant_valid = outer_arb_io_in_3_grant_valid;
  assign trackerList_3_io_outer_grant_bits_addr_beat = outer_arb_io_in_3_grant_bits_addr_beat;
  assign trackerList_3_io_outer_grant_bits_client_xact_id = outer_arb_io_in_3_grant_bits_client_xact_id;
  assign trackerList_3_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_3_grant_bits_manager_xact_id;
  assign trackerList_3_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_3_grant_bits_is_builtin_type;
  assign trackerList_3_io_outer_grant_bits_g_type = outer_arb_io_in_3_grant_bits_g_type;
  assign trackerList_3_io_outer_grant_bits_data = outer_arb_io_in_3_grant_bits_data;
  assign trackerList_3_io_outer_grant_bits_manager_id = outer_arb_io_in_3_grant_bits_manager_id;
  assign trackerList_3_io_outer_finish_ready = outer_arb_io_in_3_finish_ready;
  assign trackerList_3_io_alloc_iacq_should = T_1278;
  assign trackerList_3_io_alloc_irel_should = T_1343;
  assign trackerList_3_io_alloc_oprb_should = GEN_3;
  assign trackerList_4_clk = clk;
  assign trackerList_4_reset = reset;
  assign trackerList_4_io_inner_acquire_valid = T_1260;
  assign trackerList_4_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign trackerList_4_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign trackerList_4_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign trackerList_4_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign trackerList_4_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign trackerList_4_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign trackerList_4_io_inner_acquire_bits_data = io_inner_acquire_bits_data;
  assign trackerList_4_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign trackerList_4_io_inner_grant_ready = LockingRRArbiter_8_1_io_in_4_ready;
  assign trackerList_4_io_inner_finish_valid = T_1364;
  assign trackerList_4_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign trackerList_4_io_inner_probe_ready = LockingRRArbiter_7_1_io_in_4_ready;
  assign trackerList_4_io_inner_release_valid = io_inner_release_valid;
  assign trackerList_4_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign trackerList_4_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign trackerList_4_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign trackerList_4_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign trackerList_4_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign trackerList_4_io_inner_release_bits_data = io_inner_release_bits_data;
  assign trackerList_4_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign trackerList_4_io_incoherent_0 = io_incoherent_0;
  assign trackerList_4_io_outer_acquire_ready = outer_arb_io_in_4_acquire_ready;
  assign trackerList_4_io_outer_probe_valid = outer_arb_io_in_4_probe_valid;
  assign trackerList_4_io_outer_probe_bits_addr_block = outer_arb_io_in_4_probe_bits_addr_block;
  assign trackerList_4_io_outer_probe_bits_p_type = outer_arb_io_in_4_probe_bits_p_type;
  assign trackerList_4_io_outer_release_ready = outer_arb_io_in_4_release_ready;
  assign trackerList_4_io_outer_grant_valid = outer_arb_io_in_4_grant_valid;
  assign trackerList_4_io_outer_grant_bits_addr_beat = outer_arb_io_in_4_grant_bits_addr_beat;
  assign trackerList_4_io_outer_grant_bits_client_xact_id = outer_arb_io_in_4_grant_bits_client_xact_id;
  assign trackerList_4_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_4_grant_bits_manager_xact_id;
  assign trackerList_4_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_4_grant_bits_is_builtin_type;
  assign trackerList_4_io_outer_grant_bits_g_type = outer_arb_io_in_4_grant_bits_g_type;
  assign trackerList_4_io_outer_grant_bits_data = outer_arb_io_in_4_grant_bits_data;
  assign trackerList_4_io_outer_grant_bits_manager_id = outer_arb_io_in_4_grant_bits_manager_id;
  assign trackerList_4_io_outer_finish_ready = outer_arb_io_in_4_finish_ready;
  assign trackerList_4_io_alloc_iacq_should = T_1283;
  assign trackerList_4_io_alloc_irel_should = T_1348;
  assign trackerList_4_io_alloc_oprb_should = GEN_4;
  assign outer_arb_clk = clk;
  assign outer_arb_reset = reset;
  assign outer_arb_io_in_0_acquire_valid = trackerList_0_io_outer_acquire_valid;
  assign outer_arb_io_in_0_acquire_bits_addr_block = trackerList_0_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_0_acquire_bits_client_xact_id = trackerList_0_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_0_acquire_bits_addr_beat = trackerList_0_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_0_acquire_bits_is_builtin_type = trackerList_0_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_0_acquire_bits_a_type = trackerList_0_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_0_acquire_bits_union = trackerList_0_io_outer_acquire_bits_union;
  assign outer_arb_io_in_0_acquire_bits_data = trackerList_0_io_outer_acquire_bits_data;
  assign outer_arb_io_in_0_probe_ready = trackerList_0_io_outer_probe_ready;
  assign outer_arb_io_in_0_release_valid = trackerList_0_io_outer_release_valid;
  assign outer_arb_io_in_0_release_bits_addr_beat = trackerList_0_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_0_release_bits_addr_block = trackerList_0_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_0_release_bits_client_xact_id = trackerList_0_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_0_release_bits_voluntary = trackerList_0_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_0_release_bits_r_type = trackerList_0_io_outer_release_bits_r_type;
  assign outer_arb_io_in_0_release_bits_data = trackerList_0_io_outer_release_bits_data;
  assign outer_arb_io_in_0_grant_ready = trackerList_0_io_outer_grant_ready;
  assign outer_arb_io_in_0_finish_valid = trackerList_0_io_outer_finish_valid;
  assign outer_arb_io_in_0_finish_bits_manager_xact_id = trackerList_0_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_0_finish_bits_manager_id = trackerList_0_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_1_acquire_valid = trackerList_1_io_outer_acquire_valid;
  assign outer_arb_io_in_1_acquire_bits_addr_block = trackerList_1_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_1_acquire_bits_client_xact_id = trackerList_1_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_1_acquire_bits_addr_beat = trackerList_1_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_1_acquire_bits_is_builtin_type = trackerList_1_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_1_acquire_bits_a_type = trackerList_1_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_1_acquire_bits_union = trackerList_1_io_outer_acquire_bits_union;
  assign outer_arb_io_in_1_acquire_bits_data = trackerList_1_io_outer_acquire_bits_data;
  assign outer_arb_io_in_1_probe_ready = trackerList_1_io_outer_probe_ready;
  assign outer_arb_io_in_1_release_valid = trackerList_1_io_outer_release_valid;
  assign outer_arb_io_in_1_release_bits_addr_beat = trackerList_1_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_1_release_bits_addr_block = trackerList_1_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_1_release_bits_client_xact_id = trackerList_1_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_1_release_bits_voluntary = trackerList_1_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_1_release_bits_r_type = trackerList_1_io_outer_release_bits_r_type;
  assign outer_arb_io_in_1_release_bits_data = trackerList_1_io_outer_release_bits_data;
  assign outer_arb_io_in_1_grant_ready = trackerList_1_io_outer_grant_ready;
  assign outer_arb_io_in_1_finish_valid = trackerList_1_io_outer_finish_valid;
  assign outer_arb_io_in_1_finish_bits_manager_xact_id = trackerList_1_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_1_finish_bits_manager_id = trackerList_1_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_2_acquire_valid = trackerList_2_io_outer_acquire_valid;
  assign outer_arb_io_in_2_acquire_bits_addr_block = trackerList_2_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_2_acquire_bits_client_xact_id = trackerList_2_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_2_acquire_bits_addr_beat = trackerList_2_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_2_acquire_bits_is_builtin_type = trackerList_2_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_2_acquire_bits_a_type = trackerList_2_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_2_acquire_bits_union = trackerList_2_io_outer_acquire_bits_union;
  assign outer_arb_io_in_2_acquire_bits_data = trackerList_2_io_outer_acquire_bits_data;
  assign outer_arb_io_in_2_probe_ready = trackerList_2_io_outer_probe_ready;
  assign outer_arb_io_in_2_release_valid = trackerList_2_io_outer_release_valid;
  assign outer_arb_io_in_2_release_bits_addr_beat = trackerList_2_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_2_release_bits_addr_block = trackerList_2_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_2_release_bits_client_xact_id = trackerList_2_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_2_release_bits_voluntary = trackerList_2_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_2_release_bits_r_type = trackerList_2_io_outer_release_bits_r_type;
  assign outer_arb_io_in_2_release_bits_data = trackerList_2_io_outer_release_bits_data;
  assign outer_arb_io_in_2_grant_ready = trackerList_2_io_outer_grant_ready;
  assign outer_arb_io_in_2_finish_valid = trackerList_2_io_outer_finish_valid;
  assign outer_arb_io_in_2_finish_bits_manager_xact_id = trackerList_2_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_2_finish_bits_manager_id = trackerList_2_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_3_acquire_valid = trackerList_3_io_outer_acquire_valid;
  assign outer_arb_io_in_3_acquire_bits_addr_block = trackerList_3_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_3_acquire_bits_client_xact_id = trackerList_3_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_3_acquire_bits_addr_beat = trackerList_3_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_3_acquire_bits_is_builtin_type = trackerList_3_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_3_acquire_bits_a_type = trackerList_3_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_3_acquire_bits_union = trackerList_3_io_outer_acquire_bits_union;
  assign outer_arb_io_in_3_acquire_bits_data = trackerList_3_io_outer_acquire_bits_data;
  assign outer_arb_io_in_3_probe_ready = trackerList_3_io_outer_probe_ready;
  assign outer_arb_io_in_3_release_valid = trackerList_3_io_outer_release_valid;
  assign outer_arb_io_in_3_release_bits_addr_beat = trackerList_3_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_3_release_bits_addr_block = trackerList_3_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_3_release_bits_client_xact_id = trackerList_3_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_3_release_bits_voluntary = trackerList_3_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_3_release_bits_r_type = trackerList_3_io_outer_release_bits_r_type;
  assign outer_arb_io_in_3_release_bits_data = trackerList_3_io_outer_release_bits_data;
  assign outer_arb_io_in_3_grant_ready = trackerList_3_io_outer_grant_ready;
  assign outer_arb_io_in_3_finish_valid = trackerList_3_io_outer_finish_valid;
  assign outer_arb_io_in_3_finish_bits_manager_xact_id = trackerList_3_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_3_finish_bits_manager_id = trackerList_3_io_outer_finish_bits_manager_id;
  assign outer_arb_io_in_4_acquire_valid = trackerList_4_io_outer_acquire_valid;
  assign outer_arb_io_in_4_acquire_bits_addr_block = trackerList_4_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_4_acquire_bits_client_xact_id = trackerList_4_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_4_acquire_bits_addr_beat = trackerList_4_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_4_acquire_bits_is_builtin_type = trackerList_4_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_4_acquire_bits_a_type = trackerList_4_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_4_acquire_bits_union = trackerList_4_io_outer_acquire_bits_union;
  assign outer_arb_io_in_4_acquire_bits_data = trackerList_4_io_outer_acquire_bits_data;
  assign outer_arb_io_in_4_probe_ready = trackerList_4_io_outer_probe_ready;
  assign outer_arb_io_in_4_release_valid = trackerList_4_io_outer_release_valid;
  assign outer_arb_io_in_4_release_bits_addr_beat = trackerList_4_io_outer_release_bits_addr_beat;
  assign outer_arb_io_in_4_release_bits_addr_block = trackerList_4_io_outer_release_bits_addr_block;
  assign outer_arb_io_in_4_release_bits_client_xact_id = trackerList_4_io_outer_release_bits_client_xact_id;
  assign outer_arb_io_in_4_release_bits_voluntary = trackerList_4_io_outer_release_bits_voluntary;
  assign outer_arb_io_in_4_release_bits_r_type = trackerList_4_io_outer_release_bits_r_type;
  assign outer_arb_io_in_4_release_bits_data = trackerList_4_io_outer_release_bits_data;
  assign outer_arb_io_in_4_grant_ready = trackerList_4_io_outer_grant_ready;
  assign outer_arb_io_in_4_finish_valid = trackerList_4_io_outer_finish_valid;
  assign outer_arb_io_in_4_finish_bits_manager_xact_id = trackerList_4_io_outer_finish_bits_manager_xact_id;
  assign outer_arb_io_in_4_finish_bits_manager_id = trackerList_4_io_outer_finish_bits_manager_id;
  assign outer_arb_io_out_acquire_ready = io_outer_acquire_ready;
  assign outer_arb_io_out_probe_valid = io_outer_probe_valid;
  assign outer_arb_io_out_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign outer_arb_io_out_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign outer_arb_io_out_release_ready = io_outer_release_ready;
  assign outer_arb_io_out_grant_valid = io_outer_grant_valid;
  assign outer_arb_io_out_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign outer_arb_io_out_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign outer_arb_io_out_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign outer_arb_io_out_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign outer_arb_io_out_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign outer_arb_io_out_grant_bits_data = io_outer_grant_bits_data;
  assign outer_arb_io_out_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign outer_arb_io_out_finish_ready = io_outer_finish_ready;
  assign T_1215 = io_inner_acquire_valid & io_inner_release_valid;
  assign T_1216 = io_inner_release_bits_addr_block == io_inner_acquire_bits_addr_block;
  assign irel_vs_iacq_conflict = T_1215 & T_1216;
  assign T_1218 = irel_vs_iacq_conflict == 1'h0;
  assign T_1219 = {trackerList_1_io_inner_acquire_ready,trackerList_0_io_inner_acquire_ready};
  assign T_1220 = {trackerList_4_io_inner_acquire_ready,trackerList_3_io_inner_acquire_ready};
  assign T_1221 = {T_1220,trackerList_2_io_inner_acquire_ready};
  assign T_1222 = {T_1221,T_1219};
  assign T_1223 = {trackerList_1_io_alloc_iacq_can,trackerList_0_io_alloc_iacq_can};
  assign T_1224 = {trackerList_4_io_alloc_iacq_can,trackerList_3_io_alloc_iacq_can};
  assign T_1225 = {T_1224,trackerList_2_io_alloc_iacq_can};
  assign T_1226 = {T_1225,T_1223};
  assign T_1227 = T_1226[0];
  assign T_1228 = T_1226[1];
  assign T_1229 = T_1226[2];
  assign T_1230 = T_1226[3];
  assign T_1231 = T_1226[4];
  assign T_1239 = T_1231 ? 5'h10 : 5'h0;
  assign T_1240 = T_1230 ? 5'h8 : T_1239;
  assign T_1241 = T_1229 ? 5'h4 : T_1240;
  assign T_1242 = T_1228 ? 5'h2 : T_1241;
  assign T_1243 = T_1227 ? 5'h1 : T_1242;
  assign T_1244 = {trackerList_1_io_alloc_iacq_matches,trackerList_0_io_alloc_iacq_matches};
  assign T_1245 = {trackerList_4_io_alloc_iacq_matches,trackerList_3_io_alloc_iacq_matches};
  assign T_1246 = {T_1245,trackerList_2_io_alloc_iacq_matches};
  assign T_1247 = {T_1246,T_1244};
  assign T_1249 = T_1247 != 5'h0;
  assign T_1251 = T_1249 == 1'h0;
  assign T_1253 = T_1251 ? T_1226 : T_1247;
  assign T_1254 = T_1253 & T_1222;
  assign T_1256 = T_1254 != 5'h0;
  assign T_1257 = T_1256 & T_1218;
  assign T_1260 = io_inner_acquire_valid & T_1218;
  assign T_1261 = T_1243[0];
  assign T_1262 = T_1261 & T_1251;
  assign T_1263 = T_1262 & T_1218;
  assign T_1266 = T_1243[1];
  assign T_1267 = T_1266 & T_1251;
  assign T_1268 = T_1267 & T_1218;
  assign T_1271 = T_1243[2];
  assign T_1272 = T_1271 & T_1251;
  assign T_1273 = T_1272 & T_1218;
  assign T_1276 = T_1243[3];
  assign T_1277 = T_1276 & T_1251;
  assign T_1278 = T_1277 & T_1218;
  assign T_1281 = T_1243[4];
  assign T_1282 = T_1281 & T_1251;
  assign T_1283 = T_1282 & T_1218;
  assign T_1284 = {trackerList_1_io_inner_release_ready,trackerList_0_io_inner_release_ready};
  assign T_1285 = {trackerList_4_io_inner_release_ready,trackerList_3_io_inner_release_ready};
  assign T_1286 = {T_1285,trackerList_2_io_inner_release_ready};
  assign T_1287 = {T_1286,T_1284};
  assign T_1288 = {trackerList_1_io_alloc_irel_can,trackerList_0_io_alloc_irel_can};
  assign T_1289 = {trackerList_4_io_alloc_irel_can,trackerList_3_io_alloc_irel_can};
  assign T_1290 = {T_1289,trackerList_2_io_alloc_irel_can};
  assign T_1291 = {T_1290,T_1288};
  assign T_1292 = T_1291[0];
  assign T_1293 = T_1291[1];
  assign T_1294 = T_1291[2];
  assign T_1295 = T_1291[3];
  assign T_1296 = T_1291[4];
  assign T_1304 = T_1296 ? 5'h10 : 5'h0;
  assign T_1305 = T_1295 ? 5'h8 : T_1304;
  assign T_1306 = T_1294 ? 5'h4 : T_1305;
  assign T_1307 = T_1293 ? 5'h2 : T_1306;
  assign T_1308 = T_1292 ? 5'h1 : T_1307;
  assign T_1309 = {trackerList_1_io_alloc_irel_matches,trackerList_0_io_alloc_irel_matches};
  assign T_1310 = {trackerList_4_io_alloc_irel_matches,trackerList_3_io_alloc_irel_matches};
  assign T_1311 = {T_1310,trackerList_2_io_alloc_irel_matches};
  assign T_1312 = {T_1311,T_1309};
  assign T_1314 = T_1312 != 5'h0;
  assign T_1316 = T_1314 == 1'h0;
  assign T_1319 = T_1316 ? T_1291 : T_1312;
  assign T_1320 = T_1319 & T_1287;
  assign T_1322 = T_1320 != 5'h0;
  assign T_1327 = T_1308[0];
  assign T_1328 = T_1327 & T_1316;
  assign T_1332 = T_1308[1];
  assign T_1333 = T_1332 & T_1316;
  assign T_1337 = T_1308[2];
  assign T_1338 = T_1337 & T_1316;
  assign T_1342 = T_1308[3];
  assign T_1343 = T_1342 & T_1316;
  assign T_1347 = T_1308[4];
  assign T_1348 = T_1347 & T_1316;
  assign LockingRRArbiter_7_1_clk = clk;
  assign LockingRRArbiter_7_1_reset = reset;
  assign LockingRRArbiter_7_1_io_in_0_valid = trackerList_0_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_0_bits_addr_block = trackerList_0_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_0_bits_p_type = trackerList_0_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_0_bits_client_id = trackerList_0_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_1_valid = trackerList_1_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_1_bits_addr_block = trackerList_1_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_1_bits_p_type = trackerList_1_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_1_bits_client_id = trackerList_1_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_2_valid = trackerList_2_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_2_bits_addr_block = trackerList_2_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_2_bits_p_type = trackerList_2_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_2_bits_client_id = trackerList_2_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_3_valid = trackerList_3_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_3_bits_addr_block = trackerList_3_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_3_bits_p_type = trackerList_3_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_3_bits_client_id = trackerList_3_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_in_4_valid = trackerList_4_io_inner_probe_valid;
  assign LockingRRArbiter_7_1_io_in_4_bits_addr_block = trackerList_4_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_7_1_io_in_4_bits_p_type = trackerList_4_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_7_1_io_in_4_bits_client_id = trackerList_4_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_7_1_io_out_ready = io_inner_probe_ready;
  assign LockingRRArbiter_8_1_clk = clk;
  assign LockingRRArbiter_8_1_reset = reset;
  assign LockingRRArbiter_8_1_io_in_0_valid = trackerList_0_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_0_bits_addr_beat = trackerList_0_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_xact_id = trackerList_0_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_manager_xact_id = trackerList_0_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_0_bits_is_builtin_type = trackerList_0_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_g_type = trackerList_0_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_0_bits_data = trackerList_0_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_0_bits_client_id = trackerList_0_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_1_valid = trackerList_1_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_1_bits_addr_beat = trackerList_1_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_xact_id = trackerList_1_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_manager_xact_id = trackerList_1_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_1_bits_is_builtin_type = trackerList_1_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_g_type = trackerList_1_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_1_bits_data = trackerList_1_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_1_bits_client_id = trackerList_1_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_2_valid = trackerList_2_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_2_bits_addr_beat = trackerList_2_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_xact_id = trackerList_2_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_manager_xact_id = trackerList_2_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_2_bits_is_builtin_type = trackerList_2_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_g_type = trackerList_2_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_2_bits_data = trackerList_2_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_2_bits_client_id = trackerList_2_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_3_valid = trackerList_3_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_3_bits_addr_beat = trackerList_3_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_3_bits_client_xact_id = trackerList_3_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_3_bits_manager_xact_id = trackerList_3_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_3_bits_is_builtin_type = trackerList_3_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_3_bits_g_type = trackerList_3_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_3_bits_data = trackerList_3_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_3_bits_client_id = trackerList_3_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_in_4_valid = trackerList_4_io_inner_grant_valid;
  assign LockingRRArbiter_8_1_io_in_4_bits_addr_beat = trackerList_4_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_8_1_io_in_4_bits_client_xact_id = trackerList_4_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_8_1_io_in_4_bits_manager_xact_id = trackerList_4_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_8_1_io_in_4_bits_is_builtin_type = trackerList_4_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_8_1_io_in_4_bits_g_type = trackerList_4_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_8_1_io_in_4_bits_data = trackerList_4_io_inner_grant_bits_data;
  assign LockingRRArbiter_8_1_io_in_4_bits_client_id = trackerList_4_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_8_1_io_out_ready = io_inner_grant_ready;
  assign T_1351 = io_inner_finish_bits_manager_xact_id == 3'h0;
  assign T_1352 = io_inner_finish_valid & T_1351;
  assign T_1354 = io_inner_finish_bits_manager_xact_id == 3'h1;
  assign T_1355 = io_inner_finish_valid & T_1354;
  assign T_1357 = io_inner_finish_bits_manager_xact_id == 3'h2;
  assign T_1358 = io_inner_finish_valid & T_1357;
  assign T_1360 = io_inner_finish_bits_manager_xact_id == 3'h3;
  assign T_1361 = io_inner_finish_valid & T_1360;
  assign T_1363 = io_inner_finish_bits_manager_xact_id == 3'h4;
  assign T_1364 = io_inner_finish_valid & T_1363;
  assign T_1366 = io_inner_finish_bits_manager_xact_id & 3'h3;
  assign T_1368 = io_inner_finish_bits_manager_xact_id >= 3'h4;
  assign T_1370 = T_1366 & 3'h1;
  assign T_1372 = T_1366 >= 3'h2;
  assign T_1376 = T_1370 >= 3'h1;
  assign T_1377 = T_1376 ? trackerList_3_io_inner_finish_ready : trackerList_2_io_inner_finish_ready;
  assign T_1382 = T_1376 ? trackerList_1_io_inner_finish_ready : trackerList_0_io_inner_finish_ready;
  assign T_1383 = T_1372 ? T_1377 : T_1382;
  assign T_1384 = T_1368 ? trackerList_4_io_inner_finish_ready : T_1383;
  assign T_1388 = io_outer_probe_valid == 1'h0;
  assign T_1389 = T_1388 | reset;
  assign T_1391 = T_1389 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_4 = GEN_9[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_5 = {1{$random}};
  GEN_6 = {1{$random}};
  GEN_7 = {1{$random}};
  GEN_8 = {1{$random}};
  GEN_9 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1391) begin
          $fwrite(32'h80000002,"Assertion failed: L2 agent got illegal probe\n    at Agents.scala:160 assert(!io.outer.probe.valid, \"L2 agent got illegal probe\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1391) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module MMIOTileLinkManager(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  T_880;
  wire [2:0] T_889_0;
  wire  T_891;
  wire  T_892;
  wire  multibeat_fire;
  wire  T_894;
  wire  multibeat_start;
  wire  T_896;
  wire  multibeat_end;
  reg [5:0] xact_pending;
  reg [31:0] GEN_44;
  wire [5:0] T_898;
  wire  T_899;
  wire  T_900;
  wire  T_901;
  wire  T_902;
  wire  T_903;
  wire [2:0] T_911;
  wire [2:0] T_912;
  wire [2:0] T_913;
  wire [2:0] T_914;
  wire [2:0] xact_id_sel;
  reg [2:0] xact_id_reg;
  reg [31:0] GEN_45;
  wire [2:0] GEN_4;
  reg  xact_multibeat;
  reg [31:0] GEN_46;
  wire [2:0] outer_xact_id;
  wire  T_918;
  wire  xact_free;
  reg  xact_buffer_0_client_id;
  reg [31:0] GEN_47;
  reg [1:0] xact_buffer_0_client_xact_id;
  reg [31:0] GEN_48;
  reg  xact_buffer_1_client_id;
  reg [31:0] GEN_49;
  reg [1:0] xact_buffer_1_client_xact_id;
  reg [31:0] GEN_50;
  reg  xact_buffer_2_client_id;
  reg [31:0] GEN_51;
  reg [1:0] xact_buffer_2_client_xact_id;
  reg [31:0] GEN_52;
  reg  xact_buffer_3_client_id;
  reg [31:0] GEN_55;
  reg [1:0] xact_buffer_3_client_xact_id;
  reg [31:0] GEN_56;
  reg  xact_buffer_4_client_id;
  reg [31:0] GEN_57;
  reg [1:0] xact_buffer_4_client_xact_id;
  reg [31:0] GEN_58;
  reg  xact_buffer_5_client_id;
  reg [31:0] GEN_59;
  reg [1:0] xact_buffer_5_client_xact_id;
  reg [31:0] GEN_60;
  wire  T_1323;
  wire  T_1324;
  wire [2:0] T_1334_0;
  wire  T_1336;
  wire  T_1337;
  wire  T_1339;
  wire  T_1342;
  wire  T_1343;
  wire [3:0] T_1345;
  wire [3:0] T_1347;
  wire [5:0] GEN_2;
  wire [5:0] T_1348;
  wire  T_1349;
  wire [7:0] T_1351;
  wire [7:0] T_1353;
  wire [7:0] T_1354;
  wire [7:0] GEN_3;
  wire [7:0] T_1355;
  wire  T_1356;
  wire [2:0] T_1364_0;
  wire [3:0] GEN_53;
  wire  T_1366;
  wire  T_1367;
  wire  T_1368;
  wire  T_1371;
  wire  T_1373;
  wire  T_1374;
  wire  T_1375;
  wire  T_1381;
  wire  T_1383;
  wire  T_1386;
  wire  T_1387;
  wire [7:0] T_1389;
  wire [7:0] T_1391;
  wire [7:0] T_1392;
  wire [7:0] T_1393;
  wire [2:0] T_1403_0;
  wire  T_1405;
  wire  T_1406;
  wire  T_1408;
  wire  T_1411;
  wire  T_1412;
  wire  GEN_0;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] GEN_1;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [1:0] GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_2_client_id;
  wire [1:0] GEN_2_client_xact_id;
  wire  GEN_33;
  wire [1:0] GEN_34;
  wire  GEN_35;
  wire [1:0] GEN_36;
  wire  GEN_37;
  wire [1:0] GEN_38;
  wire [2:0] GEN_54;
  wire  GEN_39;
  wire [1:0] GEN_40;
  wire  GEN_41;
  wire [1:0] GEN_42;
  wire  GEN_3_client_id;
  wire [1:0] GEN_3_client_xact_id;
  wire [25:0] GEN_17;
  reg [31:0] GEN_61;
  wire [1:0] GEN_24;
  reg [31:0] GEN_62;
  wire  GEN_43;
  reg [31:0] GEN_63;
  assign io_inner_acquire_ready = T_1323;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = GEN_3_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = GEN_2_client_id;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_17;
  assign io_inner_probe_bits_p_type = GEN_24;
  assign io_inner_probe_bits_client_id = GEN_43;
  assign io_inner_release_ready = 1'h0;
  assign io_outer_acquire_valid = T_1324;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id[1:0];
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign T_880 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_889_0 = 3'h3;
  assign T_891 = io_outer_acquire_bits_a_type == T_889_0;
  assign T_892 = io_outer_acquire_bits_is_builtin_type & T_891;
  assign multibeat_fire = T_880 & T_892;
  assign T_894 = io_outer_acquire_bits_addr_beat == 3'h0;
  assign multibeat_start = multibeat_fire & T_894;
  assign T_896 = io_outer_acquire_bits_addr_beat == 3'h7;
  assign multibeat_end = multibeat_fire & T_896;
  assign T_898 = ~ xact_pending;
  assign T_899 = T_898[0];
  assign T_900 = T_898[1];
  assign T_901 = T_898[2];
  assign T_902 = T_898[3];
  assign T_903 = T_898[4];
  assign T_911 = T_903 ? 3'h4 : 3'h5;
  assign T_912 = T_902 ? 3'h3 : T_911;
  assign T_913 = T_901 ? 3'h2 : T_912;
  assign T_914 = T_900 ? 3'h1 : T_913;
  assign xact_id_sel = T_899 ? 3'h0 : T_914;
  assign GEN_4 = multibeat_start ? xact_id_sel : xact_id_reg;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : xact_id_sel;
  assign T_918 = T_898 == 6'h0;
  assign xact_free = T_918 == 1'h0;
  assign T_1323 = io_outer_acquire_ready & xact_free;
  assign T_1324 = io_inner_acquire_valid & xact_free;
  assign T_1334_0 = 3'h3;
  assign T_1336 = io_outer_acquire_bits_a_type == T_1334_0;
  assign T_1337 = io_outer_acquire_bits_is_builtin_type & T_1336;
  assign T_1339 = T_1337 == 1'h0;
  assign T_1342 = T_1339 | T_896;
  assign T_1343 = T_880 & T_1342;
  assign T_1345 = 4'h1 << io_outer_acquire_bits_client_xact_id;
  assign T_1347 = T_1343 ? T_1345 : 4'h0;
  assign GEN_2 = {{2'd0}, T_1347};
  assign T_1348 = xact_pending | GEN_2;
  assign T_1349 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_1351 = 8'h1 << io_inner_finish_bits_manager_xact_id;
  assign T_1353 = T_1349 ? T_1351 : 8'h0;
  assign T_1354 = ~ T_1353;
  assign GEN_3 = {{2'd0}, T_1348};
  assign T_1355 = GEN_3 & T_1354;
  assign T_1356 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1364_0 = 3'h5;
  assign GEN_53 = {{1'd0}, T_1364_0};
  assign T_1366 = io_inner_grant_bits_g_type == GEN_53;
  assign T_1367 = io_inner_grant_bits_g_type == 4'h0;
  assign T_1368 = io_inner_grant_bits_is_builtin_type ? T_1366 : T_1367;
  assign T_1371 = T_1368 == 1'h0;
  assign T_1373 = io_inner_grant_bits_addr_beat == 3'h7;
  assign T_1374 = T_1371 | T_1373;
  assign T_1375 = T_1356 & T_1374;
  assign T_1381 = io_inner_grant_bits_is_builtin_type & T_1367;
  assign T_1383 = T_1381 == 1'h0;
  assign T_1386 = T_1383 == 1'h0;
  assign T_1387 = T_1375 & T_1386;
  assign T_1389 = 8'h1 << io_inner_grant_bits_manager_xact_id;
  assign T_1391 = T_1387 ? T_1389 : 8'h0;
  assign T_1392 = ~ T_1391;
  assign T_1393 = T_1355 & T_1392;
  assign T_1403_0 = 3'h3;
  assign T_1405 = io_outer_acquire_bits_a_type == T_1403_0;
  assign T_1406 = io_outer_acquire_bits_is_builtin_type & T_1405;
  assign T_1408 = T_1406 == 1'h0;
  assign T_1411 = T_1408 | T_896;
  assign T_1412 = T_880 & T_1411;
  assign GEN_0 = io_inner_acquire_bits_client_id;
  assign GEN_5 = 3'h0 == outer_xact_id ? GEN_0 : xact_buffer_0_client_id;
  assign GEN_6 = 3'h1 == outer_xact_id ? GEN_0 : xact_buffer_1_client_id;
  assign GEN_7 = 3'h2 == outer_xact_id ? GEN_0 : xact_buffer_2_client_id;
  assign GEN_8 = 3'h3 == outer_xact_id ? GEN_0 : xact_buffer_3_client_id;
  assign GEN_9 = 3'h4 == outer_xact_id ? GEN_0 : xact_buffer_4_client_id;
  assign GEN_10 = 3'h5 == outer_xact_id ? GEN_0 : xact_buffer_5_client_id;
  assign GEN_1 = io_inner_acquire_bits_client_xact_id;
  assign GEN_11 = 3'h0 == outer_xact_id ? GEN_1 : xact_buffer_0_client_xact_id;
  assign GEN_12 = 3'h1 == outer_xact_id ? GEN_1 : xact_buffer_1_client_xact_id;
  assign GEN_13 = 3'h2 == outer_xact_id ? GEN_1 : xact_buffer_2_client_xact_id;
  assign GEN_14 = 3'h3 == outer_xact_id ? GEN_1 : xact_buffer_3_client_xact_id;
  assign GEN_15 = 3'h4 == outer_xact_id ? GEN_1 : xact_buffer_4_client_xact_id;
  assign GEN_16 = 3'h5 == outer_xact_id ? GEN_1 : xact_buffer_5_client_xact_id;
  assign GEN_18 = T_1412 ? GEN_5 : xact_buffer_0_client_id;
  assign GEN_19 = T_1412 ? GEN_6 : xact_buffer_1_client_id;
  assign GEN_20 = T_1412 ? GEN_7 : xact_buffer_2_client_id;
  assign GEN_21 = T_1412 ? GEN_8 : xact_buffer_3_client_id;
  assign GEN_22 = T_1412 ? GEN_9 : xact_buffer_4_client_id;
  assign GEN_23 = T_1412 ? GEN_10 : xact_buffer_5_client_id;
  assign GEN_25 = T_1412 ? GEN_11 : xact_buffer_0_client_xact_id;
  assign GEN_26 = T_1412 ? GEN_12 : xact_buffer_1_client_xact_id;
  assign GEN_27 = T_1412 ? GEN_13 : xact_buffer_2_client_xact_id;
  assign GEN_28 = T_1412 ? GEN_14 : xact_buffer_3_client_xact_id;
  assign GEN_29 = T_1412 ? GEN_15 : xact_buffer_4_client_xact_id;
  assign GEN_30 = T_1412 ? GEN_16 : xact_buffer_5_client_xact_id;
  assign GEN_31 = multibeat_start ? 1'h1 : xact_multibeat;
  assign GEN_32 = multibeat_end ? 1'h0 : GEN_31;
  assign GEN_2_client_id = GEN_41;
  assign GEN_2_client_xact_id = GEN_42;
  assign GEN_33 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign GEN_34 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign GEN_35 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_id : GEN_33;
  assign GEN_36 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_xact_id : GEN_34;
  assign GEN_37 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_id : GEN_35;
  assign GEN_38 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_xact_id : GEN_36;
  assign GEN_54 = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign GEN_39 = 3'h4 == GEN_54 ? xact_buffer_4_client_id : GEN_37;
  assign GEN_40 = 3'h4 == GEN_54 ? xact_buffer_4_client_xact_id : GEN_38;
  assign GEN_41 = 3'h5 == GEN_54 ? xact_buffer_5_client_id : GEN_39;
  assign GEN_42 = 3'h5 == GEN_54 ? xact_buffer_5_client_xact_id : GEN_40;
  assign GEN_3_client_id = GEN_41;
  assign GEN_3_client_xact_id = GEN_42;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_17 = GEN_61[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_24 = GEN_62[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_43 = GEN_63[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  xact_pending = GEN_44[5:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_45 = {1{$random}};
  xact_id_reg = GEN_45[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_46 = {1{$random}};
  xact_multibeat = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_47 = {1{$random}};
  xact_buffer_0_client_id = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  xact_buffer_0_client_xact_id = GEN_48[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_49 = {1{$random}};
  xact_buffer_1_client_id = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  xact_buffer_1_client_xact_id = GEN_50[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_51 = {1{$random}};
  xact_buffer_2_client_id = GEN_51[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  xact_buffer_2_client_xact_id = GEN_52[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_55 = {1{$random}};
  xact_buffer_3_client_id = GEN_55[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_56 = {1{$random}};
  xact_buffer_3_client_xact_id = GEN_56[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  xact_buffer_4_client_id = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  xact_buffer_4_client_xact_id = GEN_58[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  xact_buffer_5_client_id = GEN_59[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_60 = {1{$random}};
  xact_buffer_5_client_xact_id = GEN_60[1:0];
  `endif
  GEN_61 = {1{$random}};
  GEN_62 = {1{$random}};
  GEN_63 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      xact_pending <= 6'h0;
    end else begin
      xact_pending <= T_1393[5:0];
    end
    if(1'h0) begin
    end else begin
      if(multibeat_start) begin
        if(T_899) begin
          xact_id_reg <= 3'h0;
        end else begin
          if(T_900) begin
            xact_id_reg <= 3'h1;
          end else begin
            if(T_901) begin
              xact_id_reg <= 3'h2;
            end else begin
              if(T_902) begin
                xact_id_reg <= 3'h3;
              end else begin
                if(T_903) begin
                  xact_id_reg <= 3'h4;
                end else begin
                  xact_id_reg <= 3'h5;
                end
              end
            end
          end
        end
      end
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else begin
      if(multibeat_end) begin
        xact_multibeat <= 1'h0;
      end else begin
        if(multibeat_start) begin
          xact_multibeat <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h0 == outer_xact_id) begin
          xact_buffer_0_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h0 == outer_xact_id) begin
          xact_buffer_0_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h1 == outer_xact_id) begin
          xact_buffer_1_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h1 == outer_xact_id) begin
          xact_buffer_1_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h2 == outer_xact_id) begin
          xact_buffer_2_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h2 == outer_xact_id) begin
          xact_buffer_2_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h3 == outer_xact_id) begin
          xact_buffer_3_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h3 == outer_xact_id) begin
          xact_buffer_3_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h4 == outer_xact_id) begin
          xact_buffer_4_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h4 == outer_xact_id) begin
          xact_buffer_4_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h5 == outer_xact_id) begin
          xact_buffer_5_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1412) begin
        if(3'h5 == outer_xact_id) begin
          xact_buffer_5_client_xact_id <= GEN_1;
        end
      end
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module TileLinkMemoryInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [2:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [2:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIOArbiter_1_1_clk;
  wire  ClientUncachedTileLinkIOArbiter_1_1_reset;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data;
  wire [25:0] T_3009;
  ClientUncachedTileLinkIOArbiter_1 ClientUncachedTileLinkIOArbiter_1_1 (
    .clk(ClientUncachedTileLinkIOArbiter_1_1_clk),
    .reset(ClientUncachedTileLinkIOArbiter_1_1_reset),
    .io_in_0_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data),
    .io_out_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready),
    .io_out_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = T_3009;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_clk = clk;
  assign ClientUncachedTileLinkIOArbiter_1_1_reset = reset;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data = io_out_0_grant_bits_data;
  assign T_3009 = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block >> 1'h0;
endmodule
module LockingRRArbiter_9(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [10:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [10:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [10:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [25:0] GEN_0_bits_addr_block;
  wire [2:0] GEN_0_bits_client_xact_id;
  wire [2:0] GEN_0_bits_addr_beat;
  wire  GEN_0_bits_is_builtin_type;
  wire [2:0] GEN_0_bits_a_type;
  wire [10:0] GEN_0_bits_union;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_10;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire [10:0] GEN_15;
  wire [63:0] GEN_16;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [25:0] GEN_1_bits_addr_block;
  wire [2:0] GEN_1_bits_client_xact_id;
  wire [2:0] GEN_1_bits_addr_beat;
  wire  GEN_1_bits_is_builtin_type;
  wire [2:0] GEN_1_bits_a_type;
  wire [10:0] GEN_1_bits_union;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [25:0] GEN_2_bits_addr_block;
  wire [2:0] GEN_2_bits_client_xact_id;
  wire [2:0] GEN_2_bits_addr_beat;
  wire  GEN_2_bits_is_builtin_type;
  wire [2:0] GEN_2_bits_a_type;
  wire [10:0] GEN_2_bits_union;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [25:0] GEN_3_bits_addr_block;
  wire [2:0] GEN_3_bits_client_xact_id;
  wire [2:0] GEN_3_bits_addr_beat;
  wire  GEN_3_bits_is_builtin_type;
  wire [2:0] GEN_3_bits_a_type;
  wire [10:0] GEN_3_bits_union;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [25:0] GEN_4_bits_addr_block;
  wire [2:0] GEN_4_bits_client_xact_id;
  wire [2:0] GEN_4_bits_addr_beat;
  wire  GEN_4_bits_is_builtin_type;
  wire [2:0] GEN_4_bits_a_type;
  wire [10:0] GEN_4_bits_union;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [25:0] GEN_5_bits_addr_block;
  wire [2:0] GEN_5_bits_client_xact_id;
  wire [2:0] GEN_5_bits_addr_beat;
  wire  GEN_5_bits_is_builtin_type;
  wire [2:0] GEN_5_bits_a_type;
  wire [10:0] GEN_5_bits_union;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [25:0] GEN_6_bits_addr_block;
  wire [2:0] GEN_6_bits_client_xact_id;
  wire [2:0] GEN_6_bits_addr_beat;
  wire  GEN_6_bits_is_builtin_type;
  wire [2:0] GEN_6_bits_a_type;
  wire [10:0] GEN_6_bits_union;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [25:0] GEN_7_bits_addr_block;
  wire [2:0] GEN_7_bits_client_xact_id;
  wire [2:0] GEN_7_bits_addr_beat;
  wire  GEN_7_bits_is_builtin_type;
  wire [2:0] GEN_7_bits_a_type;
  wire [10:0] GEN_7_bits_union;
  wire [63:0] GEN_7_bits_data;
  reg [2:0] T_766;
  reg [31:0] GEN_0;
  reg  T_768;
  reg [31:0] GEN_1;
  wire  T_770;
  wire [2:0] T_779_0;
  wire  T_781;
  wire  T_782;
  wire  T_783;
  wire  T_784;
  wire [3:0] T_788;
  wire [2:0] T_789;
  wire  GEN_80;
  wire [2:0] GEN_81;
  wire  GEN_82;
  reg  lastGrant;
  reg [31:0] GEN_2;
  wire  GEN_83;
  wire  grantMask_1;
  wire  validMask_1;
  wire  T_795;
  wire  T_799;
  wire  T_801;
  wire  T_805;
  wire  T_807;
  wire  T_808;
  wire  T_809;
  wire  T_812;
  wire  T_813;
  wire  GEN_84;
  wire  GEN_85;
  assign io_in_0_ready = T_809;
  assign io_in_1_ready = T_813;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_block = GEN_1_bits_addr_block;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_addr_beat = GEN_3_bits_addr_beat;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_a_type = GEN_5_bits_a_type;
  assign io_out_bits_union = GEN_6_bits_union;
  assign io_out_bits_data = GEN_7_bits_data;
  assign io_chosen = GEN_82;
  assign choice = GEN_85;
  assign GEN_0_ready = GEN_8;
  assign GEN_0_valid = GEN_9;
  assign GEN_0_bits_addr_block = GEN_10;
  assign GEN_0_bits_client_xact_id = GEN_11;
  assign GEN_0_bits_addr_beat = GEN_12;
  assign GEN_0_bits_is_builtin_type = GEN_13;
  assign GEN_0_bits_a_type = GEN_14;
  assign GEN_0_bits_union = GEN_15;
  assign GEN_0_bits_data = GEN_16;
  assign GEN_8 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_15 = io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_16 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_1_ready = GEN_8;
  assign GEN_1_valid = GEN_9;
  assign GEN_1_bits_addr_block = GEN_10;
  assign GEN_1_bits_client_xact_id = GEN_11;
  assign GEN_1_bits_addr_beat = GEN_12;
  assign GEN_1_bits_is_builtin_type = GEN_13;
  assign GEN_1_bits_a_type = GEN_14;
  assign GEN_1_bits_union = GEN_15;
  assign GEN_1_bits_data = GEN_16;
  assign GEN_2_ready = GEN_8;
  assign GEN_2_valid = GEN_9;
  assign GEN_2_bits_addr_block = GEN_10;
  assign GEN_2_bits_client_xact_id = GEN_11;
  assign GEN_2_bits_addr_beat = GEN_12;
  assign GEN_2_bits_is_builtin_type = GEN_13;
  assign GEN_2_bits_a_type = GEN_14;
  assign GEN_2_bits_union = GEN_15;
  assign GEN_2_bits_data = GEN_16;
  assign GEN_3_ready = GEN_8;
  assign GEN_3_valid = GEN_9;
  assign GEN_3_bits_addr_block = GEN_10;
  assign GEN_3_bits_client_xact_id = GEN_11;
  assign GEN_3_bits_addr_beat = GEN_12;
  assign GEN_3_bits_is_builtin_type = GEN_13;
  assign GEN_3_bits_a_type = GEN_14;
  assign GEN_3_bits_union = GEN_15;
  assign GEN_3_bits_data = GEN_16;
  assign GEN_4_ready = GEN_8;
  assign GEN_4_valid = GEN_9;
  assign GEN_4_bits_addr_block = GEN_10;
  assign GEN_4_bits_client_xact_id = GEN_11;
  assign GEN_4_bits_addr_beat = GEN_12;
  assign GEN_4_bits_is_builtin_type = GEN_13;
  assign GEN_4_bits_a_type = GEN_14;
  assign GEN_4_bits_union = GEN_15;
  assign GEN_4_bits_data = GEN_16;
  assign GEN_5_ready = GEN_8;
  assign GEN_5_valid = GEN_9;
  assign GEN_5_bits_addr_block = GEN_10;
  assign GEN_5_bits_client_xact_id = GEN_11;
  assign GEN_5_bits_addr_beat = GEN_12;
  assign GEN_5_bits_is_builtin_type = GEN_13;
  assign GEN_5_bits_a_type = GEN_14;
  assign GEN_5_bits_union = GEN_15;
  assign GEN_5_bits_data = GEN_16;
  assign GEN_6_ready = GEN_8;
  assign GEN_6_valid = GEN_9;
  assign GEN_6_bits_addr_block = GEN_10;
  assign GEN_6_bits_client_xact_id = GEN_11;
  assign GEN_6_bits_addr_beat = GEN_12;
  assign GEN_6_bits_is_builtin_type = GEN_13;
  assign GEN_6_bits_a_type = GEN_14;
  assign GEN_6_bits_union = GEN_15;
  assign GEN_6_bits_data = GEN_16;
  assign GEN_7_ready = GEN_8;
  assign GEN_7_valid = GEN_9;
  assign GEN_7_bits_addr_block = GEN_10;
  assign GEN_7_bits_client_xact_id = GEN_11;
  assign GEN_7_bits_addr_beat = GEN_12;
  assign GEN_7_bits_is_builtin_type = GEN_13;
  assign GEN_7_bits_a_type = GEN_14;
  assign GEN_7_bits_union = GEN_15;
  assign GEN_7_bits_data = GEN_16;
  assign T_770 = T_766 != 3'h0;
  assign T_779_0 = 3'h3;
  assign T_781 = io_out_bits_a_type == T_779_0;
  assign T_782 = io_out_bits_is_builtin_type & T_781;
  assign T_783 = io_out_ready & io_out_valid;
  assign T_784 = T_783 & T_782;
  assign T_788 = T_766 + 3'h1;
  assign T_789 = T_788[2:0];
  assign GEN_80 = T_784 ? io_chosen : T_768;
  assign GEN_81 = T_784 ? T_789 : T_766;
  assign GEN_82 = T_770 ? T_768 : choice;
  assign GEN_83 = T_783 ? io_chosen : lastGrant;
  assign grantMask_1 = 1'h1 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign T_795 = validMask_1 | io_in_0_valid;
  assign T_799 = validMask_1 == 1'h0;
  assign T_801 = T_795 == 1'h0;
  assign T_805 = grantMask_1 | T_801;
  assign T_807 = T_768 == 1'h0;
  assign T_808 = T_770 ? T_807 : T_799;
  assign T_809 = T_808 & io_out_ready;
  assign T_812 = T_770 ? T_768 : T_805;
  assign T_813 = T_812 & io_out_ready;
  assign GEN_84 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_85 = validMask_1 ? 1'h1 : GEN_84;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_0 = {1{$random}};
  T_766 = GEN_0[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_768 = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  lastGrant = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_784) begin
        T_766 <= T_789;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_784) begin
        T_768 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_783) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ReorderQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_data,
  input  [2:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [2:0] io_deq_tag,
  output  io_deq_data,
  output  io_deq_matches
);
  reg  T_31 [0:7];
  reg [31:0] GEN_26;
  wire  T_31_T_51_data;
  wire [2:0] T_31_T_51_addr;
  wire  T_31_T_51_en;
  wire  T_31_T_55_data;
  wire [2:0] T_31_T_55_addr;
  wire  T_31_T_55_mask;
  wire  T_31_T_55_en;
  wire  T_45_0;
  wire  T_45_1;
  wire  T_45_2;
  wire  T_45_3;
  wire  T_45_4;
  wire  T_45_5;
  wire  T_45_6;
  wire  T_45_7;
  reg  T_49_0;
  reg [31:0] GEN_27;
  reg  T_49_1;
  reg [31:0] GEN_28;
  reg  T_49_2;
  reg [31:0] GEN_29;
  reg  T_49_3;
  reg [31:0] GEN_30;
  reg  T_49_4;
  reg [31:0] GEN_31;
  reg  T_49_5;
  reg [31:0] GEN_48;
  reg  T_49_6;
  reg [31:0] GEN_57;
  reg  T_49_7;
  reg [31:0] GEN_58;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_1;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  T_53;
  wire  T_54;
  wire  GEN_2;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_3;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  assign io_enq_ready = GEN_0;
  assign io_deq_data = T_31_T_51_data;
  assign io_deq_matches = T_53;
  assign T_31_T_51_addr = io_deq_tag;
  assign T_31_T_51_en = 1'h1;
  assign T_31_T_51_data = T_31[T_31_T_51_addr];
  assign T_31_T_55_data = io_enq_bits_data;
  assign T_31_T_55_addr = io_enq_bits_tag;
  assign T_31_T_55_mask = T_54;
  assign T_31_T_55_en = T_54;
  assign T_45_0 = 1'h1;
  assign T_45_1 = 1'h1;
  assign T_45_2 = 1'h1;
  assign T_45_3 = 1'h1;
  assign T_45_4 = 1'h1;
  assign T_45_5 = 1'h1;
  assign T_45_6 = 1'h1;
  assign T_45_7 = 1'h1;
  assign GEN_0 = GEN_10;
  assign GEN_4 = 3'h1 == io_enq_bits_tag ? T_49_1 : T_49_0;
  assign GEN_5 = 3'h2 == io_enq_bits_tag ? T_49_2 : GEN_4;
  assign GEN_6 = 3'h3 == io_enq_bits_tag ? T_49_3 : GEN_5;
  assign GEN_7 = 3'h4 == io_enq_bits_tag ? T_49_4 : GEN_6;
  assign GEN_8 = 3'h5 == io_enq_bits_tag ? T_49_5 : GEN_7;
  assign GEN_9 = 3'h6 == io_enq_bits_tag ? T_49_6 : GEN_8;
  assign GEN_10 = 3'h7 == io_enq_bits_tag ? T_49_7 : GEN_9;
  assign GEN_1 = GEN_17;
  assign GEN_11 = 3'h1 == io_deq_tag ? T_49_1 : T_49_0;
  assign GEN_12 = 3'h2 == io_deq_tag ? T_49_2 : GEN_11;
  assign GEN_13 = 3'h3 == io_deq_tag ? T_49_3 : GEN_12;
  assign GEN_14 = 3'h4 == io_deq_tag ? T_49_4 : GEN_13;
  assign GEN_15 = 3'h5 == io_deq_tag ? T_49_5 : GEN_14;
  assign GEN_16 = 3'h6 == io_deq_tag ? T_49_6 : GEN_15;
  assign GEN_17 = 3'h7 == io_deq_tag ? T_49_7 : GEN_16;
  assign T_53 = GEN_1 == 1'h0;
  assign T_54 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_18 = 3'h0 == io_enq_bits_tag ? GEN_2 : T_49_0;
  assign GEN_19 = 3'h1 == io_enq_bits_tag ? GEN_2 : T_49_1;
  assign GEN_20 = 3'h2 == io_enq_bits_tag ? GEN_2 : T_49_2;
  assign GEN_21 = 3'h3 == io_enq_bits_tag ? GEN_2 : T_49_3;
  assign GEN_22 = 3'h4 == io_enq_bits_tag ? GEN_2 : T_49_4;
  assign GEN_23 = 3'h5 == io_enq_bits_tag ? GEN_2 : T_49_5;
  assign GEN_24 = 3'h6 == io_enq_bits_tag ? GEN_2 : T_49_6;
  assign GEN_25 = 3'h7 == io_enq_bits_tag ? GEN_2 : T_49_7;
  assign GEN_32 = T_54 ? GEN_18 : T_49_0;
  assign GEN_33 = T_54 ? GEN_19 : T_49_1;
  assign GEN_34 = T_54 ? GEN_20 : T_49_2;
  assign GEN_35 = T_54 ? GEN_21 : T_49_3;
  assign GEN_36 = T_54 ? GEN_22 : T_49_4;
  assign GEN_37 = T_54 ? GEN_23 : T_49_5;
  assign GEN_38 = T_54 ? GEN_24 : T_49_6;
  assign GEN_39 = T_54 ? GEN_25 : T_49_7;
  assign GEN_3 = 1'h1;
  assign GEN_40 = 3'h0 == io_deq_tag ? GEN_3 : GEN_32;
  assign GEN_41 = 3'h1 == io_deq_tag ? GEN_3 : GEN_33;
  assign GEN_42 = 3'h2 == io_deq_tag ? GEN_3 : GEN_34;
  assign GEN_43 = 3'h3 == io_deq_tag ? GEN_3 : GEN_35;
  assign GEN_44 = 3'h4 == io_deq_tag ? GEN_3 : GEN_36;
  assign GEN_45 = 3'h5 == io_deq_tag ? GEN_3 : GEN_37;
  assign GEN_46 = 3'h6 == io_deq_tag ? GEN_3 : GEN_38;
  assign GEN_47 = 3'h7 == io_deq_tag ? GEN_3 : GEN_39;
  assign GEN_49 = io_deq_valid ? GEN_40 : GEN_32;
  assign GEN_50 = io_deq_valid ? GEN_41 : GEN_33;
  assign GEN_51 = io_deq_valid ? GEN_42 : GEN_34;
  assign GEN_52 = io_deq_valid ? GEN_43 : GEN_35;
  assign GEN_53 = io_deq_valid ? GEN_44 : GEN_36;
  assign GEN_54 = io_deq_valid ? GEN_45 : GEN_37;
  assign GEN_55 = io_deq_valid ? GEN_46 : GEN_38;
  assign GEN_56 = io_deq_valid ? GEN_47 : GEN_39;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_26 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    T_31[initvar] = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  T_49_0 = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  T_49_1 = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  T_49_2 = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  T_49_3 = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  T_49_4 = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_48 = {1{$random}};
  T_49_5 = GEN_48[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_57 = {1{$random}};
  T_49_6 = GEN_57[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_58 = {1{$random}};
  T_49_7 = GEN_58[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_31_T_55_en & T_31_T_55_mask) begin
      T_31[T_31_T_55_addr] <= T_31_T_55_data;
    end
    if(reset) begin
      T_49_0 <= T_45_0;
    end else begin
      if(io_deq_valid) begin
        if(3'h0 == io_deq_tag) begin
          T_49_0 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h0 == io_enq_bits_tag) begin
              T_49_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h0 == io_enq_bits_tag) begin
            T_49_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_1 <= T_45_1;
    end else begin
      if(io_deq_valid) begin
        if(3'h1 == io_deq_tag) begin
          T_49_1 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h1 == io_enq_bits_tag) begin
              T_49_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h1 == io_enq_bits_tag) begin
            T_49_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_2 <= T_45_2;
    end else begin
      if(io_deq_valid) begin
        if(3'h2 == io_deq_tag) begin
          T_49_2 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h2 == io_enq_bits_tag) begin
              T_49_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h2 == io_enq_bits_tag) begin
            T_49_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_3 <= T_45_3;
    end else begin
      if(io_deq_valid) begin
        if(3'h3 == io_deq_tag) begin
          T_49_3 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h3 == io_enq_bits_tag) begin
              T_49_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h3 == io_enq_bits_tag) begin
            T_49_3 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_4 <= T_45_4;
    end else begin
      if(io_deq_valid) begin
        if(3'h4 == io_deq_tag) begin
          T_49_4 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h4 == io_enq_bits_tag) begin
              T_49_4 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h4 == io_enq_bits_tag) begin
            T_49_4 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_5 <= T_45_5;
    end else begin
      if(io_deq_valid) begin
        if(3'h5 == io_deq_tag) begin
          T_49_5 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h5 == io_enq_bits_tag) begin
              T_49_5 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h5 == io_enq_bits_tag) begin
            T_49_5 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_6 <= T_45_6;
    end else begin
      if(io_deq_valid) begin
        if(3'h6 == io_deq_tag) begin
          T_49_6 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h6 == io_enq_bits_tag) begin
              T_49_6 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h6 == io_enq_bits_tag) begin
            T_49_6 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_49_7 <= T_45_7;
    end else begin
      if(io_deq_valid) begin
        if(3'h7 == io_deq_tag) begin
          T_49_7 <= GEN_3;
        end else begin
          if(T_54) begin
            if(3'h7 == io_enq_bits_tag) begin
              T_49_7 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_54) begin
          if(3'h7 == io_enq_bits_tag) begin
            T_49_7 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module ClientTileLinkIOUnwrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [2:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_probe_ready,
  output  io_in_probe_valid,
  output [25:0] io_in_probe_bits_addr_block,
  output [1:0] io_in_probe_bits_p_type,
  output  io_in_release_ready,
  input   io_in_release_valid,
  input  [2:0] io_in_release_bits_addr_beat,
  input  [25:0] io_in_release_bits_addr_block,
  input  [2:0] io_in_release_bits_client_xact_id,
  input   io_in_release_bits_voluntary,
  input  [2:0] io_in_release_bits_r_type,
  input  [63:0] io_in_release_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [2:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  output  io_in_grant_bits_manager_id,
  output  io_in_finish_ready,
  input   io_in_finish_valid,
  input   io_in_finish_bits_manager_xact_id,
  input   io_in_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [10:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  wire  acqArb_clk;
  wire  acqArb_reset;
  wire  acqArb_io_in_0_ready;
  wire  acqArb_io_in_0_valid;
  wire [25:0] acqArb_io_in_0_bits_addr_block;
  wire [2:0] acqArb_io_in_0_bits_client_xact_id;
  wire [2:0] acqArb_io_in_0_bits_addr_beat;
  wire  acqArb_io_in_0_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_0_bits_a_type;
  wire [10:0] acqArb_io_in_0_bits_union;
  wire [63:0] acqArb_io_in_0_bits_data;
  wire  acqArb_io_in_1_ready;
  wire  acqArb_io_in_1_valid;
  wire [25:0] acqArb_io_in_1_bits_addr_block;
  wire [2:0] acqArb_io_in_1_bits_client_xact_id;
  wire [2:0] acqArb_io_in_1_bits_addr_beat;
  wire  acqArb_io_in_1_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_1_bits_a_type;
  wire [10:0] acqArb_io_in_1_bits_union;
  wire [63:0] acqArb_io_in_1_bits_data;
  wire  acqArb_io_out_ready;
  wire  acqArb_io_out_valid;
  wire [25:0] acqArb_io_out_bits_addr_block;
  wire [2:0] acqArb_io_out_bits_client_xact_id;
  wire [2:0] acqArb_io_out_bits_addr_beat;
  wire  acqArb_io_out_bits_is_builtin_type;
  wire [2:0] acqArb_io_out_bits_a_type;
  wire [10:0] acqArb_io_out_bits_union;
  wire [63:0] acqArb_io_out_bits_data;
  wire  acqArb_io_chosen;
  wire  acqRoq_clk;
  wire  acqRoq_reset;
  wire  acqRoq_io_enq_ready;
  wire  acqRoq_io_enq_valid;
  wire  acqRoq_io_enq_bits_data;
  wire [2:0] acqRoq_io_enq_bits_tag;
  wire  acqRoq_io_deq_valid;
  wire [2:0] acqRoq_io_deq_tag;
  wire  acqRoq_io_deq_data;
  wire  acqRoq_io_deq_matches;
  wire  relRoq_clk;
  wire  relRoq_reset;
  wire  relRoq_io_enq_ready;
  wire  relRoq_io_enq_valid;
  wire  relRoq_io_enq_bits_data;
  wire [2:0] relRoq_io_enq_bits_tag;
  wire  relRoq_io_deq_valid;
  wire [2:0] relRoq_io_deq_tag;
  wire  relRoq_io_deq_data;
  wire  relRoq_io_deq_matches;
  wire [2:0] T_1366_0;
  wire  T_1368;
  wire  T_1369;
  wire  T_1371;
  wire  T_1373;
  wire  acq_roq_enq;
  wire  T_1375;
  wire  T_1376;
  wire  T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1382;
  wire  T_1384;
  wire  rel_roq_enq;
  wire  T_1386;
  wire  acq_roq_ready;
  wire  T_1388;
  wire  rel_roq_ready;
  wire  T_1389;
  wire  T_1390;
  wire  T_1391;
  wire [2:0] T_1394;
  wire [25:0] T_1423_addr_block;
  wire [2:0] T_1423_client_xact_id;
  wire [2:0] T_1423_addr_beat;
  wire  T_1423_is_builtin_type;
  wire [2:0] T_1423_a_type;
  wire [10:0] T_1423_union;
  wire [63:0] T_1423_data;
  wire  T_1451;
  wire  T_1452;
  wire  T_1453;
  wire  T_1454;
  wire [25:0] T_1577_addr_block;
  wire [2:0] T_1577_client_xact_id;
  wire [2:0] T_1577_addr_beat;
  wire  T_1577_is_builtin_type;
  wire [2:0] T_1577_a_type;
  wire [10:0] T_1577_union;
  wire [63:0] T_1577_data;
  wire  T_1605;
  wire  T_1606;
  wire [2:0] T_1614_0;
  wire [3:0] GEN_0;
  wire  T_1616;
  wire  T_1617;
  wire  T_1618;
  wire  T_1621;
  wire  T_1623;
  wire  T_1624;
  wire  grant_deq_roq;
  wire  T_1625;
  wire  T_1627;
  wire  T_1628;
  wire  T_1630;
  wire  T_1631;
  wire  T_1632;
  wire  T_1633;
  wire  T_1635;
  wire [3:0] T_1636;
  wire [2:0] acq_grant_addr_beat;
  wire [2:0] acq_grant_client_xact_id;
  wire  acq_grant_manager_xact_id;
  wire  acq_grant_is_builtin_type;
  wire [3:0] acq_grant_g_type;
  wire [63:0] acq_grant_data;
  wire  T_1691;
  wire  T_1692;
  wire  T_1693;
  wire  T_1695;
  wire [2:0] rel_grant_addr_beat;
  wire [2:0] rel_grant_client_xact_id;
  wire  rel_grant_manager_xact_id;
  wire  rel_grant_is_builtin_type;
  wire [3:0] rel_grant_g_type;
  wire [63:0] rel_grant_data;
  wire [2:0] T_1751_addr_beat;
  wire [2:0] T_1751_client_xact_id;
  wire  T_1751_manager_xact_id;
  wire  T_1751_is_builtin_type;
  wire [3:0] T_1751_g_type;
  wire [63:0] T_1751_data;
  wire [25:0] GEN_1;
  reg [31:0] GEN_4;
  wire [1:0] GEN_2;
  reg [31:0] GEN_5;
  wire  GEN_3;
  reg [31:0] GEN_6;
  LockingRRArbiter_9 acqArb (
    .clk(acqArb_clk),
    .reset(acqArb_reset),
    .io_in_0_ready(acqArb_io_in_0_ready),
    .io_in_0_valid(acqArb_io_in_0_valid),
    .io_in_0_bits_addr_block(acqArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(acqArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(acqArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(acqArb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(acqArb_io_in_0_bits_a_type),
    .io_in_0_bits_union(acqArb_io_in_0_bits_union),
    .io_in_0_bits_data(acqArb_io_in_0_bits_data),
    .io_in_1_ready(acqArb_io_in_1_ready),
    .io_in_1_valid(acqArb_io_in_1_valid),
    .io_in_1_bits_addr_block(acqArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(acqArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(acqArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(acqArb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(acqArb_io_in_1_bits_a_type),
    .io_in_1_bits_union(acqArb_io_in_1_bits_union),
    .io_in_1_bits_data(acqArb_io_in_1_bits_data),
    .io_out_ready(acqArb_io_out_ready),
    .io_out_valid(acqArb_io_out_valid),
    .io_out_bits_addr_block(acqArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(acqArb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(acqArb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(acqArb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(acqArb_io_out_bits_a_type),
    .io_out_bits_union(acqArb_io_out_bits_union),
    .io_out_bits_data(acqArb_io_out_bits_data),
    .io_chosen(acqArb_io_chosen)
  );
  ReorderQueue acqRoq (
    .clk(acqRoq_clk),
    .reset(acqRoq_reset),
    .io_enq_ready(acqRoq_io_enq_ready),
    .io_enq_valid(acqRoq_io_enq_valid),
    .io_enq_bits_data(acqRoq_io_enq_bits_data),
    .io_enq_bits_tag(acqRoq_io_enq_bits_tag),
    .io_deq_valid(acqRoq_io_deq_valid),
    .io_deq_tag(acqRoq_io_deq_tag),
    .io_deq_data(acqRoq_io_deq_data),
    .io_deq_matches(acqRoq_io_deq_matches)
  );
  ReorderQueue relRoq (
    .clk(relRoq_clk),
    .reset(relRoq_reset),
    .io_enq_ready(relRoq_io_enq_ready),
    .io_enq_valid(relRoq_io_enq_valid),
    .io_enq_bits_data(relRoq_io_enq_bits_data),
    .io_enq_bits_tag(relRoq_io_enq_bits_tag),
    .io_deq_valid(relRoq_io_deq_valid),
    .io_deq_tag(relRoq_io_deq_tag),
    .io_deq_data(relRoq_io_deq_data),
    .io_deq_matches(relRoq_io_deq_matches)
  );
  assign io_in_acquire_ready = T_1451;
  assign io_in_probe_valid = 1'h0;
  assign io_in_probe_bits_addr_block = GEN_1;
  assign io_in_probe_bits_p_type = GEN_2;
  assign io_in_release_ready = T_1605;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = T_1751_addr_beat;
  assign io_in_grant_bits_client_xact_id = T_1751_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = T_1751_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = T_1751_is_builtin_type;
  assign io_in_grant_bits_g_type = T_1751_g_type;
  assign io_in_grant_bits_data = T_1751_data;
  assign io_in_grant_bits_manager_id = GEN_3;
  assign io_in_finish_ready = 1'h0;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_grant_ready = io_in_grant_ready;
  assign acqArb_clk = clk;
  assign acqArb_reset = reset;
  assign acqArb_io_in_0_valid = T_1391;
  assign acqArb_io_in_0_bits_addr_block = T_1423_addr_block;
  assign acqArb_io_in_0_bits_client_xact_id = T_1423_client_xact_id;
  assign acqArb_io_in_0_bits_addr_beat = T_1423_addr_beat;
  assign acqArb_io_in_0_bits_is_builtin_type = T_1423_is_builtin_type;
  assign acqArb_io_in_0_bits_a_type = T_1423_a_type;
  assign acqArb_io_in_0_bits_union = T_1423_union;
  assign acqArb_io_in_0_bits_data = T_1423_data;
  assign acqArb_io_in_1_valid = T_1454;
  assign acqArb_io_in_1_bits_addr_block = T_1577_addr_block;
  assign acqArb_io_in_1_bits_client_xact_id = T_1577_client_xact_id;
  assign acqArb_io_in_1_bits_addr_beat = T_1577_addr_beat;
  assign acqArb_io_in_1_bits_is_builtin_type = T_1577_is_builtin_type;
  assign acqArb_io_in_1_bits_a_type = T_1577_a_type;
  assign acqArb_io_in_1_bits_union = T_1577_union;
  assign acqArb_io_in_1_bits_data = T_1577_data;
  assign acqArb_io_out_ready = io_out_acquire_ready;
  assign acqRoq_clk = clk;
  assign acqRoq_reset = reset;
  assign acqRoq_io_enq_valid = T_1390;
  assign acqRoq_io_enq_bits_data = io_in_acquire_bits_is_builtin_type;
  assign acqRoq_io_enq_bits_tag = io_in_acquire_bits_client_xact_id;
  assign acqRoq_io_deq_valid = T_1625;
  assign acqRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign relRoq_clk = clk;
  assign relRoq_reset = reset;
  assign relRoq_io_enq_valid = T_1453;
  assign relRoq_io_enq_bits_data = io_in_release_bits_voluntary;
  assign relRoq_io_enq_bits_tag = io_in_release_bits_client_xact_id;
  assign relRoq_io_deq_valid = T_1628;
  assign relRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign T_1366_0 = 3'h3;
  assign T_1368 = io_in_acquire_bits_a_type == T_1366_0;
  assign T_1369 = io_in_acquire_bits_is_builtin_type & T_1368;
  assign T_1371 = T_1369 == 1'h0;
  assign T_1373 = io_in_acquire_bits_addr_beat == 3'h0;
  assign acq_roq_enq = T_1371 | T_1373;
  assign T_1375 = io_in_release_bits_r_type == 3'h0;
  assign T_1376 = io_in_release_bits_r_type == 3'h1;
  assign T_1377 = io_in_release_bits_r_type == 3'h2;
  assign T_1378 = T_1375 | T_1376;
  assign T_1379 = T_1378 | T_1377;
  assign T_1382 = T_1379 == 1'h0;
  assign T_1384 = io_in_release_bits_addr_beat == 3'h0;
  assign rel_roq_enq = T_1382 | T_1384;
  assign T_1386 = acq_roq_enq == 1'h0;
  assign acq_roq_ready = T_1386 | acqRoq_io_enq_ready;
  assign T_1388 = rel_roq_enq == 1'h0;
  assign rel_roq_ready = T_1388 | relRoq_io_enq_ready;
  assign T_1389 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T_1390 = T_1389 & acq_roq_enq;
  assign T_1391 = io_in_acquire_valid & acq_roq_ready;
  assign T_1394 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T_1423_addr_block = io_in_acquire_bits_addr_block;
  assign T_1423_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign T_1423_addr_beat = io_in_acquire_bits_addr_beat;
  assign T_1423_is_builtin_type = 1'h1;
  assign T_1423_a_type = T_1394;
  assign T_1423_union = io_in_acquire_bits_union;
  assign T_1423_data = io_in_acquire_bits_data;
  assign T_1451 = acq_roq_ready & acqArb_io_in_0_ready;
  assign T_1452 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T_1453 = T_1452 & rel_roq_enq;
  assign T_1454 = io_in_release_valid & rel_roq_ready;
  assign T_1577_addr_block = io_in_release_bits_addr_block;
  assign T_1577_client_xact_id = io_in_release_bits_client_xact_id;
  assign T_1577_addr_beat = io_in_release_bits_addr_beat;
  assign T_1577_is_builtin_type = 1'h1;
  assign T_1577_a_type = 3'h3;
  assign T_1577_union = 11'h1ff;
  assign T_1577_data = io_in_release_bits_data;
  assign T_1605 = rel_roq_ready & acqArb_io_in_1_ready;
  assign T_1606 = io_out_grant_ready & io_out_grant_valid;
  assign T_1614_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1614_0};
  assign T_1616 = io_out_grant_bits_g_type == GEN_0;
  assign T_1617 = io_out_grant_bits_g_type == 4'h0;
  assign T_1618 = io_out_grant_bits_is_builtin_type ? T_1616 : T_1617;
  assign T_1621 = T_1618 == 1'h0;
  assign T_1623 = io_out_grant_bits_addr_beat == 3'h7;
  assign T_1624 = T_1621 | T_1623;
  assign grant_deq_roq = T_1606 & T_1624;
  assign T_1625 = acqRoq_io_deq_matches & grant_deq_roq;
  assign T_1627 = acqRoq_io_deq_matches == 1'h0;
  assign T_1628 = T_1627 & grant_deq_roq;
  assign T_1630 = grant_deq_roq == 1'h0;
  assign T_1631 = T_1630 | acqRoq_io_deq_matches;
  assign T_1632 = T_1631 | relRoq_io_deq_matches;
  assign T_1633 = T_1632 | reset;
  assign T_1635 = T_1633 == 1'h0;
  assign T_1636 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign acq_grant_g_type = T_1636;
  assign acq_grant_data = io_out_grant_bits_data;
  assign T_1691 = io_in_release_valid == 1'h0;
  assign T_1692 = T_1691 | io_in_release_bits_voluntary;
  assign T_1693 = T_1692 | reset;
  assign T_1695 = T_1693 == 1'h0;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign rel_grant_is_builtin_type = 1'h1;
  assign rel_grant_g_type = 4'h0;
  assign rel_grant_data = io_out_grant_bits_data;
  assign T_1751_addr_beat = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign T_1751_client_xact_id = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign T_1751_manager_xact_id = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign T_1751_is_builtin_type = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign T_1751_g_type = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign T_1751_data = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_4[25:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_2 = GEN_5[1:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_3 = GEN_6[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_4 = {1{$random}};
  GEN_5 = {1{$random}};
  GEN_6 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1635) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink Unwrapper: client_xact_id mismatch\n    at Tilelink.scala:120 assert(!grant_deq_roq || acqRoq.io.deq.matches || relRoq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1635) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1695) begin
          $fwrite(32'h80000002,"Assertion failed: Unwrapper can only process voluntary releases.\n    at Tilelink.scala:134 assert(!io.in.release.valid || io.in.release.bits.isVoluntary(), \"Unwrapper can only process voluntary releases.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1695) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [2:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [2:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [2:0] io_inner_grant_bits_client_xact_id,
  output  io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_manager_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input   io_inner_finish_bits_manager_xact_id,
  input   io_inner_finish_bits_manager_id,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign io_inner_finish_ready = io_outer_finish_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = io_inner_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = io_inner_finish_bits_manager_id;
endmodule
module Queue_14(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [10:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [10:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_304_data;
  wire  ram_addr_block_T_304_addr;
  wire  ram_addr_block_T_304_en;
  wire [25:0] ram_addr_block_T_269_data;
  wire  ram_addr_block_T_269_addr;
  wire  ram_addr_block_T_269_mask;
  wire  ram_addr_block_T_269_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_304_data;
  wire  ram_client_xact_id_T_304_addr;
  wire  ram_client_xact_id_T_304_en;
  wire [1:0] ram_client_xact_id_T_269_data;
  wire  ram_client_xact_id_T_269_addr;
  wire  ram_client_xact_id_T_269_mask;
  wire  ram_client_xact_id_T_269_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_304_data;
  wire  ram_addr_beat_T_304_addr;
  wire  ram_addr_beat_T_304_en;
  wire [2:0] ram_addr_beat_T_269_data;
  wire  ram_addr_beat_T_269_addr;
  wire  ram_addr_beat_T_269_mask;
  wire  ram_addr_beat_T_269_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_304_data;
  wire  ram_is_builtin_type_T_304_addr;
  wire  ram_is_builtin_type_T_304_en;
  wire  ram_is_builtin_type_T_269_data;
  wire  ram_is_builtin_type_T_269_addr;
  wire  ram_is_builtin_type_T_269_mask;
  wire  ram_is_builtin_type_T_269_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_304_data;
  wire  ram_a_type_T_304_addr;
  wire  ram_a_type_T_304_en;
  wire [2:0] ram_a_type_T_269_data;
  wire  ram_a_type_T_269_addr;
  wire  ram_a_type_T_269_mask;
  wire  ram_a_type_T_269_en;
  reg [10:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [10:0] ram_union_T_304_data;
  wire  ram_union_T_304_addr;
  wire  ram_union_T_304_en;
  wire [10:0] ram_union_T_269_data;
  wire  ram_union_T_269_addr;
  wire  ram_union_T_269_mask;
  wire  ram_union_T_269_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_304_data;
  wire  ram_data_T_304_addr;
  wire  ram_data_T_304_en;
  wire [63:0] ram_data_T_269_data;
  wire  ram_data_T_269_addr;
  wire  ram_data_T_269_mask;
  wire  ram_data_T_269_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_266;
  wire  T_267;
  wire  do_enq;
  wire  T_268;
  wire  do_deq;
  wire  T_299;
  wire  GEN_17;
  wire  T_301;
  wire [1:0] T_332;
  wire  ptr_diff;
  wire [1:0] T_334;
  assign io_enq_ready = T_266;
  assign io_deq_valid = T_301;
  assign io_deq_bits_addr_block = ram_addr_block_T_304_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_304_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_304_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_304_data;
  assign io_deq_bits_a_type = ram_a_type_T_304_data;
  assign io_deq_bits_union = ram_union_T_304_data;
  assign io_deq_bits_data = ram_data_T_304_data;
  assign io_count = T_334[0];
  assign ram_addr_block_T_304_addr = 1'h0;
  assign ram_addr_block_T_304_en = 1'h1;
  assign ram_addr_block_T_304_data = ram_addr_block[ram_addr_block_T_304_addr];
  assign ram_addr_block_T_269_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_269_addr = 1'h0;
  assign ram_addr_block_T_269_mask = do_enq;
  assign ram_addr_block_T_269_en = do_enq;
  assign ram_client_xact_id_T_304_addr = 1'h0;
  assign ram_client_xact_id_T_304_en = 1'h1;
  assign ram_client_xact_id_T_304_data = ram_client_xact_id[ram_client_xact_id_T_304_addr];
  assign ram_client_xact_id_T_269_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_269_addr = 1'h0;
  assign ram_client_xact_id_T_269_mask = do_enq;
  assign ram_client_xact_id_T_269_en = do_enq;
  assign ram_addr_beat_T_304_addr = 1'h0;
  assign ram_addr_beat_T_304_en = 1'h1;
  assign ram_addr_beat_T_304_data = ram_addr_beat[ram_addr_beat_T_304_addr];
  assign ram_addr_beat_T_269_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_269_addr = 1'h0;
  assign ram_addr_beat_T_269_mask = do_enq;
  assign ram_addr_beat_T_269_en = do_enq;
  assign ram_is_builtin_type_T_304_addr = 1'h0;
  assign ram_is_builtin_type_T_304_en = 1'h1;
  assign ram_is_builtin_type_T_304_data = ram_is_builtin_type[ram_is_builtin_type_T_304_addr];
  assign ram_is_builtin_type_T_269_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_269_addr = 1'h0;
  assign ram_is_builtin_type_T_269_mask = do_enq;
  assign ram_is_builtin_type_T_269_en = do_enq;
  assign ram_a_type_T_304_addr = 1'h0;
  assign ram_a_type_T_304_en = 1'h1;
  assign ram_a_type_T_304_data = ram_a_type[ram_a_type_T_304_addr];
  assign ram_a_type_T_269_data = io_enq_bits_a_type;
  assign ram_a_type_T_269_addr = 1'h0;
  assign ram_a_type_T_269_mask = do_enq;
  assign ram_a_type_T_269_en = do_enq;
  assign ram_union_T_304_addr = 1'h0;
  assign ram_union_T_304_en = 1'h1;
  assign ram_union_T_304_data = ram_union[ram_union_T_304_addr];
  assign ram_union_T_269_data = io_enq_bits_union;
  assign ram_union_T_269_addr = 1'h0;
  assign ram_union_T_269_mask = do_enq;
  assign ram_union_T_269_en = do_enq;
  assign ram_data_T_304_addr = 1'h0;
  assign ram_data_T_304_en = 1'h1;
  assign ram_data_T_304_data = ram_data[ram_data_T_304_addr];
  assign ram_data_T_269_data = io_enq_bits_data;
  assign ram_data_T_269_addr = 1'h0;
  assign ram_data_T_269_mask = do_enq;
  assign ram_data_T_269_en = do_enq;
  assign T_266 = maybe_full == 1'h0;
  assign T_267 = io_enq_ready & io_enq_valid;
  assign do_enq = T_267;
  assign T_268 = io_deq_ready & io_deq_valid;
  assign do_deq = T_268;
  assign T_299 = do_enq != do_deq;
  assign GEN_17 = T_299 ? do_enq : maybe_full;
  assign T_301 = T_266 == 1'h0;
  assign T_332 = 1'h0 - 1'h0;
  assign ptr_diff = T_332[0:0];
  assign T_334 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[10:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_269_en & ram_addr_block_T_269_mask) begin
      ram_addr_block[ram_addr_block_T_269_addr] <= ram_addr_block_T_269_data;
    end
    if(ram_client_xact_id_T_269_en & ram_client_xact_id_T_269_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_269_addr] <= ram_client_xact_id_T_269_data;
    end
    if(ram_addr_beat_T_269_en & ram_addr_beat_T_269_mask) begin
      ram_addr_beat[ram_addr_beat_T_269_addr] <= ram_addr_beat_T_269_data;
    end
    if(ram_is_builtin_type_T_269_en & ram_is_builtin_type_T_269_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_269_addr] <= ram_is_builtin_type_T_269_data;
    end
    if(ram_a_type_T_269_en & ram_a_type_T_269_mask) begin
      ram_a_type[ram_a_type_T_269_addr] <= ram_a_type_T_269_data;
    end
    if(ram_union_T_269_en & ram_union_T_269_mask) begin
      ram_union[ram_union_T_269_addr] <= ram_union_T_269_data;
    end
    if(ram_data_T_269_en & ram_data_T_269_mask) begin
      ram_data[ram_data_T_269_addr] <= ram_data_T_269_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_299) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_15(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_addr_beat,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_is_builtin_type,
  input  [3:0] io_enq_bits_g_type,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_addr_beat,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_is_builtin_type,
  output [3:0] io_deq_bits_g_type,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_addr_beat_T_294_data;
  wire  ram_addr_beat_T_294_addr;
  wire  ram_addr_beat_T_294_en;
  wire [2:0] ram_addr_beat_T_260_data;
  wire  ram_addr_beat_T_260_addr;
  wire  ram_addr_beat_T_260_mask;
  wire  ram_addr_beat_T_260_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_294_data;
  wire  ram_client_xact_id_T_294_addr;
  wire  ram_client_xact_id_T_294_en;
  wire [1:0] ram_client_xact_id_T_260_data;
  wire  ram_client_xact_id_T_260_addr;
  wire  ram_client_xact_id_T_260_mask;
  wire  ram_client_xact_id_T_260_en;
  reg [2:0] ram_manager_xact_id [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_manager_xact_id_T_294_data;
  wire  ram_manager_xact_id_T_294_addr;
  wire  ram_manager_xact_id_T_294_en;
  wire [2:0] ram_manager_xact_id_T_260_data;
  wire  ram_manager_xact_id_T_260_addr;
  wire  ram_manager_xact_id_T_260_mask;
  wire  ram_manager_xact_id_T_260_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_294_data;
  wire  ram_is_builtin_type_T_294_addr;
  wire  ram_is_builtin_type_T_294_en;
  wire  ram_is_builtin_type_T_260_data;
  wire  ram_is_builtin_type_T_260_addr;
  wire  ram_is_builtin_type_T_260_mask;
  wire  ram_is_builtin_type_T_260_en;
  reg [3:0] ram_g_type [0:0];
  reg [31:0] GEN_4;
  wire [3:0] ram_g_type_T_294_data;
  wire  ram_g_type_T_294_addr;
  wire  ram_g_type_T_294_en;
  wire [3:0] ram_g_type_T_260_data;
  wire  ram_g_type_T_260_addr;
  wire  ram_g_type_T_260_mask;
  wire  ram_g_type_T_260_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_5;
  wire [63:0] ram_data_T_294_data;
  wire  ram_data_T_294_addr;
  wire  ram_data_T_294_en;
  wire [63:0] ram_data_T_260_data;
  wire  ram_data_T_260_addr;
  wire  ram_data_T_260_mask;
  wire  ram_data_T_260_en;
  reg  maybe_full;
  reg [31:0] GEN_6;
  wire  T_257;
  wire  T_258;
  wire  do_enq;
  wire  T_259;
  wire  do_deq;
  wire  T_289;
  wire  GEN_15;
  wire  T_291;
  wire [1:0] T_321;
  wire  ptr_diff;
  wire [1:0] T_323;
  assign io_enq_ready = T_257;
  assign io_deq_valid = T_291;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_294_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_294_data;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_294_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_294_data;
  assign io_deq_bits_g_type = ram_g_type_T_294_data;
  assign io_deq_bits_data = ram_data_T_294_data;
  assign io_count = T_323[0];
  assign ram_addr_beat_T_294_addr = 1'h0;
  assign ram_addr_beat_T_294_en = 1'h1;
  assign ram_addr_beat_T_294_data = ram_addr_beat[ram_addr_beat_T_294_addr];
  assign ram_addr_beat_T_260_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_260_addr = 1'h0;
  assign ram_addr_beat_T_260_mask = do_enq;
  assign ram_addr_beat_T_260_en = do_enq;
  assign ram_client_xact_id_T_294_addr = 1'h0;
  assign ram_client_xact_id_T_294_en = 1'h1;
  assign ram_client_xact_id_T_294_data = ram_client_xact_id[ram_client_xact_id_T_294_addr];
  assign ram_client_xact_id_T_260_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_260_addr = 1'h0;
  assign ram_client_xact_id_T_260_mask = do_enq;
  assign ram_client_xact_id_T_260_en = do_enq;
  assign ram_manager_xact_id_T_294_addr = 1'h0;
  assign ram_manager_xact_id_T_294_en = 1'h1;
  assign ram_manager_xact_id_T_294_data = ram_manager_xact_id[ram_manager_xact_id_T_294_addr];
  assign ram_manager_xact_id_T_260_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_260_addr = 1'h0;
  assign ram_manager_xact_id_T_260_mask = do_enq;
  assign ram_manager_xact_id_T_260_en = do_enq;
  assign ram_is_builtin_type_T_294_addr = 1'h0;
  assign ram_is_builtin_type_T_294_en = 1'h1;
  assign ram_is_builtin_type_T_294_data = ram_is_builtin_type[ram_is_builtin_type_T_294_addr];
  assign ram_is_builtin_type_T_260_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_260_addr = 1'h0;
  assign ram_is_builtin_type_T_260_mask = do_enq;
  assign ram_is_builtin_type_T_260_en = do_enq;
  assign ram_g_type_T_294_addr = 1'h0;
  assign ram_g_type_T_294_en = 1'h1;
  assign ram_g_type_T_294_data = ram_g_type[ram_g_type_T_294_addr];
  assign ram_g_type_T_260_data = io_enq_bits_g_type;
  assign ram_g_type_T_260_addr = 1'h0;
  assign ram_g_type_T_260_mask = do_enq;
  assign ram_g_type_T_260_en = do_enq;
  assign ram_data_T_294_addr = 1'h0;
  assign ram_data_T_294_en = 1'h1;
  assign ram_data_T_294_data = ram_data[ram_data_T_294_addr];
  assign ram_data_T_260_data = io_enq_bits_data;
  assign ram_data_T_260_addr = 1'h0;
  assign ram_data_T_260_mask = do_enq;
  assign ram_data_T_260_en = do_enq;
  assign T_257 = maybe_full == 1'h0;
  assign T_258 = io_enq_ready & io_enq_valid;
  assign do_enq = T_258;
  assign T_259 = io_deq_ready & io_deq_valid;
  assign do_deq = T_259;
  assign T_289 = do_enq != do_deq;
  assign GEN_15 = T_289 ? do_enq : maybe_full;
  assign T_291 = T_257 == 1'h0;
  assign T_321 = 1'h0 - 1'h0;
  assign ptr_diff = T_321[0:0];
  assign T_323 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_0[2:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_g_type[initvar] = GEN_4[3:0];
  `endif
  GEN_5 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_5[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  maybe_full = GEN_6[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_beat_T_260_en & ram_addr_beat_T_260_mask) begin
      ram_addr_beat[ram_addr_beat_T_260_addr] <= ram_addr_beat_T_260_data;
    end
    if(ram_client_xact_id_T_260_en & ram_client_xact_id_T_260_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_260_addr] <= ram_client_xact_id_T_260_data;
    end
    if(ram_manager_xact_id_T_260_en & ram_manager_xact_id_T_260_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_260_addr] <= ram_manager_xact_id_T_260_data;
    end
    if(ram_is_builtin_type_T_260_en & ram_is_builtin_type_T_260_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_260_addr] <= ram_is_builtin_type_T_260_data;
    end
    if(ram_g_type_T_260_en & ram_g_type_T_260_mask) begin
      ram_g_type[ram_g_type_T_260_addr] <= ram_g_type_T_260_data;
    end
    if(ram_data_T_260_en & ram_data_T_260_mask) begin
      ram_data[ram_data_T_260_addr] <= ram_data_T_260_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_289) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module ClientUncachedTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [10:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [10:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input  [2:0] io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  Queue_14_1_clk;
  wire  Queue_14_1_reset;
  wire  Queue_14_1_io_enq_ready;
  wire  Queue_14_1_io_enq_valid;
  wire [25:0] Queue_14_1_io_enq_bits_addr_block;
  wire [1:0] Queue_14_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_14_1_io_enq_bits_addr_beat;
  wire  Queue_14_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_14_1_io_enq_bits_a_type;
  wire [10:0] Queue_14_1_io_enq_bits_union;
  wire [63:0] Queue_14_1_io_enq_bits_data;
  wire  Queue_14_1_io_deq_ready;
  wire  Queue_14_1_io_deq_valid;
  wire [25:0] Queue_14_1_io_deq_bits_addr_block;
  wire [1:0] Queue_14_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_14_1_io_deq_bits_addr_beat;
  wire  Queue_14_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_14_1_io_deq_bits_a_type;
  wire [10:0] Queue_14_1_io_deq_bits_union;
  wire [63:0] Queue_14_1_io_deq_bits_data;
  wire  Queue_14_1_io_count;
  wire  Queue_15_1_clk;
  wire  Queue_15_1_reset;
  wire  Queue_15_1_io_enq_ready;
  wire  Queue_15_1_io_enq_valid;
  wire [2:0] Queue_15_1_io_enq_bits_addr_beat;
  wire [1:0] Queue_15_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_15_1_io_enq_bits_manager_xact_id;
  wire  Queue_15_1_io_enq_bits_is_builtin_type;
  wire [3:0] Queue_15_1_io_enq_bits_g_type;
  wire [63:0] Queue_15_1_io_enq_bits_data;
  wire  Queue_15_1_io_deq_ready;
  wire  Queue_15_1_io_deq_valid;
  wire [2:0] Queue_15_1_io_deq_bits_addr_beat;
  wire [1:0] Queue_15_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_15_1_io_deq_bits_manager_xact_id;
  wire  Queue_15_1_io_deq_bits_is_builtin_type;
  wire [3:0] Queue_15_1_io_deq_bits_g_type;
  wire [63:0] Queue_15_1_io_deq_bits_data;
  wire  Queue_15_1_io_count;
  Queue_14 Queue_14_1 (
    .clk(Queue_14_1_clk),
    .reset(Queue_14_1_reset),
    .io_enq_ready(Queue_14_1_io_enq_ready),
    .io_enq_valid(Queue_14_1_io_enq_valid),
    .io_enq_bits_addr_block(Queue_14_1_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(Queue_14_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_14_1_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(Queue_14_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_14_1_io_enq_bits_a_type),
    .io_enq_bits_union(Queue_14_1_io_enq_bits_union),
    .io_enq_bits_data(Queue_14_1_io_enq_bits_data),
    .io_deq_ready(Queue_14_1_io_deq_ready),
    .io_deq_valid(Queue_14_1_io_deq_valid),
    .io_deq_bits_addr_block(Queue_14_1_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(Queue_14_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_14_1_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(Queue_14_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_14_1_io_deq_bits_a_type),
    .io_deq_bits_union(Queue_14_1_io_deq_bits_union),
    .io_deq_bits_data(Queue_14_1_io_deq_bits_data),
    .io_count(Queue_14_1_io_count)
  );
  Queue_15 Queue_15_1 (
    .clk(Queue_15_1_clk),
    .reset(Queue_15_1_reset),
    .io_enq_ready(Queue_15_1_io_enq_ready),
    .io_enq_valid(Queue_15_1_io_enq_valid),
    .io_enq_bits_addr_beat(Queue_15_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_xact_id(Queue_15_1_io_enq_bits_client_xact_id),
    .io_enq_bits_manager_xact_id(Queue_15_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_is_builtin_type(Queue_15_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_g_type(Queue_15_1_io_enq_bits_g_type),
    .io_enq_bits_data(Queue_15_1_io_enq_bits_data),
    .io_deq_ready(Queue_15_1_io_deq_ready),
    .io_deq_valid(Queue_15_1_io_deq_valid),
    .io_deq_bits_addr_beat(Queue_15_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_xact_id(Queue_15_1_io_deq_bits_client_xact_id),
    .io_deq_bits_manager_xact_id(Queue_15_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_is_builtin_type(Queue_15_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_g_type(Queue_15_1_io_deq_bits_g_type),
    .io_deq_bits_data(Queue_15_1_io_deq_bits_data),
    .io_count(Queue_15_1_io_count)
  );
  assign io_inner_acquire_ready = Queue_14_1_io_enq_ready;
  assign io_inner_grant_valid = Queue_15_1_io_deq_valid;
  assign io_inner_grant_bits_addr_beat = Queue_15_1_io_deq_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = Queue_15_1_io_deq_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = Queue_15_1_io_deq_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = Queue_15_1_io_deq_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = Queue_15_1_io_deq_bits_g_type;
  assign io_inner_grant_bits_data = Queue_15_1_io_deq_bits_data;
  assign io_outer_acquire_valid = Queue_14_1_io_deq_valid;
  assign io_outer_acquire_bits_addr_block = Queue_14_1_io_deq_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = Queue_14_1_io_deq_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = Queue_14_1_io_deq_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = Queue_14_1_io_deq_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = Queue_14_1_io_deq_bits_a_type;
  assign io_outer_acquire_bits_union = Queue_14_1_io_deq_bits_union;
  assign io_outer_acquire_bits_data = Queue_14_1_io_deq_bits_data;
  assign io_outer_grant_ready = Queue_15_1_io_enq_ready;
  assign Queue_14_1_clk = clk;
  assign Queue_14_1_reset = reset;
  assign Queue_14_1_io_enq_valid = io_inner_acquire_valid;
  assign Queue_14_1_io_enq_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign Queue_14_1_io_enq_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign Queue_14_1_io_enq_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign Queue_14_1_io_enq_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign Queue_14_1_io_enq_bits_a_type = io_inner_acquire_bits_a_type;
  assign Queue_14_1_io_enq_bits_union = io_inner_acquire_bits_union;
  assign Queue_14_1_io_enq_bits_data = io_inner_acquire_bits_data;
  assign Queue_14_1_io_deq_ready = io_outer_acquire_ready;
  assign Queue_15_1_clk = clk;
  assign Queue_15_1_reset = reset;
  assign Queue_15_1_io_enq_valid = io_outer_grant_valid;
  assign Queue_15_1_io_enq_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign Queue_15_1_io_enq_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign Queue_15_1_io_enq_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign Queue_15_1_io_enq_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign Queue_15_1_io_enq_bits_g_type = io_outer_grant_bits_g_type;
  assign Queue_15_1_io_enq_bits_data = io_outer_grant_bits_data;
  assign Queue_15_1_io_deq_ready = io_inner_grant_ready;
endmodule
module LockingRRArbiter_10(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_518;
  reg [31:0] GEN_1;
  reg  T_520;
  reg [31:0] GEN_2;
  wire  T_522;
  wire [2:0] T_530_0;
  wire [3:0] GEN_0;
  wire  T_532;
  wire  T_533;
  wire  T_534;
  wire  T_536;
  wire  T_537;
  wire [3:0] T_541;
  wire [2:0] T_542;
  wire  GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_9;
  reg  lastGrant;
  reg [31:0] GEN_3;
  wire  GEN_10;
  wire  T_551;
  wire  T_552;
  wire  T_553;
  assign io_in_0_ready = T_553;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_9;
  assign choice = 1'h0;
  assign GEN_0_ready = io_in_0_ready;
  assign GEN_0_valid = io_in_0_valid;
  assign GEN_0_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_0_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_0_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_0_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_0_bits_g_type = io_in_0_bits_g_type;
  assign GEN_0_bits_data = io_in_0_bits_data;
  assign GEN_1_ready = io_in_0_ready;
  assign GEN_1_valid = io_in_0_valid;
  assign GEN_1_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_1_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_1_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_1_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_1_bits_g_type = io_in_0_bits_g_type;
  assign GEN_1_bits_data = io_in_0_bits_data;
  assign GEN_2_ready = io_in_0_ready;
  assign GEN_2_valid = io_in_0_valid;
  assign GEN_2_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_2_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_2_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_2_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_2_bits_g_type = io_in_0_bits_g_type;
  assign GEN_2_bits_data = io_in_0_bits_data;
  assign GEN_3_ready = io_in_0_ready;
  assign GEN_3_valid = io_in_0_valid;
  assign GEN_3_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_3_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_3_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_3_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_3_bits_g_type = io_in_0_bits_g_type;
  assign GEN_3_bits_data = io_in_0_bits_data;
  assign GEN_4_ready = io_in_0_ready;
  assign GEN_4_valid = io_in_0_valid;
  assign GEN_4_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_4_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_4_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_4_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_4_bits_g_type = io_in_0_bits_g_type;
  assign GEN_4_bits_data = io_in_0_bits_data;
  assign GEN_5_ready = io_in_0_ready;
  assign GEN_5_valid = io_in_0_valid;
  assign GEN_5_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_5_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_5_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_5_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_5_bits_g_type = io_in_0_bits_g_type;
  assign GEN_5_bits_data = io_in_0_bits_data;
  assign GEN_6_ready = io_in_0_ready;
  assign GEN_6_valid = io_in_0_valid;
  assign GEN_6_bits_addr_beat = io_in_0_bits_addr_beat;
  assign GEN_6_bits_client_xact_id = io_in_0_bits_client_xact_id;
  assign GEN_6_bits_manager_xact_id = io_in_0_bits_manager_xact_id;
  assign GEN_6_bits_is_builtin_type = io_in_0_bits_is_builtin_type;
  assign GEN_6_bits_g_type = io_in_0_bits_g_type;
  assign GEN_6_bits_data = io_in_0_bits_data;
  assign T_522 = T_518 != 3'h0;
  assign T_530_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_530_0};
  assign T_532 = io_out_bits_g_type == GEN_0;
  assign T_533 = io_out_bits_g_type == 4'h0;
  assign T_534 = io_out_bits_is_builtin_type ? T_532 : T_533;
  assign T_536 = io_out_ready & io_out_valid;
  assign T_537 = T_536 & T_534;
  assign T_541 = T_518 + 3'h1;
  assign T_542 = T_541[2:0];
  assign GEN_7 = T_537 ? io_chosen : T_520;
  assign GEN_8 = T_537 ? T_542 : T_518;
  assign GEN_9 = T_522 ? T_520 : choice;
  assign GEN_10 = T_536 ? io_chosen : lastGrant;
  assign T_551 = T_520 == 1'h0;
  assign T_552 = T_522 ? T_551 : 1'h1;
  assign T_553 = T_552 & io_out_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_518 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_520 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_518 <= 3'h0;
    end else begin
      if(T_537) begin
        T_518 <= T_542;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_537) begin
        T_520 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_536) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire [2:0] T_1246_0;
  wire [2:0] T_1246_1;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1251;
  wire [2:0] T_1252;
  wire [2:0] T_1254;
  wire [28:0] T_1255;
  wire [31:0] T_1256;
  wire  T_1260;
  wire  T_1263;
  wire  T_1265;
  wire  T_1266;
  wire  T_1268;
  wire  T_1270;
  wire  T_1271;
  wire  T_1273;
  wire  T_1275;
  wire  T_1276;
  wire  T_1277;
  wire  T_1278;
  wire  acq_route;
  wire  T_1281;
  wire  GEN_0;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_chosen;
  wire  T_1306;
  wire  T_1309;
  wire  T_1310;
  wire  T_1312;
  LockingRRArbiter_10 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_0;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1281;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign T_1246_0 = 3'h0;
  assign T_1246_1 = 3'h4;
  assign T_1248 = io_in_acquire_bits_a_type == T_1246_0;
  assign T_1249 = io_in_acquire_bits_a_type == T_1246_1;
  assign T_1250 = T_1248 | T_1249;
  assign T_1251 = io_in_acquire_bits_is_builtin_type & T_1250;
  assign T_1252 = io_in_acquire_bits_union[10:8];
  assign T_1254 = T_1251 ? T_1252 : 3'h0;
  assign T_1255 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1256 = {T_1255,T_1254};
  assign T_1260 = T_1256 < 32'h1000;
  assign T_1263 = 32'h1000 <= T_1256;
  assign T_1265 = T_1256 < 32'h2000;
  assign T_1266 = T_1263 & T_1265;
  assign T_1268 = 32'h40000000 <= T_1256;
  assign T_1270 = T_1256 < 32'h44000000;
  assign T_1271 = T_1268 & T_1270;
  assign T_1273 = 32'h44000000 <= T_1256;
  assign T_1275 = T_1256 < 32'h48000000;
  assign T_1276 = T_1273 & T_1275;
  assign T_1277 = T_1260 | T_1266;
  assign T_1278 = T_1277 | T_1271;
  assign acq_route = T_1278 | T_1276;
  assign T_1281 = io_in_acquire_valid & acq_route;
  assign GEN_0 = acq_route ? io_out_0_acquire_ready : 1'h0;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1306 = io_in_acquire_valid == 1'h0;
  assign T_1309 = T_1306 | acq_route;
  assign T_1310 = T_1309 | reset;
  assign T_1312 = T_1310 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1312) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data;
  ClientUncachedTileLinkIORouter ClientUncachedTileLinkIORouter_1 (
    .clk(ClientUncachedTileLinkIORouter_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
endmodule
module LockingRRArbiter_11(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [1:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_9;
  wire [1:0] GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [3:0] GEN_13;
  wire [63:0] GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [3:0] GEN_21;
  wire [63:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_25;
  wire [1:0] GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire [3:0] GEN_29;
  wire [63:0] GEN_30;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [1:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [1:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [1:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [1:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [1:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [1:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  reg [2:0] T_794;
  reg [31:0] GEN_1;
  reg [1:0] T_796;
  reg [31:0] GEN_2;
  wire  T_798;
  wire [2:0] T_806_0;
  wire [3:0] GEN_0;
  wire  T_808;
  wire  T_809;
  wire  T_810;
  wire  T_812;
  wire  T_813;
  wire [3:0] T_817;
  wire [2:0] T_818;
  wire [1:0] GEN_175;
  wire [2:0] GEN_176;
  wire [1:0] GEN_177;
  reg [1:0] lastGrant;
  reg [31:0] GEN_3;
  wire [1:0] GEN_178;
  wire  grantMask_1;
  wire  grantMask_2;
  wire  grantMask_3;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  T_826;
  wire  T_827;
  wire  T_828;
  wire  T_829;
  wire  T_830;
  wire  T_834;
  wire  T_836;
  wire  T_838;
  wire  T_840;
  wire  T_842;
  wire  T_844;
  wire  T_848;
  wire  T_849;
  wire  T_850;
  wire  T_851;
  wire  T_852;
  wire  T_854;
  wire  T_855;
  wire  T_856;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_866;
  wire  T_867;
  wire  T_868;
  wire [1:0] GEN_179;
  wire [1:0] GEN_180;
  wire [1:0] GEN_181;
  wire [1:0] GEN_182;
  wire [1:0] GEN_183;
  wire [1:0] GEN_184;
  assign io_in_0_ready = T_856;
  assign io_in_1_ready = T_860;
  assign io_in_2_ready = T_864;
  assign io_in_3_ready = T_868;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_chosen = GEN_177;
  assign choice = GEN_184;
  assign GEN_0_ready = GEN_23;
  assign GEN_0_valid = GEN_24;
  assign GEN_0_bits_addr_beat = GEN_25;
  assign GEN_0_bits_client_xact_id = GEN_26;
  assign GEN_0_bits_manager_xact_id = GEN_27;
  assign GEN_0_bits_is_builtin_type = GEN_28;
  assign GEN_0_bits_g_type = GEN_29;
  assign GEN_0_bits_data = GEN_30;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_ready : GEN_7;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_9;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_10;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_11;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_12;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_g_type : GEN_13;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_14;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_ready : GEN_15;
  assign GEN_24 = 2'h3 == io_chosen ? io_in_3_valid : GEN_16;
  assign GEN_25 = 2'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_17;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_18;
  assign GEN_27 = 2'h3 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_19;
  assign GEN_28 = 2'h3 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_20;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_g_type : GEN_21;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_bits_data : GEN_22;
  assign GEN_1_ready = GEN_23;
  assign GEN_1_valid = GEN_24;
  assign GEN_1_bits_addr_beat = GEN_25;
  assign GEN_1_bits_client_xact_id = GEN_26;
  assign GEN_1_bits_manager_xact_id = GEN_27;
  assign GEN_1_bits_is_builtin_type = GEN_28;
  assign GEN_1_bits_g_type = GEN_29;
  assign GEN_1_bits_data = GEN_30;
  assign GEN_2_ready = GEN_23;
  assign GEN_2_valid = GEN_24;
  assign GEN_2_bits_addr_beat = GEN_25;
  assign GEN_2_bits_client_xact_id = GEN_26;
  assign GEN_2_bits_manager_xact_id = GEN_27;
  assign GEN_2_bits_is_builtin_type = GEN_28;
  assign GEN_2_bits_g_type = GEN_29;
  assign GEN_2_bits_data = GEN_30;
  assign GEN_3_ready = GEN_23;
  assign GEN_3_valid = GEN_24;
  assign GEN_3_bits_addr_beat = GEN_25;
  assign GEN_3_bits_client_xact_id = GEN_26;
  assign GEN_3_bits_manager_xact_id = GEN_27;
  assign GEN_3_bits_is_builtin_type = GEN_28;
  assign GEN_3_bits_g_type = GEN_29;
  assign GEN_3_bits_data = GEN_30;
  assign GEN_4_ready = GEN_23;
  assign GEN_4_valid = GEN_24;
  assign GEN_4_bits_addr_beat = GEN_25;
  assign GEN_4_bits_client_xact_id = GEN_26;
  assign GEN_4_bits_manager_xact_id = GEN_27;
  assign GEN_4_bits_is_builtin_type = GEN_28;
  assign GEN_4_bits_g_type = GEN_29;
  assign GEN_4_bits_data = GEN_30;
  assign GEN_5_ready = GEN_23;
  assign GEN_5_valid = GEN_24;
  assign GEN_5_bits_addr_beat = GEN_25;
  assign GEN_5_bits_client_xact_id = GEN_26;
  assign GEN_5_bits_manager_xact_id = GEN_27;
  assign GEN_5_bits_is_builtin_type = GEN_28;
  assign GEN_5_bits_g_type = GEN_29;
  assign GEN_5_bits_data = GEN_30;
  assign GEN_6_ready = GEN_23;
  assign GEN_6_valid = GEN_24;
  assign GEN_6_bits_addr_beat = GEN_25;
  assign GEN_6_bits_client_xact_id = GEN_26;
  assign GEN_6_bits_manager_xact_id = GEN_27;
  assign GEN_6_bits_is_builtin_type = GEN_28;
  assign GEN_6_bits_g_type = GEN_29;
  assign GEN_6_bits_data = GEN_30;
  assign T_798 = T_794 != 3'h0;
  assign T_806_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_806_0};
  assign T_808 = io_out_bits_g_type == GEN_0;
  assign T_809 = io_out_bits_g_type == 4'h0;
  assign T_810 = io_out_bits_is_builtin_type ? T_808 : T_809;
  assign T_812 = io_out_ready & io_out_valid;
  assign T_813 = T_812 & T_810;
  assign T_817 = T_794 + 3'h1;
  assign T_818 = T_817[2:0];
  assign GEN_175 = T_813 ? io_chosen : T_796;
  assign GEN_176 = T_813 ? T_818 : T_794;
  assign GEN_177 = T_798 ? T_796 : choice;
  assign GEN_178 = T_812 ? io_chosen : lastGrant;
  assign grantMask_1 = 2'h1 > lastGrant;
  assign grantMask_2 = 2'h2 > lastGrant;
  assign grantMask_3 = 2'h3 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign validMask_2 = io_in_2_valid & grantMask_2;
  assign validMask_3 = io_in_3_valid & grantMask_3;
  assign T_826 = validMask_1 | validMask_2;
  assign T_827 = T_826 | validMask_3;
  assign T_828 = T_827 | io_in_0_valid;
  assign T_829 = T_828 | io_in_1_valid;
  assign T_830 = T_829 | io_in_2_valid;
  assign T_834 = validMask_1 == 1'h0;
  assign T_836 = T_826 == 1'h0;
  assign T_838 = T_827 == 1'h0;
  assign T_840 = T_828 == 1'h0;
  assign T_842 = T_829 == 1'h0;
  assign T_844 = T_830 == 1'h0;
  assign T_848 = grantMask_1 | T_840;
  assign T_849 = T_834 & grantMask_2;
  assign T_850 = T_849 | T_842;
  assign T_851 = T_836 & grantMask_3;
  assign T_852 = T_851 | T_844;
  assign T_854 = T_796 == 2'h0;
  assign T_855 = T_798 ? T_854 : T_838;
  assign T_856 = T_855 & io_out_ready;
  assign T_858 = T_796 == 2'h1;
  assign T_859 = T_798 ? T_858 : T_848;
  assign T_860 = T_859 & io_out_ready;
  assign T_862 = T_796 == 2'h2;
  assign T_863 = T_798 ? T_862 : T_850;
  assign T_864 = T_863 & io_out_ready;
  assign T_866 = T_796 == 2'h3;
  assign T_867 = T_798 ? T_866 : T_852;
  assign T_868 = T_867 & io_out_ready;
  assign GEN_179 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_180 = io_in_1_valid ? 2'h1 : GEN_179;
  assign GEN_181 = io_in_0_valid ? 2'h0 : GEN_180;
  assign GEN_182 = validMask_3 ? 2'h3 : GEN_181;
  assign GEN_183 = validMask_2 ? 2'h2 : GEN_182;
  assign GEN_184 = validMask_1 ? 2'h1 : GEN_183;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_794 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_796 = GEN_2[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  lastGrant = GEN_3[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_794 <= 3'h0;
    end else begin
      if(T_813) begin
        T_794 <= T_818;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_813) begin
        T_796 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_812) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter_1(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [10:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire [2:0] T_1855_0;
  wire [2:0] T_1855_1;
  wire  T_1857;
  wire  T_1858;
  wire  T_1859;
  wire  T_1860;
  wire [2:0] T_1861;
  wire [2:0] T_1863;
  wire [28:0] T_1864;
  wire [31:0] T_1865;
  wire  T_1869;
  wire  T_1872;
  wire  T_1874;
  wire  T_1875;
  wire  T_1877;
  wire  T_1879;
  wire  T_1880;
  wire  T_1882;
  wire  T_1884;
  wire  T_1885;
  wire [1:0] T_1886;
  wire [1:0] T_1887;
  wire [3:0] acq_route;
  wire  T_1889;
  wire  T_1890;
  wire  GEN_0;
  wire  T_1892;
  wire  T_1893;
  wire  GEN_1;
  wire  T_1895;
  wire  T_1896;
  wire  GEN_2;
  wire  T_1898;
  wire  T_1899;
  wire  GEN_3;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_2_ready;
  wire  gnt_arb_io_in_2_valid;
  wire [2:0] gnt_arb_io_in_2_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_2_bits_client_xact_id;
  wire  gnt_arb_io_in_2_bits_manager_xact_id;
  wire  gnt_arb_io_in_2_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_2_bits_g_type;
  wire [63:0] gnt_arb_io_in_2_bits_data;
  wire  gnt_arb_io_in_3_ready;
  wire  gnt_arb_io_in_3_valid;
  wire [2:0] gnt_arb_io_in_3_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_3_bits_client_xact_id;
  wire  gnt_arb_io_in_3_bits_manager_xact_id;
  wire  gnt_arb_io_in_3_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_3_bits_g_type;
  wire [63:0] gnt_arb_io_in_3_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire [1:0] gnt_arb_io_chosen;
  wire  T_1924;
  wire  T_1926;
  wire  T_1927;
  wire  T_1928;
  wire  T_1930;
  LockingRRArbiter_11 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_2_ready(gnt_arb_io_in_2_ready),
    .io_in_2_valid(gnt_arb_io_in_2_valid),
    .io_in_2_bits_addr_beat(gnt_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(gnt_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(gnt_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(gnt_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(gnt_arb_io_in_2_bits_g_type),
    .io_in_2_bits_data(gnt_arb_io_in_2_bits_data),
    .io_in_3_ready(gnt_arb_io_in_3_ready),
    .io_in_3_valid(gnt_arb_io_in_3_valid),
    .io_in_3_bits_addr_beat(gnt_arb_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(gnt_arb_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(gnt_arb_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(gnt_arb_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(gnt_arb_io_in_3_bits_g_type),
    .io_in_3_bits_data(gnt_arb_io_in_3_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_3;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1890;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1893;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign io_out_2_acquire_valid = T_1896;
  assign io_out_2_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_2_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_2_grant_ready = gnt_arb_io_in_2_ready;
  assign io_out_3_acquire_valid = T_1899;
  assign io_out_3_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_3_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_3_grant_ready = gnt_arb_io_in_3_ready;
  assign T_1855_0 = 3'h0;
  assign T_1855_1 = 3'h4;
  assign T_1857 = io_in_acquire_bits_a_type == T_1855_0;
  assign T_1858 = io_in_acquire_bits_a_type == T_1855_1;
  assign T_1859 = T_1857 | T_1858;
  assign T_1860 = io_in_acquire_bits_is_builtin_type & T_1859;
  assign T_1861 = io_in_acquire_bits_union[10:8];
  assign T_1863 = T_1860 ? T_1861 : 3'h0;
  assign T_1864 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1865 = {T_1864,T_1863};
  assign T_1869 = T_1865 < 32'h1000;
  assign T_1872 = 32'h1000 <= T_1865;
  assign T_1874 = T_1865 < 32'h2000;
  assign T_1875 = T_1872 & T_1874;
  assign T_1877 = 32'h40000000 <= T_1865;
  assign T_1879 = T_1865 < 32'h44000000;
  assign T_1880 = T_1877 & T_1879;
  assign T_1882 = 32'h44000000 <= T_1865;
  assign T_1884 = T_1865 < 32'h48000000;
  assign T_1885 = T_1882 & T_1884;
  assign T_1886 = {T_1875,T_1869};
  assign T_1887 = {T_1885,T_1880};
  assign acq_route = {T_1887,T_1886};
  assign T_1889 = acq_route[0];
  assign T_1890 = io_in_acquire_valid & T_1889;
  assign GEN_0 = T_1889 ? io_out_0_acquire_ready : 1'h0;
  assign T_1892 = acq_route[1];
  assign T_1893 = io_in_acquire_valid & T_1892;
  assign GEN_1 = T_1892 ? io_out_1_acquire_ready : GEN_0;
  assign T_1895 = acq_route[2];
  assign T_1896 = io_in_acquire_valid & T_1895;
  assign GEN_2 = T_1895 ? io_out_2_acquire_ready : GEN_1;
  assign T_1898 = acq_route[3];
  assign T_1899 = io_in_acquire_valid & T_1898;
  assign GEN_3 = T_1898 ? io_out_3_acquire_ready : GEN_2;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_in_2_valid = io_out_2_grant_valid;
  assign gnt_arb_io_in_2_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign gnt_arb_io_in_2_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign gnt_arb_io_in_2_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_2_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_2_bits_g_type = io_out_2_grant_bits_g_type;
  assign gnt_arb_io_in_2_bits_data = io_out_2_grant_bits_data;
  assign gnt_arb_io_in_3_valid = io_out_3_grant_valid;
  assign gnt_arb_io_in_3_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign gnt_arb_io_in_3_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign gnt_arb_io_in_3_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_3_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_3_bits_g_type = io_out_3_grant_bits_g_type;
  assign gnt_arb_io_in_3_bits_data = io_out_3_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1924 = io_in_acquire_valid == 1'h0;
  assign T_1926 = acq_route != 4'h0;
  assign T_1927 = T_1924 | T_1926;
  assign T_1928 = T_1927 | reset;
  assign T_1930 = T_1928 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1930) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1930) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIORouter_1 ClientUncachedTileLinkIORouter_1_1 (
    .clk(ClientUncachedTileLinkIORouter_1_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [10:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [10:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [10:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  xbar_io_out_2_acquire_ready;
  wire  xbar_io_out_2_acquire_valid;
  wire [25:0] xbar_io_out_2_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_2_acquire_bits_addr_beat;
  wire  xbar_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_2_acquire_bits_a_type;
  wire [10:0] xbar_io_out_2_acquire_bits_union;
  wire [63:0] xbar_io_out_2_acquire_bits_data;
  wire  xbar_io_out_2_grant_ready;
  wire  xbar_io_out_2_grant_valid;
  wire [2:0] xbar_io_out_2_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_2_grant_bits_client_xact_id;
  wire  xbar_io_out_2_grant_bits_manager_xact_id;
  wire  xbar_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_2_grant_bits_g_type;
  wire [63:0] xbar_io_out_2_grant_bits_data;
  wire  xbar_io_out_3_acquire_ready;
  wire  xbar_io_out_3_acquire_valid;
  wire [25:0] xbar_io_out_3_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_3_acquire_bits_addr_beat;
  wire  xbar_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_3_acquire_bits_a_type;
  wire [10:0] xbar_io_out_3_acquire_bits_union;
  wire [63:0] xbar_io_out_3_acquire_bits_data;
  wire  xbar_io_out_3_grant_ready;
  wire  xbar_io_out_3_grant_valid;
  wire [2:0] xbar_io_out_3_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_3_grant_bits_client_xact_id;
  wire  xbar_io_out_3_grant_bits_manager_xact_id;
  wire  xbar_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_3_grant_bits_g_type;
  wire [63:0] xbar_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar_1 xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(xbar_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(xbar_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(xbar_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(xbar_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(xbar_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(xbar_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(xbar_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(xbar_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(xbar_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(xbar_io_out_2_grant_ready),
    .io_out_2_grant_valid(xbar_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(xbar_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(xbar_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(xbar_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(xbar_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(xbar_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(xbar_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(xbar_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(xbar_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(xbar_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(xbar_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(xbar_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(xbar_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(xbar_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(xbar_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(xbar_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(xbar_io_out_3_grant_ready),
    .io_out_3_grant_valid(xbar_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(xbar_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(xbar_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(xbar_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(xbar_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(xbar_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(xbar_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = xbar_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = xbar_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = xbar_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = xbar_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = xbar_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = xbar_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = xbar_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = xbar_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = xbar_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = xbar_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = xbar_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = xbar_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = xbar_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = xbar_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = xbar_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = xbar_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = xbar_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = xbar_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = xbar_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = xbar_io_out_3_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = io_out_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_1_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign xbar_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign xbar_io_out_2_grant_valid = io_out_2_grant_valid;
  assign xbar_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign xbar_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign xbar_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign xbar_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign xbar_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign xbar_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign xbar_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign xbar_io_out_3_grant_valid = io_out_3_grant_valid;
  assign xbar_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign xbar_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign xbar_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign xbar_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign xbar_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign xbar_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [10:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [10:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [10:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [10:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [10:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [10:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [10:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_clk;
  wire  TileLinkRecursiveInterconnect_1_1_reset;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data)
  );
  TileLinkRecursiveInterconnect_1 TileLinkRecursiveInterconnect_1_1 (
    .clk(TileLinkRecursiveInterconnect_1_1_clk),
    .reset(TileLinkRecursiveInterconnect_1_1_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_clk = clk;
  assign TileLinkRecursiveInterconnect_1_1_reset = reset;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready = xbar_io_out_0_grant_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module Queue_16(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [10:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [10:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_254_data;
  wire  ram_addr_block_T_254_addr;
  wire  ram_addr_block_T_254_en;
  wire [25:0] ram_addr_block_T_224_data;
  wire  ram_addr_block_T_224_addr;
  wire  ram_addr_block_T_224_mask;
  wire  ram_addr_block_T_224_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_254_data;
  wire  ram_client_xact_id_T_254_addr;
  wire  ram_client_xact_id_T_254_en;
  wire [1:0] ram_client_xact_id_T_224_data;
  wire  ram_client_xact_id_T_224_addr;
  wire  ram_client_xact_id_T_224_mask;
  wire  ram_client_xact_id_T_224_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_254_data;
  wire  ram_addr_beat_T_254_addr;
  wire  ram_addr_beat_T_254_en;
  wire [2:0] ram_addr_beat_T_224_data;
  wire  ram_addr_beat_T_224_addr;
  wire  ram_addr_beat_T_224_mask;
  wire  ram_addr_beat_T_224_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_254_data;
  wire  ram_is_builtin_type_T_254_addr;
  wire  ram_is_builtin_type_T_254_en;
  wire  ram_is_builtin_type_T_224_data;
  wire  ram_is_builtin_type_T_224_addr;
  wire  ram_is_builtin_type_T_224_mask;
  wire  ram_is_builtin_type_T_224_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_254_data;
  wire  ram_a_type_T_254_addr;
  wire  ram_a_type_T_254_en;
  wire [2:0] ram_a_type_T_224_data;
  wire  ram_a_type_T_224_addr;
  wire  ram_a_type_T_224_mask;
  wire  ram_a_type_T_224_en;
  reg [10:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [10:0] ram_union_T_254_data;
  wire  ram_union_T_254_addr;
  wire  ram_union_T_254_en;
  wire [10:0] ram_union_T_224_data;
  wire  ram_union_T_224_addr;
  wire  ram_union_T_224_mask;
  wire  ram_union_T_224_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_254_data;
  wire  ram_data_T_254_addr;
  wire  ram_data_T_254_en;
  wire [63:0] ram_data_T_224_data;
  wire  ram_data_T_224_addr;
  wire  ram_data_T_224_mask;
  wire  ram_data_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_17;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_addr_block = ram_addr_block_T_254_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_254_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_254_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_254_data;
  assign io_deq_bits_a_type = ram_a_type_T_254_data;
  assign io_deq_bits_union = ram_union_T_254_data;
  assign io_deq_bits_data = ram_data_T_254_data;
  assign io_count = T_279[0];
  assign ram_addr_block_T_254_addr = 1'h0;
  assign ram_addr_block_T_254_en = 1'h1;
  assign ram_addr_block_T_254_data = ram_addr_block[ram_addr_block_T_254_addr];
  assign ram_addr_block_T_224_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_224_addr = 1'h0;
  assign ram_addr_block_T_224_mask = do_enq;
  assign ram_addr_block_T_224_en = do_enq;
  assign ram_client_xact_id_T_254_addr = 1'h0;
  assign ram_client_xact_id_T_254_en = 1'h1;
  assign ram_client_xact_id_T_254_data = ram_client_xact_id[ram_client_xact_id_T_254_addr];
  assign ram_client_xact_id_T_224_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_224_addr = 1'h0;
  assign ram_client_xact_id_T_224_mask = do_enq;
  assign ram_client_xact_id_T_224_en = do_enq;
  assign ram_addr_beat_T_254_addr = 1'h0;
  assign ram_addr_beat_T_254_en = 1'h1;
  assign ram_addr_beat_T_254_data = ram_addr_beat[ram_addr_beat_T_254_addr];
  assign ram_addr_beat_T_224_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_224_addr = 1'h0;
  assign ram_addr_beat_T_224_mask = do_enq;
  assign ram_addr_beat_T_224_en = do_enq;
  assign ram_is_builtin_type_T_254_addr = 1'h0;
  assign ram_is_builtin_type_T_254_en = 1'h1;
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  assign ram_is_builtin_type_T_224_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_224_addr = 1'h0;
  assign ram_is_builtin_type_T_224_mask = do_enq;
  assign ram_is_builtin_type_T_224_en = do_enq;
  assign ram_a_type_T_254_addr = 1'h0;
  assign ram_a_type_T_254_en = 1'h1;
  assign ram_a_type_T_254_data = ram_a_type[ram_a_type_T_254_addr];
  assign ram_a_type_T_224_data = io_enq_bits_a_type;
  assign ram_a_type_T_224_addr = 1'h0;
  assign ram_a_type_T_224_mask = do_enq;
  assign ram_a_type_T_224_en = do_enq;
  assign ram_union_T_254_addr = 1'h0;
  assign ram_union_T_254_en = 1'h1;
  assign ram_union_T_254_data = ram_union[ram_union_T_254_addr];
  assign ram_union_T_224_data = io_enq_bits_union;
  assign ram_union_T_224_addr = 1'h0;
  assign ram_union_T_224_mask = do_enq;
  assign ram_union_T_224_en = do_enq;
  assign ram_data_T_254_addr = 1'h0;
  assign ram_data_T_254_en = 1'h1;
  assign ram_data_T_254_data = ram_data[ram_data_T_254_addr];
  assign ram_data_T_224_data = io_enq_bits_data;
  assign ram_data_T_224_addr = 1'h0;
  assign ram_data_T_224_mask = do_enq;
  assign ram_data_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_17 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[10:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_224_en & ram_addr_block_T_224_mask) begin
      ram_addr_block[ram_addr_block_T_224_addr] <= ram_addr_block_T_224_data;
    end
    if(ram_client_xact_id_T_224_en & ram_client_xact_id_T_224_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_224_addr] <= ram_client_xact_id_T_224_data;
    end
    if(ram_addr_beat_T_224_en & ram_addr_beat_T_224_mask) begin
      ram_addr_beat[ram_addr_beat_T_224_addr] <= ram_addr_beat_T_224_data;
    end
    if(ram_is_builtin_type_T_224_en & ram_is_builtin_type_T_224_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_224_addr] <= ram_is_builtin_type_T_224_data;
    end
    if(ram_a_type_T_224_en & ram_a_type_T_224_mask) begin
      ram_a_type[ram_a_type_T_224_addr] <= ram_a_type_T_224_data;
    end
    if(ram_union_T_224_en & ram_union_T_224_mask) begin
      ram_union[ram_union_T_224_addr] <= ram_union_T_224_data;
    end
    if(ram_data_T_224_en & ram_data_T_224_mask) begin
      ram_data[ram_data_T_224_addr] <= ram_data_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  output  io_harts_0,
  output  io_harts_1,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_477_0;
  wire  T_477_1;
  wire  T_477_2;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  T_489_0;
  wire  T_489_1;
  wire  threshold_0;
  wire  threshold_1;
  wire  T_502_0;
  wire  T_502_1;
  wire  T_502_2;
  reg  pending_0;
  reg [31:0] GEN_8;
  reg  pending_1;
  reg [31:0] GEN_16;
  reg  pending_2;
  reg [31:0] GEN_17;
  reg  enables_0_0;
  reg [31:0] GEN_20;
  reg  enables_0_1;
  reg [31:0] GEN_21;
  reg  enables_0_2;
  reg [31:0] GEN_22;
  reg  enables_1_0;
  reg [31:0] GEN_32;
  reg  enables_1_1;
  reg [31:0] GEN_35;
  reg  enables_1_2;
  reg [31:0] GEN_36;
  wire  T_545;
  wire  GEN_12;
  wire  T_549;
  wire  GEN_13;
  wire [1:0] maxDevs_0;
  wire [1:0] maxDevs_1;
  wire  T_559;
  wire [1:0] T_560;
  wire  T_561;
  wire [1:0] T_562;
  wire  T_567;
  wire [1:0] T_568;
  wire [1:0] T_570;
  wire  T_571;
  wire  T_572;
  wire  T_574;
  wire [1:0] T_575;
  wire [2:0] T_577;
  wire [1:0] T_578;
  wire [1:0] T_579;
  reg [1:0] T_580;
  reg [31:0] GEN_39;
  reg [1:0] T_581;
  reg [31:0] GEN_40;
  wire [1:0] T_583;
  wire  T_584;
  wire  T_585;
  wire [1:0] T_586;
  wire  T_587;
  wire [1:0] T_588;
  wire  T_593;
  wire [1:0] T_594;
  wire  T_598;
  wire  T_600;
  wire [1:0] T_601;
  wire [1:0] T_605;
  reg [1:0] T_606;
  reg [31:0] GEN_43;
  reg [1:0] T_607;
  reg [31:0] GEN_44;
  wire [1:0] T_609;
  wire  T_610;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_634;
  wire  T_636;
  wire  T_637;
  wire  read;
  wire  T_640;
  wire  T_641;
  wire  write;
  wire  T_644;
  wire  T_645;
  wire  T_646;
  wire  T_647;
  wire  T_649;
  wire [2:0] T_657_0;
  wire [2:0] T_657_1;
  wire  T_659;
  wire  T_660;
  wire  T_661;
  wire  T_662;
  wire [2:0] T_663;
  wire [2:0] T_665;
  wire [28:0] T_666;
  wire [31:0] T_667;
  wire [25:0] addr;
  wire [26:0] T_669;
  wire [25:0] T_670;
  wire  claimant;
  wire  hart;
  wire [63:0] rdata;
  wire  T_676;
  wire  T_677;
  wire  T_696;
  wire  T_697;
  wire  T_701;
  wire [7:0] T_702;
  wire [7:0] T_704;
  wire [7:0] T_705;
  wire  T_706;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  T_710;
  wire  T_711;
  wire  T_712;
  wire  T_713;
  wire [7:0] T_717;
  wire [7:0] T_721;
  wire [7:0] T_725;
  wire [7:0] T_729;
  wire [7:0] T_733;
  wire [7:0] T_737;
  wire [7:0] T_741;
  wire [7:0] T_745;
  wire [15:0] T_746;
  wire [15:0] T_747;
  wire [31:0] T_748;
  wire [15:0] T_749;
  wire [15:0] T_750;
  wire [31:0] T_751;
  wire [63:0] T_752;
  wire [63:0] T_753;
  wire [63:0] T_832;
  wire [63:0] T_833;
  wire [63:0] masked_wdata;
  wire  T_835;
  wire [1:0] GEN_0;
  wire [1:0] GEN_14;
  wire [32:0] T_838;
  wire  GEN_1;
  wire  GEN_15;
  wire [33:0] T_839;
  wire [7:0] T_841;
  wire [33:0] T_842;
  wire  T_843;
  wire  T_844;
  wire [1:0] GEN_2;
  wire  GEN_3;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_23;
  wire  GEN_24;
  wire [31:0] T_878;
  wire [1:0] T_879;
  wire  GEN_4;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_25;
  wire  GEN_122;
  wire  GEN_26;
  wire  GEN_123;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [2:0] T_881;
  wire [1:0] T_882;
  wire  GEN_5;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_41;
  wire  GEN_42;
  wire [63:0] GEN_45;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_53;
  wire  GEN_54;
  wire  T_890;
  wire  T_892;
  wire  T_893;
  wire [26:0] T_895;
  wire [25:0] T_896;
  wire  T_897;
  wire  GEN_6_0;
  wire  GEN_6_1;
  wire  GEN_6_2;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_7_0;
  wire  GEN_7_1;
  wire  GEN_7_2;
  wire [1:0] T_901;
  wire  GEN_8_0;
  wire  GEN_8_1;
  wire  GEN_8_2;
  wire [2:0] T_902;
  wire  T_906;
  wire  GEN_9;
  wire  T_910;
  wire  GEN_10;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_72;
  wire  GEN_73;
  wire  T_914;
  wire  GEN_11;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_77;
  wire  GEN_78;
  wire [63:0] GEN_88;
  wire  GEN_98;
  wire [63:0] GEN_108;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_116;
  wire  GEN_117;
  wire  T_916;
  wire  T_920;
  wire  T_921;
  wire  T_922;
  wire [1:0] T_924;
  wire [2:0] T_925;
  wire [2:0] T_928;
  wire [63:0] GEN_118;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_939;
  wire [31:0] T_941;
  wire [31:0] T_943;
  wire [63:0] T_944;
  wire [63:0] GEN_119;
  wire [31:0] T_948;
  wire [63:0] GEN_120;
  wire [63:0] GEN_121;
  wire  T_969;
  wire [2:0] T_970;
  wire  T_971;
  wire [2:0] T_972;
  wire  T_973;
  wire [2:0] T_974;
  wire  T_975;
  wire [2:0] T_976;
  wire  T_977;
  wire [2:0] T_978;
  wire  T_979;
  wire [2:0] T_980;
  wire  T_981;
  wire [2:0] T_982;
  wire [2:0] T_1007_addr_beat;
  wire [1:0] T_1007_client_xact_id;
  wire  T_1007_manager_xact_id;
  wire  T_1007_is_builtin_type;
  wire [3:0] T_1007_g_type;
  wire [63:0] T_1007_data;
  Queue_16 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_545;
  assign io_devices_0_complete = GEN_53;
  assign io_devices_1_ready = T_549;
  assign io_devices_1_complete = GEN_54;
  assign io_harts_0 = T_584;
  assign io_harts_1 = T_610;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_1007_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1007_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1007_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1007_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1007_g_type;
  assign io_tl_grant_bits_data = T_1007_data;
  assign T_477_0 = 1'h1;
  assign T_477_1 = 1'h1;
  assign T_477_2 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_477_1;
  assign priority_2 = T_477_2;
  assign T_489_0 = 1'h0;
  assign T_489_1 = 1'h0;
  assign threshold_0 = T_489_0;
  assign threshold_1 = T_489_1;
  assign T_502_0 = 1'h0;
  assign T_502_1 = 1'h0;
  assign T_502_2 = 1'h0;
  assign T_545 = pending_1 == 1'h0;
  assign GEN_12 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_549 = pending_2 == 1'h0;
  assign GEN_13 = io_devices_1_valid ? 1'h1 : pending_2;
  assign maxDevs_0 = T_580;
  assign maxDevs_1 = T_606;
  assign T_559 = pending_1 & enables_0_1;
  assign T_560 = {T_559,priority_1};
  assign T_561 = pending_2 & enables_0_2;
  assign T_562 = {T_561,priority_2};
  assign T_567 = 2'h2 >= T_560;
  assign T_568 = T_567 ? 2'h2 : T_560;
  assign T_570 = 1'h1 + 1'h0;
  assign T_571 = T_570[0:0];
  assign T_572 = T_567 ? 1'h0 : T_571;
  assign T_574 = T_568 >= T_562;
  assign T_575 = T_574 ? T_568 : T_562;
  assign T_577 = 2'h2 + 2'h0;
  assign T_578 = T_577[1:0];
  assign T_579 = T_574 ? {{1'd0}, T_572} : T_578;
  assign T_583 = {1'h1,threshold_0};
  assign T_584 = T_581 > T_583;
  assign T_585 = pending_1 & enables_1_1;
  assign T_586 = {T_585,priority_1};
  assign T_587 = pending_2 & enables_1_2;
  assign T_588 = {T_587,priority_2};
  assign T_593 = 2'h2 >= T_586;
  assign T_594 = T_593 ? 2'h2 : T_586;
  assign T_598 = T_593 ? 1'h0 : T_571;
  assign T_600 = T_594 >= T_588;
  assign T_601 = T_600 ? T_594 : T_588;
  assign T_605 = T_600 ? {{1'd0}, T_598} : T_578;
  assign T_609 = {1'h1,threshold_1};
  assign T_610 = T_607 > T_609;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_634 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_636 = acq_io_deq_bits_a_type == 3'h0;
  assign T_637 = acq_io_deq_bits_is_builtin_type & T_636;
  assign read = T_634 & T_637;
  assign T_640 = acq_io_deq_bits_a_type == 3'h2;
  assign T_641 = acq_io_deq_bits_is_builtin_type & T_640;
  assign write = T_634 & T_641;
  assign T_644 = T_634 == 1'h0;
  assign T_645 = T_644 | read;
  assign T_646 = T_645 | write;
  assign T_647 = T_646 | reset;
  assign T_649 = T_647 == 1'h0;
  assign T_657_0 = 3'h0;
  assign T_657_1 = 3'h4;
  assign T_659 = acq_io_deq_bits_a_type == T_657_0;
  assign T_660 = acq_io_deq_bits_a_type == T_657_1;
  assign T_661 = T_659 | T_660;
  assign T_662 = acq_io_deq_bits_is_builtin_type & T_661;
  assign T_663 = acq_io_deq_bits_union[10:8];
  assign T_665 = T_662 ? T_663 : 3'h0;
  assign T_666 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_667 = {T_666,T_665};
  assign addr = T_667[25:0];
  assign T_669 = addr - 26'h200000;
  assign T_670 = T_669[25:0];
  assign claimant = T_670[12];
  assign hart = GEN_98;
  assign rdata = GEN_121;
  assign T_676 = acq_io_deq_bits_a_type == 3'h4;
  assign T_677 = acq_io_deq_bits_is_builtin_type & T_676;
  assign T_696 = acq_io_deq_bits_a_type == 3'h3;
  assign T_697 = acq_io_deq_bits_is_builtin_type & T_696;
  assign T_701 = T_697 | T_641;
  assign T_702 = acq_io_deq_bits_union[8:1];
  assign T_704 = T_701 ? T_702 : 8'h0;
  assign T_705 = T_677 ? 8'hff : T_704;
  assign T_706 = T_705[0];
  assign T_707 = T_705[1];
  assign T_708 = T_705[2];
  assign T_709 = T_705[3];
  assign T_710 = T_705[4];
  assign T_711 = T_705[5];
  assign T_712 = T_705[6];
  assign T_713 = T_705[7];
  assign T_717 = T_706 ? 8'hff : 8'h0;
  assign T_721 = T_707 ? 8'hff : 8'h0;
  assign T_725 = T_708 ? 8'hff : 8'h0;
  assign T_729 = T_709 ? 8'hff : 8'h0;
  assign T_733 = T_710 ? 8'hff : 8'h0;
  assign T_737 = T_711 ? 8'hff : 8'h0;
  assign T_741 = T_712 ? 8'hff : 8'h0;
  assign T_745 = T_713 ? 8'hff : 8'h0;
  assign T_746 = {T_721,T_717};
  assign T_747 = {T_729,T_725};
  assign T_748 = {T_747,T_746};
  assign T_749 = {T_737,T_733};
  assign T_750 = {T_745,T_741};
  assign T_751 = {T_750,T_749};
  assign T_752 = {T_751,T_748};
  assign T_753 = acq_io_deq_bits_data & T_752;
  assign T_832 = ~ T_752;
  assign T_833 = rdata & T_832;
  assign masked_wdata = T_753 | T_833;
  assign T_835 = addr >= 26'h200000;
  assign GEN_0 = GEN_14;
  assign GEN_14 = claimant ? maxDevs_1 : maxDevs_0;
  assign T_838 = {GEN_0,31'h0};
  assign GEN_1 = GEN_15;
  assign GEN_15 = claimant ? threshold_1 : threshold_0;
  assign T_839 = {T_838,GEN_1};
  assign T_841 = 7'h0 * 7'h40;
  assign T_842 = T_839 >> T_841;
  assign T_843 = addr[2];
  assign T_844 = read & T_843;
  assign GEN_2 = GEN_14;
  assign GEN_3 = 1'h0;
  assign GEN_18 = 2'h1 == GEN_2 ? GEN_3 : GEN_12;
  assign GEN_19 = 2'h2 == GEN_2 ? GEN_3 : GEN_13;
  assign GEN_23 = T_844 ? GEN_18 : GEN_12;
  assign GEN_24 = T_844 ? GEN_19 : GEN_13;
  assign T_878 = acq_io_deq_bits_data[63:32];
  assign T_879 = T_878[1:0];
  assign GEN_4 = GEN_29;
  assign GEN_6 = 1'h0 == hart;
  assign GEN_7 = 2'h1 == T_879;
  assign GEN_25 = GEN_6 & GEN_7 ? enables_0_1 : enables_0_0;
  assign GEN_122 = 2'h2 == T_879;
  assign GEN_26 = GEN_6 & GEN_122 ? enables_0_2 : GEN_25;
  assign GEN_123 = 2'h0 == T_879;
  assign GEN_27 = hart & GEN_123 ? enables_1_0 : GEN_26;
  assign GEN_28 = hart & GEN_7 ? enables_1_1 : GEN_27;
  assign GEN_29 = hart & GEN_122 ? enables_1_2 : GEN_28;
  assign T_881 = T_879 - 2'h1;
  assign T_882 = T_881[1:0];
  assign GEN_5 = 1'h1;
  assign GEN_30 = 2'h0 == T_882 ? GEN_5 : 1'h0;
  assign GEN_31 = 2'h1 == T_882 ? GEN_5 : 1'h0;
  assign GEN_33 = GEN_4 ? GEN_30 : 1'h0;
  assign GEN_34 = GEN_4 ? GEN_31 : 1'h0;
  assign GEN_37 = T_710 ? GEN_33 : 1'h0;
  assign GEN_38 = T_710 ? GEN_34 : 1'h0;
  assign GEN_41 = write ? GEN_37 : 1'h0;
  assign GEN_42 = write ? GEN_38 : 1'h0;
  assign GEN_45 = T_835 ? {{30'd0}, T_842} : 64'h0;
  assign GEN_49 = T_835 ? GEN_23 : GEN_12;
  assign GEN_50 = T_835 ? GEN_24 : GEN_13;
  assign GEN_53 = T_835 ? GEN_41 : 1'h0;
  assign GEN_54 = T_835 ? GEN_42 : 1'h0;
  assign T_890 = addr >= 26'h2000;
  assign T_892 = T_835 == 1'h0;
  assign T_893 = T_892 & T_890;
  assign T_895 = addr - 26'h2000;
  assign T_896 = T_895[25:0];
  assign T_897 = T_896[7];
  assign GEN_6_0 = GEN_55;
  assign GEN_6_1 = GEN_56;
  assign GEN_6_2 = GEN_57;
  assign GEN_55 = hart ? enables_1_0 : enables_0_0;
  assign GEN_56 = hart ? enables_1_1 : enables_0_1;
  assign GEN_57 = hart ? enables_1_2 : enables_0_2;
  assign GEN_7_0 = GEN_55;
  assign GEN_7_1 = GEN_56;
  assign GEN_7_2 = GEN_57;
  assign T_901 = {GEN_6_2,GEN_7_1};
  assign GEN_8_0 = GEN_55;
  assign GEN_8_1 = GEN_56;
  assign GEN_8_2 = GEN_57;
  assign T_902 = {T_901,GEN_8_0};
  assign T_906 = masked_wdata[0];
  assign GEN_9 = T_906;
  assign T_910 = masked_wdata[1];
  assign GEN_10 = T_910;
  assign GEN_69 = 1'h0 == T_897 ? GEN_10 : enables_0_1;
  assign GEN_70 = T_897 ? GEN_10 : enables_1_1;
  assign GEN_72 = write ? GEN_69 : enables_0_1;
  assign GEN_73 = write ? GEN_70 : enables_1_1;
  assign T_914 = masked_wdata[2];
  assign GEN_11 = T_914;
  assign GEN_74 = 1'h0 == T_897 ? GEN_11 : enables_0_2;
  assign GEN_75 = T_897 ? GEN_11 : enables_1_2;
  assign GEN_77 = write ? GEN_74 : enables_0_2;
  assign GEN_78 = write ? GEN_75 : enables_1_2;
  assign GEN_88 = {{61'd0}, T_902};
  assign GEN_98 = T_893 ? T_897 : claimant;
  assign GEN_108 = T_893 ? GEN_88 : GEN_45;
  assign GEN_113 = T_893 ? GEN_72 : enables_0_1;
  assign GEN_114 = T_893 ? GEN_73 : enables_1_1;
  assign GEN_116 = T_893 ? GEN_77 : enables_0_2;
  assign GEN_117 = T_893 ? GEN_78 : enables_1_2;
  assign T_916 = addr >= 26'h1000;
  assign T_920 = T_890 == 1'h0;
  assign T_921 = T_892 & T_920;
  assign T_922 = T_921 & T_916;
  assign T_924 = {pending_2,pending_1};
  assign T_925 = {T_924,pending_0};
  assign T_928 = T_925 >> T_841;
  assign GEN_118 = T_922 ? {{61'd0}, T_928} : GEN_108;
  assign T_935 = T_916 == 1'h0;
  assign T_936 = T_921 & T_935;
  assign T_937 = addr[3];
  assign T_939 = T_937 == 1'h0;
  assign T_941 = {31'h0,priority_0};
  assign T_943 = {31'h0,priority_1};
  assign T_944 = {T_943,T_941};
  assign GEN_119 = T_939 ? T_944 : GEN_118;
  assign T_948 = {31'h0,priority_2};
  assign GEN_120 = T_937 ? {{32'd0}, T_948} : GEN_119;
  assign GEN_121 = T_936 ? GEN_120 : GEN_118;
  assign T_969 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_970 = T_969 ? 3'h1 : 3'h3;
  assign T_971 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_972 = T_971 ? 3'h1 : T_970;
  assign T_973 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_974 = T_973 ? 3'h4 : T_972;
  assign T_975 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_976 = T_975 ? 3'h3 : T_974;
  assign T_977 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_978 = T_977 ? 3'h3 : T_976;
  assign T_979 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_980 = T_979 ? 3'h5 : T_978;
  assign T_981 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_982 = T_981 ? 3'h4 : T_980;
  assign T_1007_addr_beat = 3'h0;
  assign T_1007_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_1007_manager_xact_id = 1'h0;
  assign T_1007_is_builtin_type = 1'h1;
  assign T_1007_g_type = {{1'd0}, T_982};
  assign T_1007_data = rdata;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_8 = {1{$random}};
  pending_0 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_16 = {1{$random}};
  pending_1 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_17 = {1{$random}};
  pending_2 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_20 = {1{$random}};
  enables_0_0 = GEN_20[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_21 = {1{$random}};
  enables_0_1 = GEN_21[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_22 = {1{$random}};
  enables_0_2 = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  enables_1_0 = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_35 = {1{$random}};
  enables_1_1 = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_36 = {1{$random}};
  enables_1_2 = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_39 = {1{$random}};
  T_580 = GEN_39[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_40 = {1{$random}};
  T_581 = GEN_40[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_43 = {1{$random}};
  T_606 = GEN_43[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_44 = {1{$random}};
  T_607 = GEN_44[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_502_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_502_1;
    end else begin
      if(T_835) begin
        if(T_844) begin
          if(2'h1 == GEN_2) begin
            pending_1 <= GEN_3;
          end else begin
            if(io_devices_0_valid) begin
              pending_1 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_2 <= T_502_2;
    end else begin
      if(T_835) begin
        if(T_844) begin
          if(2'h2 == GEN_2) begin
            pending_2 <= GEN_3;
          end else begin
            if(io_devices_1_valid) begin
              pending_2 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_893) begin
        if(write) begin
          if(1'h0 == T_897) begin
            enables_0_1 <= GEN_10;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_893) begin
        if(write) begin
          if(1'h0 == T_897) begin
            enables_0_2 <= GEN_11;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_1_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_893) begin
        if(write) begin
          if(T_897) begin
            enables_1_1 <= GEN_10;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_893) begin
        if(write) begin
          if(T_897) begin
            enables_1_2 <= GEN_11;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_574) begin
        T_580 <= {{1'd0}, T_572};
      end else begin
        T_580 <= T_578;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_574) begin
        if(T_567) begin
          T_581 <= 2'h2;
        end else begin
          T_581 <= T_560;
        end
      end else begin
        T_581 <= T_562;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_600) begin
        T_606 <= {{1'd0}, T_598};
      end else begin
        T_606 <= T_578;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_600) begin
        if(T_593) begin
          T_607 <= 2'h2;
        end else begin
          T_607 <= T_586;
        end
      end else begin
        T_607 <= T_588;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_649) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at Plic.scala:108 assert(!acq.fire() || read || write, \"unsupported PLIC operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_649) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LevelGateway(
  input   clk,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] GEN_2;
  wire  T_6;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_10;
  wire  T_11;
  assign io_plic_valid = T_11;
  assign T_6 = io_interrupt & io_plic_ready;
  assign GEN_0 = T_6 ? 1'h1 : inFlight;
  assign GEN_1 = io_plic_complete ? 1'h0 : GEN_0;
  assign T_10 = inFlight == 1'h0;
  assign T_11 = io_interrupt & T_10;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  inFlight = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      inFlight <= 1'h0;
    end else begin
      if(io_plic_complete) begin
        inFlight <= 1'h0;
      end else begin
        if(T_6) begin
          inFlight <= 1'h1;
        end
      end
    end
  end
endmodule
module DebugModule(
  input   clk,
  input   reset,
  output  io_db_req_ready,
  input   io_db_req_valid,
  input  [4:0] io_db_req_bits_addr,
  input  [33:0] io_db_req_bits_data,
  input  [1:0] io_db_req_bits_op,
  input   io_db_resp_ready,
  output  io_db_resp_valid,
  output [33:0] io_db_resp_bits_data,
  output [1:0] io_db_resp_bits_resp,
  output  io_debugInterrupts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_ndreset,
  output  io_fullreset
);
  wire  CONTROLReset_interrupt;
  wire  CONTROLReset_haltnot;
  wire [9:0] CONTROLReset_reserved0;
  wire [2:0] CONTROLReset_buserror;
  wire [2:0] CONTROLReset_serial;
  wire  CONTROLReset_autoincrement;
  wire [2:0] CONTROLReset_access;
  wire [9:0] CONTROLReset_hartid;
  wire  CONTROLReset_ndreset;
  wire  CONTROLReset_fullreset;
  wire  CONTROLWrEn;
  reg  CONTROLReg_interrupt;
  reg [31:0] GEN_26;
  reg  CONTROLReg_haltnot;
  reg [31:0] GEN_27;
  reg [9:0] CONTROLReg_reserved0;
  reg [31:0] GEN_28;
  reg [2:0] CONTROLReg_buserror;
  reg [31:0] GEN_29;
  reg [2:0] CONTROLReg_serial;
  reg [31:0] GEN_30;
  reg  CONTROLReg_autoincrement;
  reg [31:0] GEN_52;
  reg [2:0] CONTROLReg_access;
  reg [31:0] GEN_85;
  reg [9:0] CONTROLReg_hartid;
  reg [31:0] GEN_86;
  reg  CONTROLReg_ndreset;
  reg [31:0] GEN_88;
  reg  CONTROLReg_fullreset;
  reg [31:0] GEN_89;
  wire  CONTROLWrData_interrupt;
  wire  CONTROLWrData_haltnot;
  wire [9:0] CONTROLWrData_reserved0;
  wire [2:0] CONTROLWrData_buserror;
  wire [2:0] CONTROLWrData_serial;
  wire  CONTROLWrData_autoincrement;
  wire [2:0] CONTROLWrData_access;
  wire [9:0] CONTROLWrData_hartid;
  wire  CONTROLWrData_ndreset;
  wire  CONTROLWrData_fullreset;
  wire  CONTROLRdData_interrupt;
  wire  CONTROLRdData_haltnot;
  wire [9:0] CONTROLRdData_reserved0;
  wire [2:0] CONTROLRdData_buserror;
  wire [2:0] CONTROLRdData_serial;
  wire  CONTROLRdData_autoincrement;
  wire [2:0] CONTROLRdData_access;
  wire [9:0] CONTROLRdData_hartid;
  wire  CONTROLRdData_ndreset;
  wire  CONTROLRdData_fullreset;
  reg  ndresetCtrReg;
  reg [31:0] GEN_90;
  wire [1:0] DMINFORdData_reserved0;
  wire [6:0] DMINFORdData_abussize;
  wire [3:0] DMINFORdData_serialcount;
  wire  DMINFORdData_access128;
  wire  DMINFORdData_access64;
  wire  DMINFORdData_access32;
  wire  DMINFORdData_access16;
  wire  DMINFORdData_accesss8;
  wire [5:0] DMINFORdData_dramsize;
  wire  DMINFORdData_haltsum;
  wire [2:0] DMINFORdData_reserved1;
  wire  DMINFORdData_authenticated;
  wire  DMINFORdData_authbusy;
  wire [1:0] DMINFORdData_authtype;
  wire [1:0] DMINFORdData_version;
  wire  HALTSUMRdData_serialfull;
  wire  HALTSUMRdData_serialvalid;
  wire [31:0] HALTSUMRdData_acks;
  wire  RAMWrData_interrupt;
  wire  RAMWrData_haltnot;
  wire [31:0] RAMWrData_data;
  wire  RAMRdData_interrupt;
  wire  RAMRdData_haltnot;
  wire [31:0] RAMRdData_data;
  wire  SETHALTNOTWrEn;
  wire [9:0] SETHALTNOTWrData;
  wire  CLEARDEBINTWrEn;
  wire [9:0] CLEARDEBINTWrData;
  wire  T_655_0;
  reg  interruptRegs_0;
  reg [31:0] GEN_109;
  wire  T_666_0;
  reg  haltnotRegs_0;
  reg [31:0] GEN_110;
  wire [31:0] haltnotStatus_0;
  wire [31:0] rdHaltnotStatus;
  wire  haltnotSummary;
  reg [63:0] ramMem [0:7];
  reg [63:0] GEN_111;
  wire [63:0] ramMem_T_850_data;
  wire [2:0] ramMem_T_850_addr;
  wire  ramMem_T_850_en;
  wire [63:0] ramMem_T_851_data;
  wire [2:0] ramMem_T_851_addr;
  wire  ramMem_T_851_mask;
  wire  ramMem_T_851_en;
  wire [2:0] ramAddr;
  wire [63:0] ramRdData;
  wire [63:0] ramWrData;
  wire [63:0] ramWrMask;
  wire  ramWrEn;
  wire [3:0] dbRamAddr;
  wire [31:0] dbRamRdData;
  wire [31:0] dbRamWrData;
  wire  dbRamWrEn;
  wire  dbRamRdEn;
  wire [2:0] sbRamAddr;
  wire [63:0] sbRamRdData;
  wire [63:0] sbRamWrData;
  wire  sbRamWrEn;
  wire  sbRamRdEn;
  wire [63:0] sbRomRdData;
  wire  dbRdEn;
  wire  dbWrEn;
  wire [33:0] dbRdData;
  reg  dbStateReg;
  reg [31:0] GEN_112;
  wire [33:0] dbResult_data;
  wire [1:0] dbResult_resp;
  wire [4:0] dbReq_addr;
  wire [33:0] dbReq_data;
  wire [1:0] dbReq_op;
  reg [33:0] dbRespReg_data;
  reg [63:0] GEN_113;
  reg [1:0] dbRespReg_resp;
  reg [31:0] GEN_114;
  wire  rdCondWrFailure;
  wire  dbWrNeeded;
  wire [11:0] sbAddr;
  wire [63:0] sbRdData;
  wire [63:0] sbWrData;
  wire [63:0] sbWrMask;
  wire  sbWrEn;
  wire  sbRdEn;
  wire  stallFromDb;
  wire  stallFromSb;
  wire  T_720;
  wire  T_721;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_723;
  wire  T_724;
  wire  T_726;
  wire  T_727;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_735;
  wire  GEN_15;
  wire  GEN_16;
  wire  T_738;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_741;
  wire  T_742;
  wire  T_745;
  wire  GEN_19;
  wire  GEN_20;
  wire  T_750;
  wire  T_751;
  wire  T_754;
  wire  GEN_21;
  wire  GEN_22;
  wire [3:0] T_782;
  wire [2:0] T_783;
  wire [31:0] T_799_0;
  wire [31:0] T_799_1;
  wire [31:0] dbRamWrMask_0;
  wire [31:0] dbRamWrMask_1;
  wire  T_804;
  wire [31:0] T_805;
  wire [31:0] T_806;
  wire [31:0] T_812_0;
  wire [31:0] T_812_1;
  wire [31:0] T_821_0;
  wire [31:0] T_821_1;
  wire [31:0] GEN_0;
  wire [31:0] GEN_23;
  wire [31:0] GEN_24;
  wire [31:0] GEN_1;
  wire [31:0] GEN_25;
  wire [63:0] T_828;
  wire [63:0] T_829;
  wire  T_830;
  wire  T_831;
  wire  T_832;
  wire  T_834;
  wire  T_835;
  wire  T_837;
  wire [63:0] dbRamWrDataVec;
  wire [63:0] T_838;
  wire [63:0] T_839;
  wire [63:0] T_840;
  wire [63:0] T_841;
  wire [63:0] T_842;
  wire [63:0] T_845;
  wire [63:0] T_846;
  wire  T_847;
  wire [2:0] T_848;
  wire [2:0] T_849;
  wire  T_852;
  wire  T_875_interrupt;
  wire  T_875_haltnot;
  wire [9:0] T_875_reserved0;
  wire [2:0] T_875_buserror;
  wire [2:0] T_875_serial;
  wire  T_875_autoincrement;
  wire [2:0] T_875_access;
  wire [9:0] T_875_hartid;
  wire  T_875_ndreset;
  wire  T_875_fullreset;
  wire  T_886;
  wire  T_887;
  wire [9:0] T_888;
  wire [2:0] T_889;
  wire  T_890;
  wire [2:0] T_891;
  wire [2:0] T_892;
  wire [9:0] T_893;
  wire  T_894;
  wire  T_895;
  wire  T_904_interrupt;
  wire  T_904_haltnot;
  wire [31:0] T_904_data;
  wire [31:0] T_908;
  wire  T_913;
  wire  T_915;
  wire  GEN_31;
  wire  T_917;
  wire  T_919;
  wire  T_920;
  wire  GEN_32;
  wire  T_924;
  wire  T_925;
  wire  GEN_33;
  wire  GEN_34;
  wire [9:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire [2:0] GEN_39;
  wire [9:0] GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  GEN_44;
  wire  T_933;
  wire  T_935;
  wire [1:0] T_938;
  wire  T_939;
  wire  T_940;
  wire  GEN_45;
  wire [9:0] GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_945;
  wire  GEN_49;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_958;
  wire [31:0] GEN_50;
  wire [1:0] T_963;
  wire [33:0] T_964;
  wire [33:0] GEN_51;
  wire [1:0] T_970;
  wire [3:0] T_971;
  wire [13:0] T_972;
  wire [15:0] T_973;
  wire [5:0] T_974;
  wire [1:0] T_975;
  wire [11:0] T_976;
  wire [17:0] T_977;
  wire [33:0] T_978;
  wire [33:0] GEN_53;
  wire  T_980;
  wire  T_986;
  wire [2:0] T_987;
  wire [4:0] T_988;
  wire [3:0] T_989;
  wire [6:0] T_990;
  wire [10:0] T_991;
  wire [15:0] T_992;
  wire [1:0] T_993;
  wire [1:0] T_994;
  wire [3:0] T_995;
  wire [4:0] T_996;
  wire [8:0] T_997;
  wire [13:0] T_998;
  wire [17:0] T_999;
  wire [33:0] T_1000;
  wire [33:0] GEN_54;
  wire  T_1002;
  wire  T_1009;
  wire  T_1010;
  wire  T_1011;
  wire [33:0] GEN_55;
  wire [2:0] T_1013;
  wire  T_1015;
  wire  T_1025;
  wire  T_1026;
  wire  T_1027;
  wire [33:0] GEN_56;
  wire  T_1040;
  wire  T_1041;
  wire [33:0] GEN_57;
  wire  T_1043;
  wire  T_1045;
  wire  T_1046;
  wire  T_1048;
  wire  T_1051;
  wire  T_1052;
  wire  T_1053;
  wire [1:0] T_1056;
  wire  T_1058;
  wire  T_1059;
  wire  T_1061;
  wire  T_1062;
  wire  T_1063;
  wire  T_1064;
  wire  T_1066;
  wire  T_1068;
  wire  GEN_58;
  wire [33:0] GEN_59;
  wire [1:0] GEN_60;
  wire  GEN_61;
  wire [33:0] GEN_62;
  wire [1:0] GEN_63;
  wire  T_1073;
  wire  T_1074;
  wire  GEN_64;
  wire [33:0] GEN_65;
  wire [1:0] GEN_66;
  wire  T_1078;
  wire  T_1079;
  wire  GEN_67;
  wire  GEN_68;
  wire [33:0] GEN_69;
  wire [1:0] GEN_70;
  wire [63:0] T_1101_0;
  wire [63:0] T_1101_1;
  wire [63:0] T_1101_2;
  wire [63:0] T_1101_3;
  wire [63:0] T_1101_4;
  wire [63:0] T_1101_5;
  wire [63:0] T_1101_6;
  wire [63:0] T_1101_7;
  wire [63:0] T_1101_8;
  wire [63:0] T_1101_9;
  wire [63:0] T_1101_10;
  wire [63:0] T_1101_11;
  wire [63:0] T_1101_12;
  wire [63:0] T_1101_13;
  wire [63:0] T_1101_14;
  wire [3:0] T_1104;
  wire [3:0] T_1105;
  wire [63:0] GEN_6;
  wire [63:0] GEN_71;
  wire [63:0] GEN_72;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire [63:0] GEN_75;
  wire [63:0] GEN_76;
  wire [63:0] GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] GEN_79;
  wire [63:0] GEN_80;
  wire [63:0] GEN_81;
  wire [63:0] GEN_82;
  wire [63:0] GEN_83;
  wire [63:0] GEN_84;
  wire [31:0] T_1109;
  wire [31:0] T_1110;
  wire [31:0] T_1116_0;
  wire [31:0] T_1116_1;
  wire [31:0] T_1118;
  wire [31:0] T_1119;
  wire [31:0] T_1125_0;
  wire [31:0] T_1125_1;
  wire [31:0] GEN_7;
  wire [31:0] GEN_8;
  wire [3:0] T_1131;
  wire  T_1133;
  wire  GEN_87;
  wire [8:0] T_1134;
  wire  T_1137;
  wire [31:0] GEN_9;
  wire  T_1141;
  wire  T_1142;
  wire  T_1143;
  wire  T_1147;
  wire [31:0] GEN_10;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire [63:0] GEN_91;
  wire  GEN_92;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1167;
  wire  T_1168;
  wire [63:0] GEN_93;
  wire  T_1172;
  wire  T_1173;
  wire [63:0] GEN_94;
  reg [25:0] sbAcqReg_addr_block;
  reg [31:0] GEN_115;
  reg [1:0] sbAcqReg_client_xact_id;
  reg [31:0] GEN_116;
  reg [2:0] sbAcqReg_addr_beat;
  reg [31:0] GEN_117;
  reg  sbAcqReg_is_builtin_type;
  reg [31:0] GEN_118;
  reg [2:0] sbAcqReg_a_type;
  reg [31:0] GEN_119;
  reg [10:0] sbAcqReg_union;
  reg [31:0] GEN_120;
  reg [63:0] sbAcqReg_data;
  reg [63:0] GEN_121;
  reg  sbAcqValidReg;
  reg [31:0] GEN_122;
  wire  T_1202;
  wire  sbReg_get;
  wire  T_1203;
  wire  sbReg_getblk;
  wire  T_1204;
  wire  sbReg_put;
  wire  T_1205;
  wire  sbReg_putblk;
  wire  sbMultibeat;
  wire [3:0] T_1207;
  wire [2:0] sbBeatInc1;
  wire  sbLast;
  wire [2:0] T_1216_0;
  wire [2:0] T_1216_1;
  wire  T_1218;
  wire  T_1219;
  wire  T_1220;
  wire  T_1221;
  wire [2:0] T_1222;
  wire [2:0] T_1224;
  wire [28:0] T_1225;
  wire [31:0] T_1226;
  wire  T_1227;
  wire  T_1228;
  wire  T_1229;
  wire  T_1230;
  wire  T_1232;
  wire  T_1233;
  wire  T_1257;
  wire [7:0] T_1258;
  wire [7:0] T_1260;
  wire [7:0] T_1261;
  wire  T_1262;
  wire  T_1263;
  wire  T_1264;
  wire  T_1265;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire  T_1269;
  wire [7:0] T_1273;
  wire [7:0] T_1277;
  wire [7:0] T_1281;
  wire [7:0] T_1285;
  wire [7:0] T_1289;
  wire [7:0] T_1293;
  wire [7:0] T_1297;
  wire [7:0] T_1301;
  wire [15:0] T_1302;
  wire [15:0] T_1303;
  wire [31:0] T_1304;
  wire [15:0] T_1305;
  wire [15:0] T_1306;
  wire [31:0] T_1307;
  wire [63:0] T_1308;
  wire  T_1309;
  wire [25:0] GEN_95;
  wire [1:0] GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire [2:0] GEN_99;
  wire [10:0] GEN_100;
  wire [63:0] GEN_101;
  wire  GEN_102;
  wire  T_1311;
  wire  T_1313;
  wire  T_1314;
  wire  GEN_103;
  wire [2:0] GEN_104;
  wire  GEN_105;
  wire  T_1317;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_1335;
  wire [2:0] T_1336;
  wire  T_1337;
  wire [2:0] T_1338;
  wire  T_1339;
  wire [2:0] T_1340;
  wire  T_1341;
  wire [2:0] T_1342;
  wire  T_1343;
  wire [2:0] T_1344;
  wire  T_1345;
  wire [2:0] T_1346;
  wire  T_1347;
  wire [2:0] T_1348;
  wire [2:0] T_1372_addr_beat;
  wire [1:0] T_1372_client_xact_id;
  wire  T_1372_manager_xact_id;
  wire  T_1372_is_builtin_type;
  wire [3:0] T_1372_g_type;
  wire [63:0] T_1372_data;
  wire  T_1397;
  wire  T_1398;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire  sbStall;
  wire  T_1404;
  assign io_db_req_ready = T_1064;
  assign io_db_resp_valid = dbStateReg;
  assign io_db_resp_bits_data = dbRespReg_data;
  assign io_db_resp_bits_resp = dbRespReg_resp;
  assign io_debugInterrupts_0 = interruptRegs_0;
  assign io_tl_acquire_ready = T_1404;
  assign io_tl_grant_valid = sbAcqValidReg;
  assign io_tl_grant_bits_addr_beat = T_1372_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1372_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1372_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1372_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1372_g_type;
  assign io_tl_grant_bits_data = T_1372_data;
  assign io_ndreset = ndresetCtrReg;
  assign io_fullreset = CONTROLReg_fullreset;
  assign CONTROLReset_interrupt = 1'h0;
  assign CONTROLReset_haltnot = 1'h0;
  assign CONTROLReset_reserved0 = 10'h0;
  assign CONTROLReset_buserror = 3'h0;
  assign CONTROLReset_serial = 3'h0;
  assign CONTROLReset_autoincrement = 1'h0;
  assign CONTROLReset_access = 3'h2;
  assign CONTROLReset_hartid = 10'h0;
  assign CONTROLReset_ndreset = 1'h0;
  assign CONTROLReset_fullreset = 1'h0;
  assign CONTROLWrEn = GEN_32;
  assign CONTROLWrData_interrupt = T_875_interrupt;
  assign CONTROLWrData_haltnot = T_875_haltnot;
  assign CONTROLWrData_reserved0 = T_875_reserved0;
  assign CONTROLWrData_buserror = T_875_buserror;
  assign CONTROLWrData_serial = T_875_serial;
  assign CONTROLWrData_autoincrement = T_875_autoincrement;
  assign CONTROLWrData_access = T_875_access;
  assign CONTROLWrData_hartid = T_875_hartid;
  assign CONTROLWrData_ndreset = T_875_ndreset;
  assign CONTROLWrData_fullreset = T_875_fullreset;
  assign CONTROLRdData_interrupt = GEN_2;
  assign CONTROLRdData_haltnot = GEN_3;
  assign CONTROLRdData_reserved0 = CONTROLReg_reserved0;
  assign CONTROLRdData_buserror = CONTROLReg_buserror;
  assign CONTROLRdData_serial = CONTROLReg_serial;
  assign CONTROLRdData_autoincrement = CONTROLReg_autoincrement;
  assign CONTROLRdData_access = CONTROLReg_access;
  assign CONTROLRdData_hartid = CONTROLReg_hartid;
  assign CONTROLRdData_ndreset = ndresetCtrReg;
  assign CONTROLRdData_fullreset = CONTROLReg_fullreset;
  assign DMINFORdData_reserved0 = 2'h0;
  assign DMINFORdData_abussize = 7'h0;
  assign DMINFORdData_serialcount = 4'h0;
  assign DMINFORdData_access128 = 1'h0;
  assign DMINFORdData_access64 = 1'h0;
  assign DMINFORdData_access32 = 1'h0;
  assign DMINFORdData_access16 = 1'h0;
  assign DMINFORdData_accesss8 = 1'h0;
  assign DMINFORdData_dramsize = 6'hf;
  assign DMINFORdData_haltsum = 1'h0;
  assign DMINFORdData_reserved1 = 3'h0;
  assign DMINFORdData_authenticated = 1'h1;
  assign DMINFORdData_authbusy = 1'h0;
  assign DMINFORdData_authtype = 2'h0;
  assign DMINFORdData_version = 2'h1;
  assign HALTSUMRdData_serialfull = 1'h0;
  assign HALTSUMRdData_serialvalid = 1'h0;
  assign HALTSUMRdData_acks = {{31'd0}, haltnotSummary};
  assign RAMWrData_interrupt = T_904_interrupt;
  assign RAMWrData_haltnot = T_904_haltnot;
  assign RAMWrData_data = T_904_data;
  assign RAMRdData_interrupt = GEN_4;
  assign RAMRdData_haltnot = GEN_5;
  assign RAMRdData_data = dbRamRdData;
  assign SETHALTNOTWrEn = T_1143;
  assign SETHALTNOTWrData = GEN_7[9:0];
  assign CLEARDEBINTWrEn = T_1153;
  assign CLEARDEBINTWrData = GEN_8[9:0];
  assign T_655_0 = 1'h0;
  assign T_666_0 = 1'h0;
  assign haltnotStatus_0 = {{31'd0}, haltnotRegs_0};
  assign rdHaltnotStatus = GEN_50;
  assign haltnotSummary = haltnotStatus_0 != 32'h0;
  assign ramMem_T_850_addr = ramAddr;
  assign ramMem_T_850_en = 1'h1;
  assign ramMem_T_850_data = ramMem[ramMem_T_850_addr];
  assign ramMem_T_851_data = ramWrData;
  assign ramMem_T_851_addr = ramAddr;
  assign ramMem_T_851_mask = ramWrEn;
  assign ramMem_T_851_en = ramWrEn;
  assign ramAddr = T_849;
  assign ramRdData = ramMem_T_850_data;
  assign ramWrData = T_846;
  assign ramWrMask = T_829;
  assign ramWrEn = T_852;
  assign dbRamAddr = T_782;
  assign dbRamRdData = GEN_1;
  assign dbRamWrData = dbReq_data[31:0];
  assign dbRamWrEn = GEN_31;
  assign dbRamRdEn = 1'h0;
  assign sbRamAddr = T_783;
  assign sbRamRdData = ramRdData;
  assign sbRamWrData = sbWrData;
  assign sbRamWrEn = GEN_87;
  assign sbRamRdEn = GEN_92;
  assign sbRomRdData = GEN_6;
  assign dbRdEn = T_1066;
  assign dbWrEn = T_1068;
  assign dbRdData = GEN_57;
  assign dbResult_data = dbRdData;
  assign dbResult_resp = T_1056;
  assign dbReq_addr = io_db_req_bits_addr;
  assign dbReq_data = io_db_req_bits_data;
  assign dbReq_op = io_db_req_bits_op;
  assign rdCondWrFailure = T_1046;
  assign dbWrNeeded = T_1053;
  assign sbAddr = T_1226[11:0];
  assign sbRdData = GEN_94;
  assign sbWrData = sbAcqReg_data;
  assign sbWrMask = T_1308;
  assign sbWrEn = T_1230;
  assign sbRdEn = T_1228;
  assign stallFromDb = 1'h0;
  assign stallFromSb = T_831;
  assign T_720 = CONTROLWrData_hartid == 10'h0;
  assign T_721 = interruptRegs_0 | CONTROLWrData_interrupt;
  assign GEN_11 = T_720 ? T_721 : interruptRegs_0;
  assign GEN_12 = CONTROLWrEn ? GEN_11 : interruptRegs_0;
  assign T_723 = CONTROLWrEn == 1'h0;
  assign T_724 = T_723 & dbRamWrEn;
  assign T_726 = CONTROLReg_hartid == 10'h0;
  assign T_727 = interruptRegs_0 | RAMWrData_interrupt;
  assign GEN_13 = T_726 ? T_727 : GEN_12;
  assign GEN_14 = T_724 ? GEN_13 : GEN_12;
  assign T_731 = dbRamWrEn == 1'h0;
  assign T_732 = T_723 & T_731;
  assign T_733 = T_732 & CLEARDEBINTWrEn;
  assign T_735 = CLEARDEBINTWrData == 10'h0;
  assign GEN_15 = T_735 ? 1'h0 : GEN_14;
  assign GEN_16 = T_733 ? GEN_15 : GEN_14;
  assign T_738 = SETHALTNOTWrData == 10'h0;
  assign GEN_17 = T_738 ? 1'h1 : haltnotRegs_0;
  assign GEN_18 = SETHALTNOTWrEn ? GEN_17 : haltnotRegs_0;
  assign T_741 = SETHALTNOTWrEn == 1'h0;
  assign T_742 = T_741 & CONTROLWrEn;
  assign T_745 = haltnotRegs_0 & CONTROLWrData_haltnot;
  assign GEN_19 = T_720 ? T_745 : GEN_18;
  assign GEN_20 = T_742 ? GEN_19 : GEN_18;
  assign T_750 = T_741 & T_723;
  assign T_751 = T_750 & dbRamWrEn;
  assign T_754 = haltnotRegs_0 & RAMWrData_haltnot;
  assign GEN_21 = T_726 ? T_754 : GEN_20;
  assign GEN_22 = T_751 ? GEN_21 : GEN_20;
  assign T_782 = dbReq_addr[3:0];
  assign T_783 = sbAddr[5:3];
  assign T_799_0 = 32'hffffffff;
  assign T_799_1 = 32'hffffffff;
  assign dbRamWrMask_0 = GEN_23;
  assign dbRamWrMask_1 = GEN_24;
  assign T_804 = dbRamAddr[0];
  assign T_805 = ramRdData[31:0];
  assign T_806 = ramRdData[63:32];
  assign T_812_0 = T_805;
  assign T_812_1 = T_806;
  assign T_821_0 = 32'h0;
  assign T_821_1 = 32'h0;
  assign GEN_0 = 32'hffffffff;
  assign GEN_23 = 1'h0 == T_804 ? GEN_0 : T_821_0;
  assign GEN_24 = T_804 ? GEN_0 : T_821_1;
  assign GEN_1 = GEN_25;
  assign GEN_25 = T_804 ? T_812_1 : T_812_0;
  assign T_828 = {dbRamWrMask_1,dbRamWrMask_0};
  assign T_829 = sbRamWrEn ? sbWrMask : T_828;
  assign T_830 = dbRamWrEn | dbRamRdEn;
  assign T_831 = sbRamRdEn | sbRamWrEn;
  assign T_832 = T_830 & T_831;
  assign T_834 = T_832 == 1'h0;
  assign T_835 = T_834 | reset;
  assign T_837 = T_835 == 1'h0;
  assign dbRamWrDataVec = {dbRamWrData,dbRamWrData};
  assign T_838 = ramWrMask & sbRamWrData;
  assign T_839 = ~ ramWrMask;
  assign T_840 = T_839 & ramRdData;
  assign T_841 = T_838 | T_840;
  assign T_842 = ramWrMask & dbRamWrDataVec;
  assign T_845 = T_842 | T_840;
  assign T_846 = sbRamWrEn ? T_841 : T_845;
  assign T_847 = sbRamWrEn | sbRamRdEn;
  assign T_848 = dbRamAddr[3:1];
  assign T_849 = T_847 ? sbRamAddr : T_848;
  assign T_852 = sbRamWrEn | dbRamWrEn;
  assign T_875_interrupt = T_895;
  assign T_875_haltnot = T_894;
  assign T_875_reserved0 = T_893;
  assign T_875_buserror = T_892;
  assign T_875_serial = T_891;
  assign T_875_autoincrement = T_890;
  assign T_875_access = T_889;
  assign T_875_hartid = T_888;
  assign T_875_ndreset = T_887;
  assign T_875_fullreset = T_886;
  assign T_886 = dbReq_data[0];
  assign T_887 = dbReq_data[1];
  assign T_888 = dbReq_data[11:2];
  assign T_889 = dbReq_data[14:12];
  assign T_890 = dbReq_data[15];
  assign T_891 = dbReq_data[18:16];
  assign T_892 = dbReq_data[21:19];
  assign T_893 = dbReq_data[31:22];
  assign T_894 = dbReq_data[32];
  assign T_895 = dbReq_data[33];
  assign T_904_interrupt = T_895;
  assign T_904_haltnot = T_894;
  assign T_904_data = T_908;
  assign T_908 = dbReq_data[31:0];
  assign T_913 = dbReq_addr[4:4];
  assign T_915 = T_913 == 1'h0;
  assign GEN_31 = T_915 ? dbWrEn : 1'h0;
  assign T_917 = dbReq_addr == 5'h10;
  assign T_919 = T_915 == 1'h0;
  assign T_920 = T_919 & T_917;
  assign GEN_32 = T_920 ? dbWrEn : 1'h0;
  assign T_924 = T_917 == 1'h0;
  assign T_925 = T_919 & T_924;
  assign GEN_33 = reset ? CONTROLReset_interrupt : CONTROLReg_interrupt;
  assign GEN_34 = reset ? CONTROLReset_haltnot : CONTROLReg_haltnot;
  assign GEN_35 = reset ? CONTROLReset_reserved0 : CONTROLReg_reserved0;
  assign GEN_36 = reset ? CONTROLReset_buserror : CONTROLReg_buserror;
  assign GEN_37 = reset ? CONTROLReset_serial : CONTROLReg_serial;
  assign GEN_38 = reset ? CONTROLReset_autoincrement : CONTROLReg_autoincrement;
  assign GEN_39 = reset ? CONTROLReset_access : CONTROLReg_access;
  assign GEN_40 = reset ? CONTROLReset_hartid : CONTROLReg_hartid;
  assign GEN_41 = reset ? CONTROLReset_ndreset : CONTROLReg_ndreset;
  assign GEN_42 = reset ? CONTROLReset_fullreset : CONTROLReg_fullreset;
  assign GEN_43 = reset ? 1'h0 : ndresetCtrReg;
  assign T_928 = reset == 1'h0;
  assign T_929 = T_928 & CONTROLWrEn;
  assign T_930 = CONTROLReg_fullreset | CONTROLWrData_fullreset;
  assign GEN_44 = CONTROLWrData_ndreset ? 1'h1 : GEN_43;
  assign T_933 = CONTROLWrData_ndreset == 1'h0;
  assign T_935 = ndresetCtrReg == 1'h0;
  assign T_938 = ndresetCtrReg - 1'h1;
  assign T_939 = T_938[0:0];
  assign T_940 = T_935 ? 1'h0 : T_939;
  assign GEN_45 = T_933 ? T_940 : GEN_44;
  assign GEN_46 = T_929 ? CONTROLWrData_hartid : GEN_40;
  assign GEN_47 = T_929 ? T_930 : GEN_42;
  assign GEN_48 = T_929 ? GEN_45 : GEN_43;
  assign T_945 = T_928 & T_723;
  assign GEN_49 = T_945 ? T_940 : GEN_48;
  assign GEN_2 = interruptRegs_0;
  assign GEN_3 = haltnotRegs_0;
  assign GEN_4 = interruptRegs_0;
  assign GEN_5 = haltnotRegs_0;
  assign T_958 = dbReq_addr == 5'h0;
  assign GEN_50 = T_958 ? haltnotStatus_0 : 32'h0;
  assign T_963 = {RAMRdData_interrupt,RAMRdData_haltnot};
  assign T_964 = {T_963,RAMRdData_data};
  assign GEN_51 = T_915 ? T_964 : 34'h0;
  assign T_970 = {CONTROLRdData_ndreset,CONTROLRdData_fullreset};
  assign T_971 = {CONTROLRdData_autoincrement,CONTROLRdData_access};
  assign T_972 = {T_971,CONTROLRdData_hartid};
  assign T_973 = {T_972,T_970};
  assign T_974 = {CONTROLRdData_buserror,CONTROLRdData_serial};
  assign T_975 = {CONTROLRdData_interrupt,CONTROLRdData_haltnot};
  assign T_976 = {T_975,CONTROLRdData_reserved0};
  assign T_977 = {T_976,T_974};
  assign T_978 = {T_977,T_973};
  assign GEN_53 = T_920 ? T_978 : GEN_51;
  assign T_980 = dbReq_addr == 5'h11;
  assign T_986 = T_925 & T_980;
  assign T_987 = {DMINFORdData_authbusy,DMINFORdData_authtype};
  assign T_988 = {T_987,DMINFORdData_version};
  assign T_989 = {DMINFORdData_reserved1,DMINFORdData_authenticated};
  assign T_990 = {DMINFORdData_dramsize,DMINFORdData_haltsum};
  assign T_991 = {T_990,T_989};
  assign T_992 = {T_991,T_988};
  assign T_993 = {DMINFORdData_access16,DMINFORdData_accesss8};
  assign T_994 = {DMINFORdData_access64,DMINFORdData_access32};
  assign T_995 = {T_994,T_993};
  assign T_996 = {DMINFORdData_serialcount,DMINFORdData_access128};
  assign T_997 = {DMINFORdData_reserved0,DMINFORdData_abussize};
  assign T_998 = {T_997,T_996};
  assign T_999 = {T_998,T_995};
  assign T_1000 = {T_999,T_992};
  assign GEN_54 = T_986 ? T_1000 : GEN_53;
  assign T_1002 = dbReq_addr == 5'h1b;
  assign T_1009 = T_980 == 1'h0;
  assign T_1010 = T_925 & T_1009;
  assign T_1011 = T_1010 & T_1002;
  assign GEN_55 = T_1011 ? 34'h0 : GEN_54;
  assign T_1013 = dbReq_addr[4:2];
  assign T_1015 = T_1013 == 3'h7;
  assign T_1025 = T_1002 == 1'h0;
  assign T_1026 = T_1010 & T_1025;
  assign T_1027 = T_1026 & T_1015;
  assign GEN_56 = T_1027 ? {{2'd0}, rdHaltnotStatus} : GEN_55;
  assign T_1040 = T_1015 == 1'h0;
  assign T_1041 = T_1026 & T_1040;
  assign GEN_57 = T_1041 ? 34'h0 : GEN_56;
  assign T_1043 = dbRdData[33];
  assign T_1045 = dbReq_op == 2'h3;
  assign T_1046 = T_1043 & T_1045;
  assign T_1048 = dbReq_op == 2'h2;
  assign T_1051 = ~ rdCondWrFailure;
  assign T_1052 = T_1045 & T_1051;
  assign T_1053 = T_1048 | T_1052;
  assign T_1056 = rdCondWrFailure ? 2'h1 : 2'h0;
  assign T_1058 = stallFromSb == 1'h0;
  assign T_1059 = dbStateReg == 1'h0;
  assign T_1061 = io_db_resp_ready & io_db_resp_valid;
  assign T_1062 = dbStateReg & T_1061;
  assign T_1063 = T_1059 | T_1062;
  assign T_1064 = T_1058 & T_1063;
  assign T_1066 = io_db_req_ready & io_db_req_valid;
  assign T_1068 = dbWrNeeded & T_1066;
  assign GEN_58 = T_1066 ? 1'h1 : dbStateReg;
  assign GEN_59 = T_1066 ? dbResult_data : dbRespReg_data;
  assign GEN_60 = T_1066 ? dbResult_resp : dbRespReg_resp;
  assign GEN_61 = T_1059 ? GEN_58 : dbStateReg;
  assign GEN_62 = T_1059 ? GEN_59 : dbRespReg_data;
  assign GEN_63 = T_1059 ? GEN_60 : dbRespReg_resp;
  assign T_1073 = T_1059 == 1'h0;
  assign T_1074 = T_1073 & dbStateReg;
  assign GEN_64 = T_1066 ? 1'h1 : GEN_61;
  assign GEN_65 = T_1066 ? dbResult_data : GEN_62;
  assign GEN_66 = T_1066 ? dbResult_resp : GEN_63;
  assign T_1078 = T_1066 == 1'h0;
  assign T_1079 = T_1078 & T_1061;
  assign GEN_67 = T_1079 ? 1'h0 : GEN_64;
  assign GEN_68 = T_1074 ? GEN_67 : GEN_61;
  assign GEN_69 = T_1074 ? GEN_65 : GEN_62;
  assign GEN_70 = T_1074 ? GEN_66 : GEN_63;
  assign T_1101_0 = 64'hc0006f03c0006f;
  assign T_1101_1 = 64'h80006ffff00413;
  assign T_1101_2 = 64'hff0000f00000413;
  assign T_1101_3 = 64'h42802e2343803483;
  assign T_1101_4 = 64'h10802023f1402473;
  assign T_1101_5 = 64'h8474137b002473;
  assign T_1101_6 = 64'h7b20247302041a63;
  assign T_1101_7 = 64'h7b2410737b200073;
  assign T_1101_8 = 64'h1c0474137b002473;
  assign T_1101_9 = 64'h41663f4040413;
  assign T_1101_10 = 64'h4000006742903c23;
  assign T_1101_11 = 64'h10802623f1402473;
  assign T_1101_12 = 64'h7b0024737b046073;
  assign T_1101_13 = 64'hfe040ce302047413;
  assign T_1101_14 = 64'hfe1ff06f;
  assign T_1104 = T_1105;
  assign T_1105 = sbAddr[6:3];
  assign GEN_6 = GEN_84;
  assign GEN_71 = 4'h1 == T_1104 ? T_1101_1 : T_1101_0;
  assign GEN_72 = 4'h2 == T_1104 ? T_1101_2 : GEN_71;
  assign GEN_73 = 4'h3 == T_1104 ? T_1101_3 : GEN_72;
  assign GEN_74 = 4'h4 == T_1104 ? T_1101_4 : GEN_73;
  assign GEN_75 = 4'h5 == T_1104 ? T_1101_5 : GEN_74;
  assign GEN_76 = 4'h6 == T_1104 ? T_1101_6 : GEN_75;
  assign GEN_77 = 4'h7 == T_1104 ? T_1101_7 : GEN_76;
  assign GEN_78 = 4'h8 == T_1104 ? T_1101_8 : GEN_77;
  assign GEN_79 = 4'h9 == T_1104 ? T_1101_9 : GEN_78;
  assign GEN_80 = 4'ha == T_1104 ? T_1101_10 : GEN_79;
  assign GEN_81 = 4'hb == T_1104 ? T_1101_11 : GEN_80;
  assign GEN_82 = 4'hc == T_1104 ? T_1101_12 : GEN_81;
  assign GEN_83 = 4'hd == T_1104 ? T_1101_13 : GEN_82;
  assign GEN_84 = 4'he == T_1104 ? T_1101_14 : GEN_83;
  assign T_1109 = sbWrData[31:0];
  assign T_1110 = sbWrData[63:32];
  assign T_1116_0 = T_1109;
  assign T_1116_1 = T_1110;
  assign T_1118 = sbWrMask[31:0];
  assign T_1119 = sbWrMask[63:32];
  assign T_1125_0 = T_1118;
  assign T_1125_1 = T_1119;
  assign GEN_7 = T_1116_1;
  assign GEN_8 = T_1116_0;
  assign T_1131 = sbAddr[11:8];
  assign T_1133 = T_1131 == 4'h4;
  assign GEN_87 = T_1133 ? sbWrEn : 1'h0;
  assign T_1134 = sbAddr[11:3];
  assign T_1137 = T_1134 == 9'h21;
  assign GEN_9 = T_1125_1;
  assign T_1141 = GEN_9 != 32'h0;
  assign T_1142 = T_1137 & T_1141;
  assign T_1143 = T_1142 & sbWrEn;
  assign T_1147 = T_1134 == 9'h20;
  assign GEN_10 = T_1125_0;
  assign T_1151 = GEN_10 != 32'h0;
  assign T_1152 = T_1147 & T_1151;
  assign T_1153 = T_1152 & sbWrEn;
  assign GEN_91 = T_1133 ? sbRamRdData : 64'h0;
  assign GEN_92 = T_1133 ? sbRdEn : 1'h0;
  assign T_1163 = T_1131 == 4'h8;
  assign T_1164 = T_1131 == 4'h9;
  assign T_1165 = T_1163 | T_1164;
  assign T_1167 = T_1133 == 1'h0;
  assign T_1168 = T_1167 & T_1165;
  assign GEN_93 = T_1168 ? sbRomRdData : GEN_91;
  assign T_1172 = T_1165 == 1'h0;
  assign T_1173 = T_1167 & T_1172;
  assign GEN_94 = T_1173 ? 64'h0 : GEN_93;
  assign T_1202 = sbAcqReg_a_type == 3'h0;
  assign sbReg_get = sbAcqReg_is_builtin_type & T_1202;
  assign T_1203 = sbAcqReg_a_type == 3'h1;
  assign sbReg_getblk = sbAcqReg_is_builtin_type & T_1203;
  assign T_1204 = sbAcqReg_a_type == 3'h2;
  assign sbReg_put = sbAcqReg_is_builtin_type & T_1204;
  assign T_1205 = sbAcqReg_a_type == 3'h3;
  assign sbReg_putblk = sbAcqReg_is_builtin_type & T_1205;
  assign sbMultibeat = sbReg_getblk & sbAcqValidReg;
  assign T_1207 = sbAcqReg_addr_beat + 3'h1;
  assign sbBeatInc1 = T_1207[2:0];
  assign sbLast = sbAcqReg_addr_beat == 3'h7;
  assign T_1216_0 = 3'h0;
  assign T_1216_1 = 3'h4;
  assign T_1218 = sbAcqReg_a_type == T_1216_0;
  assign T_1219 = sbAcqReg_a_type == T_1216_1;
  assign T_1220 = T_1218 | T_1219;
  assign T_1221 = sbAcqReg_is_builtin_type & T_1220;
  assign T_1222 = sbAcqReg_union[10:8];
  assign T_1224 = T_1221 ? T_1222 : 3'h0;
  assign T_1225 = {sbAcqReg_addr_block,sbAcqReg_addr_beat};
  assign T_1226 = {T_1225,T_1224};
  assign T_1227 = sbReg_get | sbReg_getblk;
  assign T_1228 = sbAcqValidReg & T_1227;
  assign T_1229 = sbReg_put | sbReg_putblk;
  assign T_1230 = sbAcqValidReg & T_1229;
  assign T_1232 = sbAcqReg_a_type == 3'h4;
  assign T_1233 = sbAcqReg_is_builtin_type & T_1232;
  assign T_1257 = sbReg_putblk | sbReg_put;
  assign T_1258 = sbAcqReg_union[8:1];
  assign T_1260 = T_1257 ? T_1258 : 8'h0;
  assign T_1261 = T_1233 ? 8'hff : T_1260;
  assign T_1262 = T_1261[0];
  assign T_1263 = T_1261[1];
  assign T_1264 = T_1261[2];
  assign T_1265 = T_1261[3];
  assign T_1266 = T_1261[4];
  assign T_1267 = T_1261[5];
  assign T_1268 = T_1261[6];
  assign T_1269 = T_1261[7];
  assign T_1273 = T_1262 ? 8'hff : 8'h0;
  assign T_1277 = T_1263 ? 8'hff : 8'h0;
  assign T_1281 = T_1264 ? 8'hff : 8'h0;
  assign T_1285 = T_1265 ? 8'hff : 8'h0;
  assign T_1289 = T_1266 ? 8'hff : 8'h0;
  assign T_1293 = T_1267 ? 8'hff : 8'h0;
  assign T_1297 = T_1268 ? 8'hff : 8'h0;
  assign T_1301 = T_1269 ? 8'hff : 8'h0;
  assign T_1302 = {T_1277,T_1273};
  assign T_1303 = {T_1285,T_1281};
  assign T_1304 = {T_1303,T_1302};
  assign T_1305 = {T_1293,T_1289};
  assign T_1306 = {T_1301,T_1297};
  assign T_1307 = {T_1306,T_1305};
  assign T_1308 = {T_1307,T_1304};
  assign T_1309 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign GEN_95 = T_1309 ? io_tl_acquire_bits_addr_block : sbAcqReg_addr_block;
  assign GEN_96 = T_1309 ? io_tl_acquire_bits_client_xact_id : sbAcqReg_client_xact_id;
  assign GEN_97 = T_1309 ? io_tl_acquire_bits_addr_beat : sbAcqReg_addr_beat;
  assign GEN_98 = T_1309 ? io_tl_acquire_bits_is_builtin_type : sbAcqReg_is_builtin_type;
  assign GEN_99 = T_1309 ? io_tl_acquire_bits_a_type : sbAcqReg_a_type;
  assign GEN_100 = T_1309 ? io_tl_acquire_bits_union : sbAcqReg_union;
  assign GEN_101 = T_1309 ? io_tl_acquire_bits_data : sbAcqReg_data;
  assign GEN_102 = T_1309 ? 1'h1 : sbAcqValidReg;
  assign T_1311 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1313 = T_1309 == 1'h0;
  assign T_1314 = T_1313 & T_1311;
  assign GEN_103 = sbLast ? 1'h0 : GEN_102;
  assign GEN_104 = sbMultibeat ? sbBeatInc1 : GEN_97;
  assign GEN_105 = sbMultibeat ? GEN_103 : GEN_102;
  assign T_1317 = sbMultibeat == 1'h0;
  assign GEN_106 = T_1317 ? 1'h0 : GEN_105;
  assign GEN_107 = T_1314 ? GEN_104 : GEN_97;
  assign GEN_108 = T_1314 ? GEN_106 : GEN_102;
  assign T_1335 = 3'h6 == sbAcqReg_a_type;
  assign T_1336 = T_1335 ? 3'h1 : 3'h3;
  assign T_1337 = 3'h5 == sbAcqReg_a_type;
  assign T_1338 = T_1337 ? 3'h1 : T_1336;
  assign T_1339 = 3'h4 == sbAcqReg_a_type;
  assign T_1340 = T_1339 ? 3'h4 : T_1338;
  assign T_1341 = 3'h3 == sbAcqReg_a_type;
  assign T_1342 = T_1341 ? 3'h3 : T_1340;
  assign T_1343 = 3'h2 == sbAcqReg_a_type;
  assign T_1344 = T_1343 ? 3'h3 : T_1342;
  assign T_1345 = 3'h1 == sbAcqReg_a_type;
  assign T_1346 = T_1345 ? 3'h5 : T_1344;
  assign T_1347 = 3'h0 == sbAcqReg_a_type;
  assign T_1348 = T_1347 ? 3'h4 : T_1346;
  assign T_1372_addr_beat = sbAcqReg_addr_beat;
  assign T_1372_client_xact_id = sbAcqReg_client_xact_id;
  assign T_1372_manager_xact_id = 1'h0;
  assign T_1372_is_builtin_type = 1'h1;
  assign T_1372_g_type = {{1'd0}, T_1348};
  assign T_1372_data = sbRdData;
  assign T_1397 = sbLast == 1'h0;
  assign T_1398 = sbMultibeat & T_1397;
  assign T_1400 = io_tl_grant_ready == 1'h0;
  assign T_1401 = io_tl_grant_valid & T_1400;
  assign T_1402 = T_1398 | T_1401;
  assign sbStall = T_1402 | stallFromDb;
  assign T_1404 = sbStall == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_26 = {1{$random}};
  CONTROLReg_interrupt = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_27 = {1{$random}};
  CONTROLReg_haltnot = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  CONTROLReg_reserved0 = GEN_28[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  CONTROLReg_buserror = GEN_29[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  CONTROLReg_serial = GEN_30[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_52 = {1{$random}};
  CONTROLReg_autoincrement = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_85 = {1{$random}};
  CONTROLReg_access = GEN_85[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_86 = {1{$random}};
  CONTROLReg_hartid = GEN_86[9:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_88 = {1{$random}};
  CONTROLReg_ndreset = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_89 = {1{$random}};
  CONTROLReg_fullreset = GEN_89[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_90 = {1{$random}};
  ndresetCtrReg = GEN_90[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_109 = {1{$random}};
  interruptRegs_0 = GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_110 = {1{$random}};
  haltnotRegs_0 = GEN_110[0:0];
  `endif
  GEN_111 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ramMem[initvar] = GEN_111[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_112 = {1{$random}};
  dbStateReg = GEN_112[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_113 = {2{$random}};
  dbRespReg_data = GEN_113[33:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_114 = {1{$random}};
  dbRespReg_resp = GEN_114[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_115 = {1{$random}};
  sbAcqReg_addr_block = GEN_115[25:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_116 = {1{$random}};
  sbAcqReg_client_xact_id = GEN_116[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_117 = {1{$random}};
  sbAcqReg_addr_beat = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_118 = {1{$random}};
  sbAcqReg_is_builtin_type = GEN_118[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_119 = {1{$random}};
  sbAcqReg_a_type = GEN_119[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_120 = {1{$random}};
  sbAcqReg_union = GEN_120[10:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_121 = {2{$random}};
  sbAcqReg_data = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_122 = {1{$random}};
  sbAcqValidReg = GEN_122[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_interrupt <= CONTROLReset_interrupt;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_haltnot <= CONTROLReset_haltnot;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_reserved0 <= CONTROLReset_reserved0;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_buserror <= CONTROLReset_buserror;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_serial <= CONTROLReset_serial;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_autoincrement <= CONTROLReset_autoincrement;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_access <= CONTROLReset_access;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_hartid <= CONTROLWrData_hartid;
      end else begin
        if(reset) begin
          CONTROLReg_hartid <= CONTROLReset_hartid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_ndreset <= CONTROLReset_ndreset;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_fullreset <= T_930;
      end else begin
        if(reset) begin
          CONTROLReg_fullreset <= CONTROLReset_fullreset;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_945) begin
        if(T_935) begin
          ndresetCtrReg <= 1'h0;
        end else begin
          ndresetCtrReg <= T_939;
        end
      end else begin
        if(T_929) begin
          if(T_933) begin
            if(T_935) begin
              ndresetCtrReg <= 1'h0;
            end else begin
              ndresetCtrReg <= T_939;
            end
          end else begin
            if(CONTROLWrData_ndreset) begin
              ndresetCtrReg <= 1'h1;
            end else begin
              if(reset) begin
                ndresetCtrReg <= 1'h0;
              end
            end
          end
        end else begin
          if(reset) begin
            ndresetCtrReg <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      interruptRegs_0 <= T_655_0;
    end else begin
      if(T_733) begin
        if(T_735) begin
          interruptRegs_0 <= 1'h0;
        end else begin
          if(T_724) begin
            if(T_726) begin
              interruptRegs_0 <= T_727;
            end else begin
              if(CONTROLWrEn) begin
                if(T_720) begin
                  interruptRegs_0 <= T_721;
                end
              end
            end
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end
      end else begin
        if(T_724) begin
          if(T_726) begin
            interruptRegs_0 <= T_727;
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end else begin
          if(CONTROLWrEn) begin
            if(T_720) begin
              interruptRegs_0 <= T_721;
            end
          end
        end
      end
    end
    if(reset) begin
      haltnotRegs_0 <= T_666_0;
    end else begin
      if(T_751) begin
        if(T_726) begin
          haltnotRegs_0 <= T_754;
        end else begin
          if(T_742) begin
            if(T_720) begin
              haltnotRegs_0 <= T_745;
            end else begin
              if(SETHALTNOTWrEn) begin
                if(T_738) begin
                  haltnotRegs_0 <= 1'h1;
                end
              end
            end
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_742) begin
          if(T_720) begin
            haltnotRegs_0 <= T_745;
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end else begin
          if(SETHALTNOTWrEn) begin
            if(T_738) begin
              haltnotRegs_0 <= 1'h1;
            end
          end
        end
      end
    end
    if(ramMem_T_851_en & ramMem_T_851_mask) begin
      ramMem[ramMem_T_851_addr] <= ramMem_T_851_data;
    end
    if(reset) begin
      dbStateReg <= 1'h0;
    end else begin
      if(T_1074) begin
        if(T_1079) begin
          dbStateReg <= 1'h0;
        end else begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end else begin
            if(T_1059) begin
              if(T_1066) begin
                dbStateReg <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_data <= dbResult_data;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_data <= dbResult_data;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_data <= dbResult_data;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_resp <= dbResult_resp;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_resp <= dbResult_resp;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_resp <= dbResult_resp;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_addr_block <= io_tl_acquire_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_client_xact_id <= io_tl_acquire_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1314) begin
        if(sbMultibeat) begin
          sbAcqReg_addr_beat <= sbBeatInc1;
        end else begin
          if(T_1309) begin
            sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
          end
        end
      end else begin
        if(T_1309) begin
          sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_is_builtin_type <= io_tl_acquire_bits_is_builtin_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_a_type <= io_tl_acquire_bits_a_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_union <= io_tl_acquire_bits_union;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1309) begin
        sbAcqReg_data <= io_tl_acquire_bits_data;
      end
    end
    if(reset) begin
      sbAcqValidReg <= 1'h0;
    end else begin
      if(T_1314) begin
        if(T_1317) begin
          sbAcqValidReg <= 1'h0;
        end else begin
          if(sbMultibeat) begin
            if(sbLast) begin
              sbAcqValidReg <= 1'h0;
            end else begin
              if(T_1309) begin
                sbAcqValidReg <= 1'h1;
              end
            end
          end else begin
            if(T_1309) begin
              sbAcqValidReg <= 1'h1;
            end
          end
        end
      end else begin
        if(T_1309) begin
          sbAcqValidReg <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_837) begin
          $fwrite(32'h80000002,"Assertion failed: Stall logic should have prevented concurrent SB/DB RAM Access\n    at Debug.scala:650 assert (!((dbRamWrEn | dbRamRdEn) & (sbRamRdEn | sbRamWrEn)), \"Stall logic should have prevented concurrent SB/DB RAM Access\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_837) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module PRCI(
  input   clk,
  input   reset,
  input   io_interrupts_0_meip,
  input   io_interrupts_0_seip,
  input   io_interrupts_0_debug,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_tiles_0_reset,
  output  io_tiles_0_id,
  output  io_tiles_0_interrupts_meip,
  output  io_tiles_0_interrupts_seip,
  output  io_tiles_0_interrupts_debug,
  output  io_tiles_0_interrupts_mtip,
  output  io_tiles_0_interrupts_msip,
  input   io_rtcTick
);
  reg [63:0] timecmp_0;
  reg [63:0] GEN_3;
  reg [63:0] time$;
  reg [63:0] GEN_4;
  wire [64:0] T_525;
  wire [63:0] T_526;
  wire [63:0] GEN_0;
  wire [31:0] T_533_0;
  reg [31:0] ipi_0;
  reg [31:0] GEN_5;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire [2:0] T_568_0;
  wire [2:0] T_568_1;
  wire  T_570;
  wire  T_571;
  wire  T_572;
  wire  T_573;
  wire [2:0] T_574;
  wire [2:0] T_576;
  wire [28:0] T_577;
  wire [31:0] T_578;
  wire [15:0] addr;
  wire [63:0] rdata;
  wire  T_598;
  wire [2:0] T_599;
  wire  T_600;
  wire [2:0] T_601;
  wire  T_602;
  wire [2:0] T_603;
  wire  T_604;
  wire [2:0] T_605;
  wire  T_606;
  wire [2:0] T_607;
  wire  T_608;
  wire [2:0] T_609;
  wire  T_610;
  wire [2:0] T_611;
  wire [2:0] T_636_addr_beat;
  wire [1:0] T_636_client_xact_id;
  wire  T_636_manager_xact_id;
  wire  T_636_is_builtin_type;
  wire [3:0] T_636_g_type;
  wire [63:0] T_636_data;
  wire  T_658;
  wire  T_659;
  wire [2:0] T_667_0;
  wire [2:0] T_667_1;
  wire [2:0] T_685_0;
  wire [2:0] T_685_1;
  wire  T_697;
  wire  T_698;
  wire  T_717;
  wire  T_718;
  wire  T_720;
  wire  T_721;
  wire  T_722;
  wire [7:0] T_723;
  wire [7:0] T_725;
  wire [7:0] T_726;
  wire  T_727;
  wire  T_728;
  wire  T_729;
  wire  T_730;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_734;
  wire [7:0] T_738;
  wire [7:0] T_742;
  wire [7:0] T_746;
  wire [7:0] T_750;
  wire [7:0] T_754;
  wire [7:0] T_758;
  wire [7:0] T_762;
  wire [7:0] T_766;
  wire [15:0] T_767;
  wire [15:0] T_768;
  wire [31:0] T_769;
  wire [15:0] T_770;
  wire [15:0] T_771;
  wire [31:0] T_772;
  wire [63:0] T_773;
  wire [63:0] T_774;
  wire [63:0] T_853;
  wire [63:0] T_854;
  wire [63:0] T_855;
  wire  T_859;
  wire [63:0] GEN_2;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire  T_865;
  wire  T_867;
  wire  T_868;
  wire [2:0] T_877_0;
  wire [2:0] T_877_1;
  wire [2:0] T_895_0;
  wire [2:0] T_895_1;
  wire [63:0] T_1064;
  wire [63:0] T_1065;
  wire [63:0] GEN_10;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire  T_1077;
  wire  T_1078;
  wire [2:0] T_1087_0;
  wire [2:0] T_1087_1;
  wire [2:0] T_1105_0;
  wire [2:0] T_1105_1;
  wire [63:0] GEN_25;
  wire [63:0] T_1274;
  wire [63:0] T_1275;
  wire [63:0] GEN_18;
  wire [63:0] T_1286;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire  T_1287;
  wire  T_1288;
  wire  GEN_1;
  reg [31:0] GEN_6;
  Queue_16 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_636_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_636_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_636_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_636_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_636_g_type;
  assign io_tl_grant_bits_data = T_636_data;
  assign io_tiles_0_reset = GEN_1;
  assign io_tiles_0_id = 1'h0;
  assign io_tiles_0_interrupts_meip = io_interrupts_0_meip;
  assign io_tiles_0_interrupts_seip = io_interrupts_0_seip;
  assign io_tiles_0_interrupts_debug = io_interrupts_0_debug;
  assign io_tiles_0_interrupts_mtip = T_1288;
  assign io_tiles_0_interrupts_msip = T_1287;
  assign T_525 = time$ + 64'h1;
  assign T_526 = T_525[63:0];
  assign GEN_0 = io_rtcTick ? T_526 : time$;
  assign T_533_0 = 32'h0;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_568_0 = 3'h0;
  assign T_568_1 = 3'h4;
  assign T_570 = acq_io_deq_bits_a_type == T_568_0;
  assign T_571 = acq_io_deq_bits_a_type == T_568_1;
  assign T_572 = T_570 | T_571;
  assign T_573 = acq_io_deq_bits_is_builtin_type & T_572;
  assign T_574 = acq_io_deq_bits_union[10:8];
  assign T_576 = T_573 ? T_574 : 3'h0;
  assign T_577 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_578 = {T_577,T_576};
  assign addr = T_578[15:0];
  assign rdata = GEN_24;
  assign T_598 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_599 = T_598 ? 3'h1 : 3'h3;
  assign T_600 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_601 = T_600 ? 3'h1 : T_599;
  assign T_602 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_603 = T_602 ? 3'h4 : T_601;
  assign T_604 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_605 = T_604 ? 3'h3 : T_603;
  assign T_606 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_607 = T_606 ? 3'h3 : T_605;
  assign T_608 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_609 = T_608 ? 3'h5 : T_607;
  assign T_610 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_611 = T_610 ? 3'h4 : T_609;
  assign T_636_addr_beat = 3'h0;
  assign T_636_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_636_manager_xact_id = 1'h0;
  assign T_636_is_builtin_type = 1'h1;
  assign T_636_g_type = {{1'd0}, T_611};
  assign T_636_data = rdata;
  assign T_658 = addr[15];
  assign T_659 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_667_0 = 3'h0;
  assign T_667_1 = 3'h4;
  assign T_685_0 = 3'h0;
  assign T_685_1 = 3'h4;
  assign T_697 = acq_io_deq_bits_a_type == 3'h4;
  assign T_698 = acq_io_deq_bits_is_builtin_type & T_697;
  assign T_717 = acq_io_deq_bits_a_type == 3'h3;
  assign T_718 = acq_io_deq_bits_is_builtin_type & T_717;
  assign T_720 = acq_io_deq_bits_a_type == 3'h2;
  assign T_721 = acq_io_deq_bits_is_builtin_type & T_720;
  assign T_722 = T_718 | T_721;
  assign T_723 = acq_io_deq_bits_union[8:1];
  assign T_725 = T_722 ? T_723 : 8'h0;
  assign T_726 = T_698 ? 8'hff : T_725;
  assign T_727 = T_726[0];
  assign T_728 = T_726[1];
  assign T_729 = T_726[2];
  assign T_730 = T_726[3];
  assign T_731 = T_726[4];
  assign T_732 = T_726[5];
  assign T_733 = T_726[6];
  assign T_734 = T_726[7];
  assign T_738 = T_727 ? 8'hff : 8'h0;
  assign T_742 = T_728 ? 8'hff : 8'h0;
  assign T_746 = T_729 ? 8'hff : 8'h0;
  assign T_750 = T_730 ? 8'hff : 8'h0;
  assign T_754 = T_731 ? 8'hff : 8'h0;
  assign T_758 = T_732 ? 8'hff : 8'h0;
  assign T_762 = T_733 ? 8'hff : 8'h0;
  assign T_766 = T_734 ? 8'hff : 8'h0;
  assign T_767 = {T_742,T_738};
  assign T_768 = {T_750,T_746};
  assign T_769 = {T_768,T_767};
  assign T_770 = {T_758,T_754};
  assign T_771 = {T_766,T_762};
  assign T_772 = {T_771,T_770};
  assign T_773 = {T_772,T_769};
  assign T_774 = acq_io_deq_bits_data & T_773;
  assign T_853 = ~ T_773;
  assign T_854 = time$ & T_853;
  assign T_855 = T_774 | T_854;
  assign T_859 = T_659 & T_721;
  assign GEN_2 = T_859 ? T_855 : GEN_0;
  assign GEN_7 = T_658 ? GEN_2 : GEN_0;
  assign GEN_8 = T_658 ? time$ : 64'h0;
  assign T_865 = addr >= 16'h4000;
  assign T_867 = T_658 == 1'h0;
  assign T_868 = T_867 & T_865;
  assign T_877_0 = 3'h0;
  assign T_877_1 = 3'h4;
  assign T_895_0 = 3'h0;
  assign T_895_1 = 3'h4;
  assign T_1064 = timecmp_0 & T_853;
  assign T_1065 = T_774 | T_1064;
  assign GEN_10 = T_859 ? T_1065 : timecmp_0;
  assign GEN_15 = T_868 ? GEN_10 : timecmp_0;
  assign GEN_16 = T_868 ? timecmp_0 : GEN_8;
  assign T_1077 = T_865 == 1'h0;
  assign T_1078 = T_867 & T_1077;
  assign T_1087_0 = 3'h0;
  assign T_1087_1 = 3'h4;
  assign T_1105_0 = 3'h0;
  assign T_1105_1 = 3'h4;
  assign GEN_25 = {{32'd0}, ipi_0};
  assign T_1274 = GEN_25 & T_853;
  assign T_1275 = T_774 | T_1274;
  assign GEN_18 = T_859 ? T_1275 : {{32'd0}, ipi_0};
  assign T_1286 = GEN_25 & 64'h100000001;
  assign GEN_23 = T_1078 ? GEN_18 : {{32'd0}, ipi_0};
  assign GEN_24 = T_1078 ? T_1286 : GEN_16;
  assign T_1287 = ipi_0[0];
  assign T_1288 = time$ >= timecmp_0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_1 = GEN_6[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {2{$random}};
  timecmp_0 = GEN_3[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_4 = {2{$random}};
  time$ = GEN_4[63:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  ipi_0 = GEN_5[31:0];
  `endif
  GEN_6 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_868) begin
        if(T_859) begin
          timecmp_0 <= T_1065;
        end
      end
    end
    if(reset) begin
      time$ <= 64'h0;
    end else begin
      if(T_658) begin
        if(T_859) begin
          time$ <= T_855;
        end else begin
          if(io_rtcTick) begin
            time$ <= T_526;
          end
        end
      end else begin
        if(io_rtcTick) begin
          time$ <= T_526;
        end
      end
    end
    if(reset) begin
      ipi_0 <= T_533_0;
    end else begin
      ipi_0 <= GEN_23[31:0];
    end
  end
endmodule
module ROMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [10:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [10:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [10:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_446;
  wire  single_beat;
  wire  T_448;
  wire  multi_beat;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_455;
  reg [2:0] addr_beat;
  reg [31:0] GEN_68;
  wire  T_457;
  wire [3:0] T_459;
  wire [2:0] T_460;
  wire [2:0] GEN_1;
  wire  T_461;
  wire [2:0] GEN_2;
  wire [63:0] rom_0;
  wire [63:0] rom_1;
  wire [63:0] rom_2;
  wire [63:0] rom_3;
  wire [63:0] rom_4;
  wire [63:0] rom_5;
  wire [63:0] rom_6;
  wire [63:0] rom_7;
  wire [63:0] rom_8;
  wire [63:0] rom_9;
  wire [63:0] rom_10;
  wire [63:0] rom_11;
  wire [63:0] rom_12;
  wire [63:0] rom_13;
  wire [63:0] rom_14;
  wire [63:0] rom_15;
  wire [63:0] rom_16;
  wire [63:0] rom_17;
  wire [63:0] rom_18;
  wire [63:0] rom_19;
  wire [63:0] rom_20;
  wire [63:0] rom_21;
  wire [63:0] rom_22;
  wire [63:0] rom_23;
  wire [63:0] rom_24;
  wire [63:0] rom_25;
  wire [63:0] rom_26;
  wire [63:0] rom_27;
  wire [63:0] rom_28;
  wire [63:0] rom_29;
  wire [63:0] rom_30;
  wire [63:0] rom_31;
  wire [63:0] rom_32;
  wire [63:0] rom_33;
  wire [63:0] rom_34;
  wire [63:0] rom_35;
  wire [63:0] rom_36;
  wire [63:0] rom_37;
  wire [63:0] rom_38;
  wire [63:0] rom_39;
  wire [63:0] rom_40;
  wire [63:0] rom_41;
  wire [63:0] rom_42;
  wire [63:0] rom_43;
  wire [63:0] rom_44;
  wire [63:0] rom_45;
  wire [63:0] rom_46;
  wire [63:0] rom_47;
  wire [63:0] rom_48;
  wire [63:0] rom_49;
  wire [63:0] rom_50;
  wire [63:0] rom_51;
  wire [63:0] rom_52;
  wire [63:0] rom_53;
  wire [63:0] rom_54;
  wire [63:0] rom_55;
  wire [63:0] rom_56;
  wire [63:0] rom_57;
  wire [63:0] rom_58;
  wire [63:0] rom_59;
  wire [63:0] rom_60;
  wire [63:0] rom_61;
  wire [63:0] rom_62;
  wire [63:0] rom_63;
  wire [63:0] rom_64;
  wire [63:0] rom_65;
  wire [28:0] raddr;
  wire [6:0] T_534;
  wire  T_536;
  wire  T_538;
  wire  last;
  wire  T_539;
  wire  T_556;
  wire [2:0] T_557;
  wire  T_558;
  wire [2:0] T_559;
  wire  T_560;
  wire [2:0] T_561;
  wire  T_562;
  wire [2:0] T_563;
  wire  T_564;
  wire [2:0] T_565;
  wire  T_566;
  wire [2:0] T_567;
  wire  T_568;
  wire [2:0] T_569;
  wire [2:0] T_593_addr_beat;
  wire [1:0] T_593_client_xact_id;
  wire  T_593_manager_xact_id;
  wire  T_593_is_builtin_type;
  wire [3:0] T_593_g_type;
  wire [63:0] T_593_data;
  wire [63:0] GEN_0;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire [63:0] GEN_9;
  wire [63:0] GEN_10;
  wire [63:0] GEN_11;
  wire [63:0] GEN_12;
  wire [63:0] GEN_13;
  wire [63:0] GEN_14;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire [63:0] GEN_17;
  wire [63:0] GEN_18;
  wire [63:0] GEN_19;
  wire [63:0] GEN_20;
  wire [63:0] GEN_21;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_29;
  wire [63:0] GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [63:0] GEN_40;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire [63:0] GEN_55;
  wire [63:0] GEN_56;
  wire [63:0] GEN_57;
  wire [63:0] GEN_58;
  wire [63:0] GEN_59;
  wire [63:0] GEN_60;
  wire [63:0] GEN_61;
  wire [63:0] GEN_62;
  wire [63:0] GEN_63;
  wire [63:0] GEN_64;
  wire [63:0] GEN_65;
  wire [63:0] GEN_66;
  wire [63:0] GEN_67;
  Queue_16 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_acquire_ready = acq_io_enq_ready;
  assign io_grant_valid = acq_io_deq_valid;
  assign io_grant_bits_addr_beat = T_593_addr_beat;
  assign io_grant_bits_client_xact_id = T_593_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_593_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_593_is_builtin_type;
  assign io_grant_bits_g_type = T_593_g_type;
  assign io_grant_bits_data = T_593_data;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_acquire_bits_union;
  assign acq_io_enq_bits_data = io_acquire_bits_data;
  assign acq_io_deq_ready = T_539;
  assign T_446 = acq_io_deq_bits_a_type == 3'h0;
  assign single_beat = acq_io_deq_bits_is_builtin_type & T_446;
  assign T_448 = acq_io_deq_bits_a_type == 3'h1;
  assign multi_beat = acq_io_deq_bits_is_builtin_type & T_448;
  assign T_450 = acq_io_deq_valid == 1'h0;
  assign T_451 = T_450 | single_beat;
  assign T_452 = T_451 | multi_beat;
  assign T_453 = T_452 | reset;
  assign T_455 = T_453 == 1'h0;
  assign T_457 = io_grant_ready & io_grant_valid;
  assign T_459 = addr_beat + 3'h1;
  assign T_460 = T_459[2:0];
  assign GEN_1 = T_457 ? T_460 : addr_beat;
  assign T_461 = io_acquire_ready & io_acquire_valid;
  assign GEN_2 = T_461 ? io_acquire_bits_addr_beat : GEN_1;
  assign rom_0 = 64'h6f;
  assign rom_1 = 64'h102000000000;
  assign rom_2 = 64'h0;
  assign rom_3 = 64'h0;
  assign rom_4 = 64'h200a7b2063696c70;
  assign rom_5 = 64'h7469726f69727020;
  assign rom_6 = 64'h3030303478302079;
  assign rom_7 = 64'h20200a3b30303030;
  assign rom_8 = 64'h20676e69646e6570;
  assign rom_9 = 64'h3031303030347830;
  assign rom_10 = 64'h646e20200a3b3030;
  assign rom_11 = 64'h7d0a3b3220737665;
  assign rom_12 = 64'ha7b206374720a3b;
  assign rom_13 = 64'h3020726464612020;
  assign rom_14 = 64'h6666623030343478;
  assign rom_15 = 64'h61720a3b7d0a3b38;
  assign rom_16 = 64'h203020200a7b206d;
  assign rom_17 = 64'h6461202020200a7b;
  assign rom_18 = 64'h3030387830207264;
  assign rom_19 = 64'h200a3b3030303030;
  assign rom_20 = 64'h20657a6973202020;
  assign rom_21 = 64'h3030303030317830;
  assign rom_22 = 64'h3b7d20200a3b3030;
  assign rom_23 = 64'h65726f630a3b7d0a;
  assign rom_24 = 64'h7b203020200a7b20;
  assign rom_25 = 64'h7b2030202020200a;
  assign rom_26 = 64'h692020202020200a;
  assign rom_27 = 64'h6934367672206173;
  assign rom_28 = 64'h200a3b736466616d;
  assign rom_29 = 64'h6d69742020202020;
  assign rom_30 = 64'h34783020706d6365;
  assign rom_31 = 64'h3b30303034303034;
  assign rom_32 = 64'h692020202020200a;
  assign rom_33 = 64'h3034347830206970;
  assign rom_34 = 64'h200a3b3030303030;
  assign rom_35 = 64'h696c702020202020;
  assign rom_36 = 64'h202020200a7b2063;
  assign rom_37 = 64'ha7b206d20202020;
  assign rom_38 = 64'h2020202020202020;
  assign rom_39 = 64'h3034783020656920;
  assign rom_40 = 64'ha3b303030323030;
  assign rom_41 = 64'h2020202020202020;
  assign rom_42 = 64'h2068736572687420;
  assign rom_43 = 64'h3030303230347830;
  assign rom_44 = 64'h202020200a3b3030;
  assign rom_45 = 64'h616c632020202020;
  assign rom_46 = 64'h3230347830206d69;
  assign rom_47 = 64'h200a3b3430303030;
  assign rom_48 = 64'h7d20202020202020;
  assign rom_49 = 64'h2020202020200a3b;
  assign rom_50 = 64'h20200a7b20732020;
  assign rom_51 = 64'h6920202020202020;
  assign rom_52 = 64'h3030303478302065;
  assign rom_53 = 64'h20200a3b30383032;
  assign rom_54 = 64'h7420202020202020;
  assign rom_55 = 64'h7830206873657268;
  assign rom_56 = 64'h3030303130323034;
  assign rom_57 = 64'h2020202020200a3b;
  assign rom_58 = 64'h6d69616c63202020;
  assign rom_59 = 64'h3130323034783020;
  assign rom_60 = 64'h2020200a3b343030;
  assign rom_61 = 64'ha3b7d2020202020;
  assign rom_62 = 64'h3b7d202020202020;
  assign rom_63 = 64'ha3b7d202020200a;
  assign rom_64 = 64'ha3b7d0a3b7d2020;
  assign rom_65 = 64'h0;
  assign raddr = {acq_io_deq_bits_addr_block,addr_beat};
  assign T_534 = raddr[6:0];
  assign T_536 = multi_beat == 1'h0;
  assign T_538 = addr_beat == 3'h7;
  assign last = T_536 | T_538;
  assign T_539 = io_grant_ready & last;
  assign T_556 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_557 = T_556 ? 3'h1 : 3'h3;
  assign T_558 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_559 = T_558 ? 3'h1 : T_557;
  assign T_560 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_561 = T_560 ? 3'h4 : T_559;
  assign T_562 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_563 = T_562 ? 3'h3 : T_561;
  assign T_564 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_565 = T_564 ? 3'h3 : T_563;
  assign T_566 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_567 = T_566 ? 3'h5 : T_565;
  assign T_568 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_569 = T_568 ? 3'h4 : T_567;
  assign T_593_addr_beat = addr_beat;
  assign T_593_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_593_manager_xact_id = 1'h0;
  assign T_593_is_builtin_type = 1'h1;
  assign T_593_g_type = {{1'd0}, T_569};
  assign T_593_data = GEN_0;
  assign GEN_0 = GEN_67;
  assign GEN_3 = 7'h1 == T_534 ? rom_1 : rom_0;
  assign GEN_4 = 7'h2 == T_534 ? rom_2 : GEN_3;
  assign GEN_5 = 7'h3 == T_534 ? rom_3 : GEN_4;
  assign GEN_6 = 7'h4 == T_534 ? rom_4 : GEN_5;
  assign GEN_7 = 7'h5 == T_534 ? rom_5 : GEN_6;
  assign GEN_8 = 7'h6 == T_534 ? rom_6 : GEN_7;
  assign GEN_9 = 7'h7 == T_534 ? rom_7 : GEN_8;
  assign GEN_10 = 7'h8 == T_534 ? rom_8 : GEN_9;
  assign GEN_11 = 7'h9 == T_534 ? rom_9 : GEN_10;
  assign GEN_12 = 7'ha == T_534 ? rom_10 : GEN_11;
  assign GEN_13 = 7'hb == T_534 ? rom_11 : GEN_12;
  assign GEN_14 = 7'hc == T_534 ? rom_12 : GEN_13;
  assign GEN_15 = 7'hd == T_534 ? rom_13 : GEN_14;
  assign GEN_16 = 7'he == T_534 ? rom_14 : GEN_15;
  assign GEN_17 = 7'hf == T_534 ? rom_15 : GEN_16;
  assign GEN_18 = 7'h10 == T_534 ? rom_16 : GEN_17;
  assign GEN_19 = 7'h11 == T_534 ? rom_17 : GEN_18;
  assign GEN_20 = 7'h12 == T_534 ? rom_18 : GEN_19;
  assign GEN_21 = 7'h13 == T_534 ? rom_19 : GEN_20;
  assign GEN_22 = 7'h14 == T_534 ? rom_20 : GEN_21;
  assign GEN_23 = 7'h15 == T_534 ? rom_21 : GEN_22;
  assign GEN_24 = 7'h16 == T_534 ? rom_22 : GEN_23;
  assign GEN_25 = 7'h17 == T_534 ? rom_23 : GEN_24;
  assign GEN_26 = 7'h18 == T_534 ? rom_24 : GEN_25;
  assign GEN_27 = 7'h19 == T_534 ? rom_25 : GEN_26;
  assign GEN_28 = 7'h1a == T_534 ? rom_26 : GEN_27;
  assign GEN_29 = 7'h1b == T_534 ? rom_27 : GEN_28;
  assign GEN_30 = 7'h1c == T_534 ? rom_28 : GEN_29;
  assign GEN_31 = 7'h1d == T_534 ? rom_29 : GEN_30;
  assign GEN_32 = 7'h1e == T_534 ? rom_30 : GEN_31;
  assign GEN_33 = 7'h1f == T_534 ? rom_31 : GEN_32;
  assign GEN_34 = 7'h20 == T_534 ? rom_32 : GEN_33;
  assign GEN_35 = 7'h21 == T_534 ? rom_33 : GEN_34;
  assign GEN_36 = 7'h22 == T_534 ? rom_34 : GEN_35;
  assign GEN_37 = 7'h23 == T_534 ? rom_35 : GEN_36;
  assign GEN_38 = 7'h24 == T_534 ? rom_36 : GEN_37;
  assign GEN_39 = 7'h25 == T_534 ? rom_37 : GEN_38;
  assign GEN_40 = 7'h26 == T_534 ? rom_38 : GEN_39;
  assign GEN_41 = 7'h27 == T_534 ? rom_39 : GEN_40;
  assign GEN_42 = 7'h28 == T_534 ? rom_40 : GEN_41;
  assign GEN_43 = 7'h29 == T_534 ? rom_41 : GEN_42;
  assign GEN_44 = 7'h2a == T_534 ? rom_42 : GEN_43;
  assign GEN_45 = 7'h2b == T_534 ? rom_43 : GEN_44;
  assign GEN_46 = 7'h2c == T_534 ? rom_44 : GEN_45;
  assign GEN_47 = 7'h2d == T_534 ? rom_45 : GEN_46;
  assign GEN_48 = 7'h2e == T_534 ? rom_46 : GEN_47;
  assign GEN_49 = 7'h2f == T_534 ? rom_47 : GEN_48;
  assign GEN_50 = 7'h30 == T_534 ? rom_48 : GEN_49;
  assign GEN_51 = 7'h31 == T_534 ? rom_49 : GEN_50;
  assign GEN_52 = 7'h32 == T_534 ? rom_50 : GEN_51;
  assign GEN_53 = 7'h33 == T_534 ? rom_51 : GEN_52;
  assign GEN_54 = 7'h34 == T_534 ? rom_52 : GEN_53;
  assign GEN_55 = 7'h35 == T_534 ? rom_53 : GEN_54;
  assign GEN_56 = 7'h36 == T_534 ? rom_54 : GEN_55;
  assign GEN_57 = 7'h37 == T_534 ? rom_55 : GEN_56;
  assign GEN_58 = 7'h38 == T_534 ? rom_56 : GEN_57;
  assign GEN_59 = 7'h39 == T_534 ? rom_57 : GEN_58;
  assign GEN_60 = 7'h3a == T_534 ? rom_58 : GEN_59;
  assign GEN_61 = 7'h3b == T_534 ? rom_59 : GEN_60;
  assign GEN_62 = 7'h3c == T_534 ? rom_60 : GEN_61;
  assign GEN_63 = 7'h3d == T_534 ? rom_61 : GEN_62;
  assign GEN_64 = 7'h3e == T_534 ? rom_62 : GEN_63;
  assign GEN_65 = 7'h3f == T_534 ? rom_63 : GEN_64;
  assign GEN_66 = 7'h40 == T_534 ? rom_64 : GEN_65;
  assign GEN_67 = 7'h41 == T_534 ? rom_65 : GEN_66;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_68 = {1{$random}};
  addr_beat = GEN_68[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_461) begin
        addr_beat <= io_acquire_bits_addr_beat;
      end else begin
        if(T_457) begin
          addr_beat <= T_460;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported ROMSlave operation\n    at Rom.scala:17 assert(!acq.valid || single_beat || multi_beat, \"unsupported ROMSlave operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module DefaultCoreplex(
  input   clk,
  input   reset,
  input   io_mem_0_acquire_ready,
  output  io_mem_0_acquire_valid,
  output [25:0] io_mem_0_acquire_bits_addr_block,
  output [2:0] io_mem_0_acquire_bits_client_xact_id,
  output [2:0] io_mem_0_acquire_bits_addr_beat,
  output  io_mem_0_acquire_bits_is_builtin_type,
  output [2:0] io_mem_0_acquire_bits_a_type,
  output [10:0] io_mem_0_acquire_bits_union,
  output [63:0] io_mem_0_acquire_bits_data,
  output  io_mem_0_grant_ready,
  input   io_mem_0_grant_valid,
  input  [2:0] io_mem_0_grant_bits_addr_beat,
  input  [2:0] io_mem_0_grant_bits_client_xact_id,
  input   io_mem_0_grant_bits_manager_xact_id,
  input   io_mem_0_grant_bits_is_builtin_type,
  input  [3:0] io_mem_0_grant_bits_g_type,
  input  [63:0] io_mem_0_grant_bits_data,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [33:0] io_debug_req_bits_data,
  input  [1:0] io_debug_req_bits_op,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [33:0] io_debug_resp_bits_data,
  output [1:0] io_debug_resp_bits_resp,
  input   io_rtcTick
);
  wire  tileResets_0;
  wire  tileList_0_clk;
  wire  tileList_0_reset;
  wire  tileList_0_io_cached_0_acquire_ready;
  wire  tileList_0_io_cached_0_acquire_valid;
  wire [25:0] tileList_0_io_cached_0_acquire_bits_addr_block;
  wire [1:0] tileList_0_io_cached_0_acquire_bits_client_xact_id;
  wire [2:0] tileList_0_io_cached_0_acquire_bits_addr_beat;
  wire  tileList_0_io_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] tileList_0_io_cached_0_acquire_bits_a_type;
  wire [10:0] tileList_0_io_cached_0_acquire_bits_union;
  wire [63:0] tileList_0_io_cached_0_acquire_bits_data;
  wire  tileList_0_io_cached_0_probe_ready;
  wire  tileList_0_io_cached_0_probe_valid;
  wire [25:0] tileList_0_io_cached_0_probe_bits_addr_block;
  wire [1:0] tileList_0_io_cached_0_probe_bits_p_type;
  wire  tileList_0_io_cached_0_release_ready;
  wire  tileList_0_io_cached_0_release_valid;
  wire [2:0] tileList_0_io_cached_0_release_bits_addr_beat;
  wire [25:0] tileList_0_io_cached_0_release_bits_addr_block;
  wire [1:0] tileList_0_io_cached_0_release_bits_client_xact_id;
  wire  tileList_0_io_cached_0_release_bits_voluntary;
  wire [2:0] tileList_0_io_cached_0_release_bits_r_type;
  wire [63:0] tileList_0_io_cached_0_release_bits_data;
  wire  tileList_0_io_cached_0_grant_ready;
  wire  tileList_0_io_cached_0_grant_valid;
  wire [2:0] tileList_0_io_cached_0_grant_bits_addr_beat;
  wire [1:0] tileList_0_io_cached_0_grant_bits_client_xact_id;
  wire [2:0] tileList_0_io_cached_0_grant_bits_manager_xact_id;
  wire  tileList_0_io_cached_0_grant_bits_is_builtin_type;
  wire [3:0] tileList_0_io_cached_0_grant_bits_g_type;
  wire [63:0] tileList_0_io_cached_0_grant_bits_data;
  wire  tileList_0_io_cached_0_grant_bits_manager_id;
  wire  tileList_0_io_cached_0_finish_ready;
  wire  tileList_0_io_cached_0_finish_valid;
  wire [2:0] tileList_0_io_cached_0_finish_bits_manager_xact_id;
  wire  tileList_0_io_cached_0_finish_bits_manager_id;
  wire  tileList_0_io_uncached_0_acquire_ready;
  wire  tileList_0_io_uncached_0_acquire_valid;
  wire [25:0] tileList_0_io_uncached_0_acquire_bits_addr_block;
  wire [1:0] tileList_0_io_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] tileList_0_io_uncached_0_acquire_bits_addr_beat;
  wire  tileList_0_io_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] tileList_0_io_uncached_0_acquire_bits_a_type;
  wire [10:0] tileList_0_io_uncached_0_acquire_bits_union;
  wire [63:0] tileList_0_io_uncached_0_acquire_bits_data;
  wire  tileList_0_io_uncached_0_grant_ready;
  wire  tileList_0_io_uncached_0_grant_valid;
  wire [2:0] tileList_0_io_uncached_0_grant_bits_addr_beat;
  wire [1:0] tileList_0_io_uncached_0_grant_bits_client_xact_id;
  wire [2:0] tileList_0_io_uncached_0_grant_bits_manager_xact_id;
  wire  tileList_0_io_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] tileList_0_io_uncached_0_grant_bits_g_type;
  wire [63:0] tileList_0_io_uncached_0_grant_bits_data;
  wire  tileList_0_io_prci_reset;
  wire  tileList_0_io_prci_id;
  wire  tileList_0_io_prci_interrupts_meip;
  wire  tileList_0_io_prci_interrupts_seip;
  wire  tileList_0_io_prci_interrupts_debug;
  wire  tileList_0_io_prci_interrupts_mtip;
  wire  tileList_0_io_prci_interrupts_msip;
  wire  PortedTileLinkCrossbar_1_clk;
  wire  PortedTileLinkCrossbar_1_reset;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat;
  wire [1:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_finish_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_0_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type;
  wire [10:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type;
  wire [3:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_finish_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_finish_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_valid;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type;
  wire  PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_ready;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_valid;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat;
  wire [25:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block;
  wire [1:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary;
  wire [2:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type;
  wire [63:0] PortedTileLinkCrossbar_1_io_managers_1_release_bits_data;
  wire  PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id;
  wire  L2BroadcastHub_1_clk;
  wire  L2BroadcastHub_1_reset;
  wire  L2BroadcastHub_1_io_inner_acquire_ready;
  wire  L2BroadcastHub_1_io_inner_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_inner_acquire_bits_a_type;
  wire [10:0] L2BroadcastHub_1_io_inner_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_inner_acquire_bits_data;
  wire  L2BroadcastHub_1_io_inner_acquire_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_grant_ready;
  wire  L2BroadcastHub_1_io_inner_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  wire [1:0] L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_inner_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_inner_grant_bits_data;
  wire  L2BroadcastHub_1_io_inner_grant_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_finish_ready;
  wire  L2BroadcastHub_1_io_inner_finish_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_inner_probe_ready;
  wire  L2BroadcastHub_1_io_inner_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_inner_probe_bits_client_id;
  wire  L2BroadcastHub_1_io_inner_release_ready;
  wire  L2BroadcastHub_1_io_inner_release_valid;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_inner_release_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_inner_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_inner_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_inner_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_inner_release_bits_data;
  wire  L2BroadcastHub_1_io_inner_release_bits_client_id;
  wire  L2BroadcastHub_1_io_incoherent_0;
  wire  L2BroadcastHub_1_io_outer_acquire_ready;
  wire  L2BroadcastHub_1_io_outer_acquire_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  wire  L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  wire [10:0] L2BroadcastHub_1_io_outer_acquire_bits_union;
  wire [63:0] L2BroadcastHub_1_io_outer_acquire_bits_data;
  wire  L2BroadcastHub_1_io_outer_probe_ready;
  wire  L2BroadcastHub_1_io_outer_probe_valid;
  wire [25:0] L2BroadcastHub_1_io_outer_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_1_io_outer_probe_bits_p_type;
  wire  L2BroadcastHub_1_io_outer_release_ready;
  wire  L2BroadcastHub_1_io_outer_release_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_1_io_outer_release_bits_addr_block;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_1_io_outer_release_bits_r_type;
  wire [63:0] L2BroadcastHub_1_io_outer_release_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_ready;
  wire  L2BroadcastHub_1_io_outer_grant_valid;
  wire [2:0] L2BroadcastHub_1_io_outer_grant_bits_addr_beat;
  wire [2:0] L2BroadcastHub_1_io_outer_grant_bits_client_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_1_io_outer_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_1_io_outer_grant_bits_data;
  wire  L2BroadcastHub_1_io_outer_grant_bits_manager_id;
  wire  L2BroadcastHub_1_io_outer_finish_ready;
  wire  L2BroadcastHub_1_io_outer_finish_valid;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  wire  MMIOTileLinkManager_1_clk;
  wire  MMIOTileLinkManager_1_reset;
  wire  MMIOTileLinkManager_1_io_inner_acquire_ready;
  wire  MMIOTileLinkManager_1_io_inner_acquire_valid;
  wire [25:0] MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat;
  wire  MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] MMIOTileLinkManager_1_io_inner_acquire_bits_a_type;
  wire [10:0] MMIOTileLinkManager_1_io_inner_acquire_bits_union;
  wire [63:0] MMIOTileLinkManager_1_io_inner_acquire_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_acquire_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_grant_ready;
  wire  MMIOTileLinkManager_1_io_inner_grant_valid;
  wire [2:0] MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat;
  wire [1:0] MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] MMIOTileLinkManager_1_io_inner_grant_bits_g_type;
  wire [63:0] MMIOTileLinkManager_1_io_inner_grant_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_grant_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_finish_ready;
  wire  MMIOTileLinkManager_1_io_inner_finish_valid;
  wire [2:0] MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_probe_ready;
  wire  MMIOTileLinkManager_1_io_inner_probe_valid;
  wire [25:0] MMIOTileLinkManager_1_io_inner_probe_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_inner_probe_bits_p_type;
  wire  MMIOTileLinkManager_1_io_inner_probe_bits_client_id;
  wire  MMIOTileLinkManager_1_io_inner_release_ready;
  wire  MMIOTileLinkManager_1_io_inner_release_valid;
  wire [2:0] MMIOTileLinkManager_1_io_inner_release_bits_addr_beat;
  wire [25:0] MMIOTileLinkManager_1_io_inner_release_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id;
  wire  MMIOTileLinkManager_1_io_inner_release_bits_voluntary;
  wire [2:0] MMIOTileLinkManager_1_io_inner_release_bits_r_type;
  wire [63:0] MMIOTileLinkManager_1_io_inner_release_bits_data;
  wire  MMIOTileLinkManager_1_io_inner_release_bits_client_id;
  wire  MMIOTileLinkManager_1_io_incoherent_0;
  wire  MMIOTileLinkManager_1_io_outer_acquire_ready;
  wire  MMIOTileLinkManager_1_io_outer_acquire_valid;
  wire [25:0] MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block;
  wire [1:0] MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat;
  wire  MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] MMIOTileLinkManager_1_io_outer_acquire_bits_a_type;
  wire [10:0] MMIOTileLinkManager_1_io_outer_acquire_bits_union;
  wire [63:0] MMIOTileLinkManager_1_io_outer_acquire_bits_data;
  wire  MMIOTileLinkManager_1_io_outer_grant_ready;
  wire  MMIOTileLinkManager_1_io_outer_grant_valid;
  wire [2:0] MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat;
  wire [1:0] MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id;
  wire  MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id;
  wire  MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] MMIOTileLinkManager_1_io_outer_grant_bits_g_type;
  wire [63:0] MMIOTileLinkManager_1_io_outer_grant_bits_data;
  wire  TileLinkMemoryInterconnect_1_clk;
  wire  TileLinkMemoryInterconnect_1_reset;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_ready;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_ready;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_valid;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat;
  wire [2:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_ready;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_ready;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_valid;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat;
  wire [2:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_clk;
  wire  ClientTileLinkIOUnwrapper_1_reset;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type;
  wire [10:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_valid;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  wire [10:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_clk;
  wire  ClientTileLinkEnqueuer_1_reset;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [10:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [10:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  wire  ClientUncachedTileLinkEnqueuer_1_clk;
  wire  ClientUncachedTileLinkEnqueuer_1_reset;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [10:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_clk;
  wire  TileLinkRecursiveInterconnect_2_reset;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  wire [10:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data;
  wire  PLIC_1_clk;
  wire  PLIC_1_reset;
  wire  PLIC_1_io_devices_0_valid;
  wire  PLIC_1_io_devices_0_ready;
  wire  PLIC_1_io_devices_0_complete;
  wire  PLIC_1_io_devices_1_valid;
  wire  PLIC_1_io_devices_1_ready;
  wire  PLIC_1_io_devices_1_complete;
  wire  PLIC_1_io_harts_0;
  wire  PLIC_1_io_harts_1;
  wire  PLIC_1_io_tl_acquire_ready;
  wire  PLIC_1_io_tl_acquire_valid;
  wire [25:0] PLIC_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PLIC_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PLIC_1_io_tl_acquire_bits_addr_beat;
  wire  PLIC_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PLIC_1_io_tl_acquire_bits_a_type;
  wire [10:0] PLIC_1_io_tl_acquire_bits_union;
  wire [63:0] PLIC_1_io_tl_acquire_bits_data;
  wire  PLIC_1_io_tl_grant_ready;
  wire  PLIC_1_io_tl_grant_valid;
  wire [2:0] PLIC_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PLIC_1_io_tl_grant_bits_client_xact_id;
  wire  PLIC_1_io_tl_grant_bits_manager_xact_id;
  wire  PLIC_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PLIC_1_io_tl_grant_bits_g_type;
  wire [63:0] PLIC_1_io_tl_grant_bits_data;
  wire  LevelGateway_2_clk;
  wire  LevelGateway_2_reset;
  wire  LevelGateway_2_io_interrupt;
  wire  LevelGateway_2_io_plic_valid;
  wire  LevelGateway_2_io_plic_ready;
  wire  LevelGateway_2_io_plic_complete;
  wire  LevelGateway_1_1_clk;
  wire  LevelGateway_1_1_reset;
  wire  LevelGateway_1_1_io_interrupt;
  wire  LevelGateway_1_1_io_plic_valid;
  wire  LevelGateway_1_1_io_plic_ready;
  wire  LevelGateway_1_1_io_plic_complete;
  wire  DebugModule_1_clk;
  wire  DebugModule_1_reset;
  wire  DebugModule_1_io_db_req_ready;
  wire  DebugModule_1_io_db_req_valid;
  wire [4:0] DebugModule_1_io_db_req_bits_addr;
  wire [33:0] DebugModule_1_io_db_req_bits_data;
  wire [1:0] DebugModule_1_io_db_req_bits_op;
  wire  DebugModule_1_io_db_resp_ready;
  wire  DebugModule_1_io_db_resp_valid;
  wire [33:0] DebugModule_1_io_db_resp_bits_data;
  wire [1:0] DebugModule_1_io_db_resp_bits_resp;
  wire  DebugModule_1_io_debugInterrupts_0;
  wire  DebugModule_1_io_tl_acquire_ready;
  wire  DebugModule_1_io_tl_acquire_valid;
  wire [25:0] DebugModule_1_io_tl_acquire_bits_addr_block;
  wire [1:0] DebugModule_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_addr_beat;
  wire  DebugModule_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_a_type;
  wire [10:0] DebugModule_1_io_tl_acquire_bits_union;
  wire [63:0] DebugModule_1_io_tl_acquire_bits_data;
  wire  DebugModule_1_io_tl_grant_ready;
  wire  DebugModule_1_io_tl_grant_valid;
  wire [2:0] DebugModule_1_io_tl_grant_bits_addr_beat;
  wire [1:0] DebugModule_1_io_tl_grant_bits_client_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_manager_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] DebugModule_1_io_tl_grant_bits_g_type;
  wire [63:0] DebugModule_1_io_tl_grant_bits_data;
  wire  DebugModule_1_io_ndreset;
  wire  DebugModule_1_io_fullreset;
  wire  PRCI_1_clk;
  wire  PRCI_1_reset;
  wire  PRCI_1_io_interrupts_0_meip;
  wire  PRCI_1_io_interrupts_0_seip;
  wire  PRCI_1_io_interrupts_0_debug;
  wire  PRCI_1_io_tl_acquire_ready;
  wire  PRCI_1_io_tl_acquire_valid;
  wire [25:0] PRCI_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PRCI_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PRCI_1_io_tl_acquire_bits_addr_beat;
  wire  PRCI_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PRCI_1_io_tl_acquire_bits_a_type;
  wire [10:0] PRCI_1_io_tl_acquire_bits_union;
  wire [63:0] PRCI_1_io_tl_acquire_bits_data;
  wire  PRCI_1_io_tl_grant_ready;
  wire  PRCI_1_io_tl_grant_valid;
  wire [2:0] PRCI_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PRCI_1_io_tl_grant_bits_client_xact_id;
  wire  PRCI_1_io_tl_grant_bits_manager_xact_id;
  wire  PRCI_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PRCI_1_io_tl_grant_bits_g_type;
  wire [63:0] PRCI_1_io_tl_grant_bits_data;
  wire  PRCI_1_io_tiles_0_reset;
  wire  PRCI_1_io_tiles_0_id;
  wire  PRCI_1_io_tiles_0_interrupts_meip;
  wire  PRCI_1_io_tiles_0_interrupts_seip;
  wire  PRCI_1_io_tiles_0_interrupts_debug;
  wire  PRCI_1_io_tiles_0_interrupts_mtip;
  wire  PRCI_1_io_tiles_0_interrupts_msip;
  wire  PRCI_1_io_rtcTick;
  wire  ROMSlave_1_clk;
  wire  ROMSlave_1_reset;
  wire  ROMSlave_1_io_acquire_ready;
  wire  ROMSlave_1_io_acquire_valid;
  wire [25:0] ROMSlave_1_io_acquire_bits_addr_block;
  wire [1:0] ROMSlave_1_io_acquire_bits_client_xact_id;
  wire [2:0] ROMSlave_1_io_acquire_bits_addr_beat;
  wire  ROMSlave_1_io_acquire_bits_is_builtin_type;
  wire [2:0] ROMSlave_1_io_acquire_bits_a_type;
  wire [10:0] ROMSlave_1_io_acquire_bits_union;
  wire [63:0] ROMSlave_1_io_acquire_bits_data;
  wire  ROMSlave_1_io_grant_ready;
  wire  ROMSlave_1_io_grant_valid;
  wire [2:0] ROMSlave_1_io_grant_bits_addr_beat;
  wire [1:0] ROMSlave_1_io_grant_bits_client_xact_id;
  wire  ROMSlave_1_io_grant_bits_manager_xact_id;
  wire  ROMSlave_1_io_grant_bits_is_builtin_type;
  wire [3:0] ROMSlave_1_io_grant_bits_g_type;
  wire [63:0] ROMSlave_1_io_grant_bits_data;
  wire  GEN_0;
  reg [31:0] GEN_1;
  RocketTile tileList_0 (
    .clk(tileList_0_clk),
    .reset(tileList_0_reset),
    .io_cached_0_acquire_ready(tileList_0_io_cached_0_acquire_ready),
    .io_cached_0_acquire_valid(tileList_0_io_cached_0_acquire_valid),
    .io_cached_0_acquire_bits_addr_block(tileList_0_io_cached_0_acquire_bits_addr_block),
    .io_cached_0_acquire_bits_client_xact_id(tileList_0_io_cached_0_acquire_bits_client_xact_id),
    .io_cached_0_acquire_bits_addr_beat(tileList_0_io_cached_0_acquire_bits_addr_beat),
    .io_cached_0_acquire_bits_is_builtin_type(tileList_0_io_cached_0_acquire_bits_is_builtin_type),
    .io_cached_0_acquire_bits_a_type(tileList_0_io_cached_0_acquire_bits_a_type),
    .io_cached_0_acquire_bits_union(tileList_0_io_cached_0_acquire_bits_union),
    .io_cached_0_acquire_bits_data(tileList_0_io_cached_0_acquire_bits_data),
    .io_cached_0_probe_ready(tileList_0_io_cached_0_probe_ready),
    .io_cached_0_probe_valid(tileList_0_io_cached_0_probe_valid),
    .io_cached_0_probe_bits_addr_block(tileList_0_io_cached_0_probe_bits_addr_block),
    .io_cached_0_probe_bits_p_type(tileList_0_io_cached_0_probe_bits_p_type),
    .io_cached_0_release_ready(tileList_0_io_cached_0_release_ready),
    .io_cached_0_release_valid(tileList_0_io_cached_0_release_valid),
    .io_cached_0_release_bits_addr_beat(tileList_0_io_cached_0_release_bits_addr_beat),
    .io_cached_0_release_bits_addr_block(tileList_0_io_cached_0_release_bits_addr_block),
    .io_cached_0_release_bits_client_xact_id(tileList_0_io_cached_0_release_bits_client_xact_id),
    .io_cached_0_release_bits_voluntary(tileList_0_io_cached_0_release_bits_voluntary),
    .io_cached_0_release_bits_r_type(tileList_0_io_cached_0_release_bits_r_type),
    .io_cached_0_release_bits_data(tileList_0_io_cached_0_release_bits_data),
    .io_cached_0_grant_ready(tileList_0_io_cached_0_grant_ready),
    .io_cached_0_grant_valid(tileList_0_io_cached_0_grant_valid),
    .io_cached_0_grant_bits_addr_beat(tileList_0_io_cached_0_grant_bits_addr_beat),
    .io_cached_0_grant_bits_client_xact_id(tileList_0_io_cached_0_grant_bits_client_xact_id),
    .io_cached_0_grant_bits_manager_xact_id(tileList_0_io_cached_0_grant_bits_manager_xact_id),
    .io_cached_0_grant_bits_is_builtin_type(tileList_0_io_cached_0_grant_bits_is_builtin_type),
    .io_cached_0_grant_bits_g_type(tileList_0_io_cached_0_grant_bits_g_type),
    .io_cached_0_grant_bits_data(tileList_0_io_cached_0_grant_bits_data),
    .io_cached_0_grant_bits_manager_id(tileList_0_io_cached_0_grant_bits_manager_id),
    .io_cached_0_finish_ready(tileList_0_io_cached_0_finish_ready),
    .io_cached_0_finish_valid(tileList_0_io_cached_0_finish_valid),
    .io_cached_0_finish_bits_manager_xact_id(tileList_0_io_cached_0_finish_bits_manager_xact_id),
    .io_cached_0_finish_bits_manager_id(tileList_0_io_cached_0_finish_bits_manager_id),
    .io_uncached_0_acquire_ready(tileList_0_io_uncached_0_acquire_ready),
    .io_uncached_0_acquire_valid(tileList_0_io_uncached_0_acquire_valid),
    .io_uncached_0_acquire_bits_addr_block(tileList_0_io_uncached_0_acquire_bits_addr_block),
    .io_uncached_0_acquire_bits_client_xact_id(tileList_0_io_uncached_0_acquire_bits_client_xact_id),
    .io_uncached_0_acquire_bits_addr_beat(tileList_0_io_uncached_0_acquire_bits_addr_beat),
    .io_uncached_0_acquire_bits_is_builtin_type(tileList_0_io_uncached_0_acquire_bits_is_builtin_type),
    .io_uncached_0_acquire_bits_a_type(tileList_0_io_uncached_0_acquire_bits_a_type),
    .io_uncached_0_acquire_bits_union(tileList_0_io_uncached_0_acquire_bits_union),
    .io_uncached_0_acquire_bits_data(tileList_0_io_uncached_0_acquire_bits_data),
    .io_uncached_0_grant_ready(tileList_0_io_uncached_0_grant_ready),
    .io_uncached_0_grant_valid(tileList_0_io_uncached_0_grant_valid),
    .io_uncached_0_grant_bits_addr_beat(tileList_0_io_uncached_0_grant_bits_addr_beat),
    .io_uncached_0_grant_bits_client_xact_id(tileList_0_io_uncached_0_grant_bits_client_xact_id),
    .io_uncached_0_grant_bits_manager_xact_id(tileList_0_io_uncached_0_grant_bits_manager_xact_id),
    .io_uncached_0_grant_bits_is_builtin_type(tileList_0_io_uncached_0_grant_bits_is_builtin_type),
    .io_uncached_0_grant_bits_g_type(tileList_0_io_uncached_0_grant_bits_g_type),
    .io_uncached_0_grant_bits_data(tileList_0_io_uncached_0_grant_bits_data),
    .io_prci_reset(tileList_0_io_prci_reset),
    .io_prci_id(tileList_0_io_prci_id),
    .io_prci_interrupts_meip(tileList_0_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(tileList_0_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(tileList_0_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(tileList_0_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(tileList_0_io_prci_interrupts_msip)
  );
  PortedTileLinkCrossbar PortedTileLinkCrossbar_1 (
    .clk(PortedTileLinkCrossbar_1_clk),
    .reset(PortedTileLinkCrossbar_1_reset),
    .io_clients_cached_0_acquire_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready),
    .io_clients_cached_0_acquire_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid),
    .io_clients_cached_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block),
    .io_clients_cached_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id),
    .io_clients_cached_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat),
    .io_clients_cached_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type),
    .io_clients_cached_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type),
    .io_clients_cached_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union),
    .io_clients_cached_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data),
    .io_clients_cached_0_probe_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready),
    .io_clients_cached_0_probe_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid),
    .io_clients_cached_0_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block),
    .io_clients_cached_0_probe_bits_p_type(PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type),
    .io_clients_cached_0_release_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready),
    .io_clients_cached_0_release_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid),
    .io_clients_cached_0_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat),
    .io_clients_cached_0_release_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block),
    .io_clients_cached_0_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id),
    .io_clients_cached_0_release_bits_voluntary(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary),
    .io_clients_cached_0_release_bits_r_type(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type),
    .io_clients_cached_0_release_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data),
    .io_clients_cached_0_grant_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready),
    .io_clients_cached_0_grant_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid),
    .io_clients_cached_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat),
    .io_clients_cached_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id),
    .io_clients_cached_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id),
    .io_clients_cached_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type),
    .io_clients_cached_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type),
    .io_clients_cached_0_grant_bits_data(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data),
    .io_clients_cached_0_grant_bits_manager_id(PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id),
    .io_clients_cached_0_finish_ready(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready),
    .io_clients_cached_0_finish_valid(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid),
    .io_clients_cached_0_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id),
    .io_clients_cached_0_finish_bits_manager_id(PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id),
    .io_clients_uncached_0_acquire_ready(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready),
    .io_clients_uncached_0_acquire_valid(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid),
    .io_clients_uncached_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block),
    .io_clients_uncached_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id),
    .io_clients_uncached_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat),
    .io_clients_uncached_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type),
    .io_clients_uncached_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type),
    .io_clients_uncached_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union),
    .io_clients_uncached_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data),
    .io_clients_uncached_0_grant_ready(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready),
    .io_clients_uncached_0_grant_valid(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid),
    .io_clients_uncached_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat),
    .io_clients_uncached_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id),
    .io_clients_uncached_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id),
    .io_clients_uncached_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type),
    .io_clients_uncached_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type),
    .io_clients_uncached_0_grant_bits_data(PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data),
    .io_managers_0_acquire_ready(PortedTileLinkCrossbar_1_io_managers_0_acquire_ready),
    .io_managers_0_acquire_valid(PortedTileLinkCrossbar_1_io_managers_0_acquire_valid),
    .io_managers_0_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block),
    .io_managers_0_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id),
    .io_managers_0_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat),
    .io_managers_0_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type),
    .io_managers_0_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type),
    .io_managers_0_acquire_bits_union(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union),
    .io_managers_0_acquire_bits_data(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data),
    .io_managers_0_acquire_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id),
    .io_managers_0_grant_ready(PortedTileLinkCrossbar_1_io_managers_0_grant_ready),
    .io_managers_0_grant_valid(PortedTileLinkCrossbar_1_io_managers_0_grant_valid),
    .io_managers_0_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat),
    .io_managers_0_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id),
    .io_managers_0_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id),
    .io_managers_0_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type),
    .io_managers_0_grant_bits_g_type(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type),
    .io_managers_0_grant_bits_data(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data),
    .io_managers_0_grant_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id),
    .io_managers_0_finish_ready(PortedTileLinkCrossbar_1_io_managers_0_finish_ready),
    .io_managers_0_finish_valid(PortedTileLinkCrossbar_1_io_managers_0_finish_valid),
    .io_managers_0_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id),
    .io_managers_0_probe_ready(PortedTileLinkCrossbar_1_io_managers_0_probe_ready),
    .io_managers_0_probe_valid(PortedTileLinkCrossbar_1_io_managers_0_probe_valid),
    .io_managers_0_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block),
    .io_managers_0_probe_bits_p_type(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type),
    .io_managers_0_probe_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id),
    .io_managers_0_release_ready(PortedTileLinkCrossbar_1_io_managers_0_release_ready),
    .io_managers_0_release_valid(PortedTileLinkCrossbar_1_io_managers_0_release_valid),
    .io_managers_0_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat),
    .io_managers_0_release_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block),
    .io_managers_0_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id),
    .io_managers_0_release_bits_voluntary(PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary),
    .io_managers_0_release_bits_r_type(PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type),
    .io_managers_0_release_bits_data(PortedTileLinkCrossbar_1_io_managers_0_release_bits_data),
    .io_managers_0_release_bits_client_id(PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id),
    .io_managers_1_acquire_ready(PortedTileLinkCrossbar_1_io_managers_1_acquire_ready),
    .io_managers_1_acquire_valid(PortedTileLinkCrossbar_1_io_managers_1_acquire_valid),
    .io_managers_1_acquire_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block),
    .io_managers_1_acquire_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id),
    .io_managers_1_acquire_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat),
    .io_managers_1_acquire_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type),
    .io_managers_1_acquire_bits_a_type(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type),
    .io_managers_1_acquire_bits_union(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union),
    .io_managers_1_acquire_bits_data(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data),
    .io_managers_1_acquire_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id),
    .io_managers_1_grant_ready(PortedTileLinkCrossbar_1_io_managers_1_grant_ready),
    .io_managers_1_grant_valid(PortedTileLinkCrossbar_1_io_managers_1_grant_valid),
    .io_managers_1_grant_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat),
    .io_managers_1_grant_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id),
    .io_managers_1_grant_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id),
    .io_managers_1_grant_bits_is_builtin_type(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type),
    .io_managers_1_grant_bits_g_type(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type),
    .io_managers_1_grant_bits_data(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data),
    .io_managers_1_grant_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id),
    .io_managers_1_finish_ready(PortedTileLinkCrossbar_1_io_managers_1_finish_ready),
    .io_managers_1_finish_valid(PortedTileLinkCrossbar_1_io_managers_1_finish_valid),
    .io_managers_1_finish_bits_manager_xact_id(PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id),
    .io_managers_1_probe_ready(PortedTileLinkCrossbar_1_io_managers_1_probe_ready),
    .io_managers_1_probe_valid(PortedTileLinkCrossbar_1_io_managers_1_probe_valid),
    .io_managers_1_probe_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block),
    .io_managers_1_probe_bits_p_type(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type),
    .io_managers_1_probe_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id),
    .io_managers_1_release_ready(PortedTileLinkCrossbar_1_io_managers_1_release_ready),
    .io_managers_1_release_valid(PortedTileLinkCrossbar_1_io_managers_1_release_valid),
    .io_managers_1_release_bits_addr_beat(PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat),
    .io_managers_1_release_bits_addr_block(PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block),
    .io_managers_1_release_bits_client_xact_id(PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id),
    .io_managers_1_release_bits_voluntary(PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary),
    .io_managers_1_release_bits_r_type(PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type),
    .io_managers_1_release_bits_data(PortedTileLinkCrossbar_1_io_managers_1_release_bits_data),
    .io_managers_1_release_bits_client_id(PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id)
  );
  L2BroadcastHub L2BroadcastHub_1 (
    .clk(L2BroadcastHub_1_clk),
    .reset(L2BroadcastHub_1_reset),
    .io_inner_acquire_ready(L2BroadcastHub_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(L2BroadcastHub_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(L2BroadcastHub_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(L2BroadcastHub_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(L2BroadcastHub_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(L2BroadcastHub_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(L2BroadcastHub_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(L2BroadcastHub_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(L2BroadcastHub_1_io_inner_grant_ready),
    .io_inner_grant_valid(L2BroadcastHub_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(L2BroadcastHub_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(L2BroadcastHub_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(L2BroadcastHub_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(L2BroadcastHub_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(L2BroadcastHub_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(L2BroadcastHub_1_io_inner_finish_ready),
    .io_inner_finish_valid(L2BroadcastHub_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(L2BroadcastHub_1_io_inner_probe_ready),
    .io_inner_probe_valid(L2BroadcastHub_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(L2BroadcastHub_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(L2BroadcastHub_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(L2BroadcastHub_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(L2BroadcastHub_1_io_inner_release_ready),
    .io_inner_release_valid(L2BroadcastHub_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(L2BroadcastHub_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(L2BroadcastHub_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(L2BroadcastHub_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(L2BroadcastHub_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(L2BroadcastHub_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(L2BroadcastHub_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(L2BroadcastHub_1_io_inner_release_bits_client_id),
    .io_incoherent_0(L2BroadcastHub_1_io_incoherent_0),
    .io_outer_acquire_ready(L2BroadcastHub_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(L2BroadcastHub_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(L2BroadcastHub_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(L2BroadcastHub_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(L2BroadcastHub_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(L2BroadcastHub_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(L2BroadcastHub_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(L2BroadcastHub_1_io_outer_probe_ready),
    .io_outer_probe_valid(L2BroadcastHub_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(L2BroadcastHub_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(L2BroadcastHub_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(L2BroadcastHub_1_io_outer_release_ready),
    .io_outer_release_valid(L2BroadcastHub_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(L2BroadcastHub_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(L2BroadcastHub_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(L2BroadcastHub_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(L2BroadcastHub_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(L2BroadcastHub_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(L2BroadcastHub_1_io_outer_release_bits_data),
    .io_outer_grant_ready(L2BroadcastHub_1_io_outer_grant_ready),
    .io_outer_grant_valid(L2BroadcastHub_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(L2BroadcastHub_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(L2BroadcastHub_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(L2BroadcastHub_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(L2BroadcastHub_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(L2BroadcastHub_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(L2BroadcastHub_1_io_outer_finish_ready),
    .io_outer_finish_valid(L2BroadcastHub_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(L2BroadcastHub_1_io_outer_finish_bits_manager_id)
  );
  MMIOTileLinkManager MMIOTileLinkManager_1 (
    .clk(MMIOTileLinkManager_1_clk),
    .reset(MMIOTileLinkManager_1_reset),
    .io_inner_acquire_ready(MMIOTileLinkManager_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(MMIOTileLinkManager_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(MMIOTileLinkManager_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(MMIOTileLinkManager_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(MMIOTileLinkManager_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(MMIOTileLinkManager_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(MMIOTileLinkManager_1_io_inner_grant_ready),
    .io_inner_grant_valid(MMIOTileLinkManager_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(MMIOTileLinkManager_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(MMIOTileLinkManager_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(MMIOTileLinkManager_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(MMIOTileLinkManager_1_io_inner_finish_ready),
    .io_inner_finish_valid(MMIOTileLinkManager_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(MMIOTileLinkManager_1_io_inner_probe_ready),
    .io_inner_probe_valid(MMIOTileLinkManager_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(MMIOTileLinkManager_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(MMIOTileLinkManager_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(MMIOTileLinkManager_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(MMIOTileLinkManager_1_io_inner_release_ready),
    .io_inner_release_valid(MMIOTileLinkManager_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(MMIOTileLinkManager_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(MMIOTileLinkManager_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(MMIOTileLinkManager_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(MMIOTileLinkManager_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(MMIOTileLinkManager_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(MMIOTileLinkManager_1_io_inner_release_bits_client_id),
    .io_incoherent_0(MMIOTileLinkManager_1_io_incoherent_0),
    .io_outer_acquire_ready(MMIOTileLinkManager_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(MMIOTileLinkManager_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(MMIOTileLinkManager_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(MMIOTileLinkManager_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(MMIOTileLinkManager_1_io_outer_acquire_bits_data),
    .io_outer_grant_ready(MMIOTileLinkManager_1_io_outer_grant_ready),
    .io_outer_grant_valid(MMIOTileLinkManager_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(MMIOTileLinkManager_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(MMIOTileLinkManager_1_io_outer_grant_bits_data)
  );
  TileLinkMemoryInterconnect TileLinkMemoryInterconnect_1 (
    .clk(TileLinkMemoryInterconnect_1_clk),
    .reset(TileLinkMemoryInterconnect_1_reset),
    .io_in_0_acquire_ready(TileLinkMemoryInterconnect_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkMemoryInterconnect_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkMemoryInterconnect_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkMemoryInterconnect_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkMemoryInterconnect_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkMemoryInterconnect_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkMemoryInterconnect_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkMemoryInterconnect_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data)
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper_1 (
    .clk(ClientTileLinkIOUnwrapper_1_clk),
    .reset(ClientTileLinkIOUnwrapper_1_reset),
    .io_in_acquire_ready(ClientTileLinkIOUnwrapper_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOUnwrapper_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data),
    .io_in_probe_ready(ClientTileLinkIOUnwrapper_1_io_in_probe_ready),
    .io_in_probe_valid(ClientTileLinkIOUnwrapper_1_io_in_probe_valid),
    .io_in_probe_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block),
    .io_in_probe_bits_p_type(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type),
    .io_in_release_ready(ClientTileLinkIOUnwrapper_1_io_in_release_ready),
    .io_in_release_valid(ClientTileLinkIOUnwrapper_1_io_in_release_valid),
    .io_in_release_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat),
    .io_in_release_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block),
    .io_in_release_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id),
    .io_in_release_bits_voluntary(ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary),
    .io_in_release_bits_r_type(ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type),
    .io_in_release_bits_data(ClientTileLinkIOUnwrapper_1_io_in_release_bits_data),
    .io_in_grant_ready(ClientTileLinkIOUnwrapper_1_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOUnwrapper_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data),
    .io_in_grant_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id),
    .io_in_finish_ready(ClientTileLinkIOUnwrapper_1_io_in_finish_ready),
    .io_in_finish_valid(ClientTileLinkIOUnwrapper_1_io_in_finish_valid),
    .io_in_finish_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id),
    .io_in_finish_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id),
    .io_out_acquire_ready(ClientTileLinkIOUnwrapper_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOUnwrapper_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientTileLinkIOUnwrapper_1_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOUnwrapper_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data)
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer_1 (
    .clk(ClientTileLinkEnqueuer_1_clk),
    .reset(ClientTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_probe_ready(ClientTileLinkEnqueuer_1_io_inner_probe_ready),
    .io_inner_probe_valid(ClientTileLinkEnqueuer_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type),
    .io_inner_release_ready(ClientTileLinkEnqueuer_1_io_inner_release_ready),
    .io_inner_release_valid(ClientTileLinkEnqueuer_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ClientTileLinkEnqueuer_1_io_inner_release_bits_data),
    .io_inner_grant_ready(ClientTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id),
    .io_inner_finish_ready(ClientTileLinkEnqueuer_1_io_inner_finish_ready),
    .io_inner_finish_valid(ClientTileLinkEnqueuer_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id),
    .io_outer_acquire_ready(ClientTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ClientTileLinkEnqueuer_1_io_outer_probe_ready),
    .io_outer_probe_valid(ClientTileLinkEnqueuer_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ClientTileLinkEnqueuer_1_io_outer_release_ready),
    .io_outer_release_valid(ClientTileLinkEnqueuer_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ClientTileLinkEnqueuer_1_io_outer_release_bits_data),
    .io_outer_grant_ready(ClientTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientTileLinkEnqueuer_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ClientTileLinkEnqueuer_1_io_outer_finish_ready),
    .io_outer_finish_valid(ClientTileLinkEnqueuer_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id)
  );
  ClientUncachedTileLinkEnqueuer ClientUncachedTileLinkEnqueuer_1 (
    .clk(ClientUncachedTileLinkEnqueuer_1_clk),
    .reset(ClientUncachedTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_grant_ready(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_outer_acquire_ready(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_grant_ready(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data)
  );
  TileLinkRecursiveInterconnect TileLinkRecursiveInterconnect_2 (
    .clk(TileLinkRecursiveInterconnect_2_clk),
    .reset(TileLinkRecursiveInterconnect_2_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_2_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_2_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_2_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_2_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_2_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_2_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_2_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_2_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_2_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_2_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data)
  );
  PLIC PLIC_1 (
    .clk(PLIC_1_clk),
    .reset(PLIC_1_reset),
    .io_devices_0_valid(PLIC_1_io_devices_0_valid),
    .io_devices_0_ready(PLIC_1_io_devices_0_ready),
    .io_devices_0_complete(PLIC_1_io_devices_0_complete),
    .io_devices_1_valid(PLIC_1_io_devices_1_valid),
    .io_devices_1_ready(PLIC_1_io_devices_1_ready),
    .io_devices_1_complete(PLIC_1_io_devices_1_complete),
    .io_harts_0(PLIC_1_io_harts_0),
    .io_harts_1(PLIC_1_io_harts_1),
    .io_tl_acquire_ready(PLIC_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PLIC_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PLIC_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PLIC_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PLIC_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PLIC_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PLIC_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PLIC_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PLIC_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PLIC_1_io_tl_grant_ready),
    .io_tl_grant_valid(PLIC_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PLIC_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PLIC_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PLIC_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PLIC_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PLIC_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PLIC_1_io_tl_grant_bits_data)
  );
  LevelGateway LevelGateway_2 (
    .clk(LevelGateway_2_clk),
    .reset(LevelGateway_2_reset),
    .io_interrupt(LevelGateway_2_io_interrupt),
    .io_plic_valid(LevelGateway_2_io_plic_valid),
    .io_plic_ready(LevelGateway_2_io_plic_ready),
    .io_plic_complete(LevelGateway_2_io_plic_complete)
  );
  LevelGateway LevelGateway_1_1 (
    .clk(LevelGateway_1_1_clk),
    .reset(LevelGateway_1_1_reset),
    .io_interrupt(LevelGateway_1_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_1_io_plic_complete)
  );
  DebugModule DebugModule_1 (
    .clk(DebugModule_1_clk),
    .reset(DebugModule_1_reset),
    .io_db_req_ready(DebugModule_1_io_db_req_ready),
    .io_db_req_valid(DebugModule_1_io_db_req_valid),
    .io_db_req_bits_addr(DebugModule_1_io_db_req_bits_addr),
    .io_db_req_bits_data(DebugModule_1_io_db_req_bits_data),
    .io_db_req_bits_op(DebugModule_1_io_db_req_bits_op),
    .io_db_resp_ready(DebugModule_1_io_db_resp_ready),
    .io_db_resp_valid(DebugModule_1_io_db_resp_valid),
    .io_db_resp_bits_data(DebugModule_1_io_db_resp_bits_data),
    .io_db_resp_bits_resp(DebugModule_1_io_db_resp_bits_resp),
    .io_debugInterrupts_0(DebugModule_1_io_debugInterrupts_0),
    .io_tl_acquire_ready(DebugModule_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(DebugModule_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(DebugModule_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(DebugModule_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(DebugModule_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(DebugModule_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(DebugModule_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(DebugModule_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(DebugModule_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(DebugModule_1_io_tl_grant_ready),
    .io_tl_grant_valid(DebugModule_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(DebugModule_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(DebugModule_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(DebugModule_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(DebugModule_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(DebugModule_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(DebugModule_1_io_tl_grant_bits_data),
    .io_ndreset(DebugModule_1_io_ndreset),
    .io_fullreset(DebugModule_1_io_fullreset)
  );
  PRCI PRCI_1 (
    .clk(PRCI_1_clk),
    .reset(PRCI_1_reset),
    .io_interrupts_0_meip(PRCI_1_io_interrupts_0_meip),
    .io_interrupts_0_seip(PRCI_1_io_interrupts_0_seip),
    .io_interrupts_0_debug(PRCI_1_io_interrupts_0_debug),
    .io_tl_acquire_ready(PRCI_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PRCI_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PRCI_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PRCI_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PRCI_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PRCI_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PRCI_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PRCI_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PRCI_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PRCI_1_io_tl_grant_ready),
    .io_tl_grant_valid(PRCI_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PRCI_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PRCI_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PRCI_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PRCI_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PRCI_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PRCI_1_io_tl_grant_bits_data),
    .io_tiles_0_reset(PRCI_1_io_tiles_0_reset),
    .io_tiles_0_id(PRCI_1_io_tiles_0_id),
    .io_tiles_0_interrupts_meip(PRCI_1_io_tiles_0_interrupts_meip),
    .io_tiles_0_interrupts_seip(PRCI_1_io_tiles_0_interrupts_seip),
    .io_tiles_0_interrupts_debug(PRCI_1_io_tiles_0_interrupts_debug),
    .io_tiles_0_interrupts_mtip(PRCI_1_io_tiles_0_interrupts_mtip),
    .io_tiles_0_interrupts_msip(PRCI_1_io_tiles_0_interrupts_msip),
    .io_rtcTick(PRCI_1_io_rtcTick)
  );
  ROMSlave ROMSlave_1 (
    .clk(ROMSlave_1_clk),
    .reset(ROMSlave_1_reset),
    .io_acquire_ready(ROMSlave_1_io_acquire_ready),
    .io_acquire_valid(ROMSlave_1_io_acquire_valid),
    .io_acquire_bits_addr_block(ROMSlave_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(ROMSlave_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(ROMSlave_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(ROMSlave_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(ROMSlave_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(ROMSlave_1_io_acquire_bits_union),
    .io_acquire_bits_data(ROMSlave_1_io_acquire_bits_data),
    .io_grant_ready(ROMSlave_1_io_grant_ready),
    .io_grant_valid(ROMSlave_1_io_grant_valid),
    .io_grant_bits_addr_beat(ROMSlave_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(ROMSlave_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(ROMSlave_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(ROMSlave_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(ROMSlave_1_io_grant_bits_g_type),
    .io_grant_bits_data(ROMSlave_1_io_grant_bits_data)
  );
  assign io_mem_0_acquire_valid = TileLinkMemoryInterconnect_1_io_out_0_acquire_valid;
  assign io_mem_0_acquire_bits_addr_block = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_block;
  assign io_mem_0_acquire_bits_client_xact_id = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_client_xact_id;
  assign io_mem_0_acquire_bits_addr_beat = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_addr_beat;
  assign io_mem_0_acquire_bits_is_builtin_type = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_mem_0_acquire_bits_a_type = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_a_type;
  assign io_mem_0_acquire_bits_union = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_union;
  assign io_mem_0_acquire_bits_data = TileLinkMemoryInterconnect_1_io_out_0_acquire_bits_data;
  assign io_mem_0_grant_ready = TileLinkMemoryInterconnect_1_io_out_0_grant_ready;
  assign io_debug_req_ready = DebugModule_1_io_db_req_ready;
  assign io_debug_resp_valid = DebugModule_1_io_db_resp_valid;
  assign io_debug_resp_bits_data = DebugModule_1_io_db_resp_bits_data;
  assign io_debug_resp_bits_resp = DebugModule_1_io_db_resp_bits_resp;
  assign tileResets_0 = reset;
  assign tileList_0_clk = clk;
  assign tileList_0_reset = tileResets_0;
  assign tileList_0_io_cached_0_acquire_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_ready;
  assign tileList_0_io_cached_0_probe_valid = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_valid;
  assign tileList_0_io_cached_0_probe_bits_addr_block = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_addr_block;
  assign tileList_0_io_cached_0_probe_bits_p_type = PortedTileLinkCrossbar_1_io_clients_cached_0_probe_bits_p_type;
  assign tileList_0_io_cached_0_release_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_release_ready;
  assign tileList_0_io_cached_0_grant_valid = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_valid;
  assign tileList_0_io_cached_0_grant_bits_addr_beat = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_addr_beat;
  assign tileList_0_io_cached_0_grant_bits_client_xact_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_client_xact_id;
  assign tileList_0_io_cached_0_grant_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_xact_id;
  assign tileList_0_io_cached_0_grant_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_is_builtin_type;
  assign tileList_0_io_cached_0_grant_bits_g_type = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_g_type;
  assign tileList_0_io_cached_0_grant_bits_data = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_data;
  assign tileList_0_io_cached_0_grant_bits_manager_id = PortedTileLinkCrossbar_1_io_clients_cached_0_grant_bits_manager_id;
  assign tileList_0_io_cached_0_finish_ready = PortedTileLinkCrossbar_1_io_clients_cached_0_finish_ready;
  assign tileList_0_io_uncached_0_acquire_ready = PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_ready;
  assign tileList_0_io_uncached_0_grant_valid = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_valid;
  assign tileList_0_io_uncached_0_grant_bits_addr_beat = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_addr_beat;
  assign tileList_0_io_uncached_0_grant_bits_client_xact_id = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_client_xact_id;
  assign tileList_0_io_uncached_0_grant_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_manager_xact_id;
  assign tileList_0_io_uncached_0_grant_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_is_builtin_type;
  assign tileList_0_io_uncached_0_grant_bits_g_type = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_g_type;
  assign tileList_0_io_uncached_0_grant_bits_data = PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_bits_data;
  assign tileList_0_io_prci_reset = PRCI_1_io_tiles_0_reset;
  assign tileList_0_io_prci_id = PRCI_1_io_tiles_0_id;
  assign tileList_0_io_prci_interrupts_meip = PRCI_1_io_tiles_0_interrupts_meip;
  assign tileList_0_io_prci_interrupts_seip = PRCI_1_io_tiles_0_interrupts_seip;
  assign tileList_0_io_prci_interrupts_debug = PRCI_1_io_tiles_0_interrupts_debug;
  assign tileList_0_io_prci_interrupts_mtip = PRCI_1_io_tiles_0_interrupts_mtip;
  assign tileList_0_io_prci_interrupts_msip = PRCI_1_io_tiles_0_interrupts_msip;
  assign PortedTileLinkCrossbar_1_clk = clk;
  assign PortedTileLinkCrossbar_1_reset = reset;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_valid = tileList_0_io_cached_0_acquire_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_block = tileList_0_io_cached_0_acquire_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_client_xact_id = tileList_0_io_cached_0_acquire_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_addr_beat = tileList_0_io_cached_0_acquire_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_is_builtin_type = tileList_0_io_cached_0_acquire_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_a_type = tileList_0_io_cached_0_acquire_bits_a_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_union = tileList_0_io_cached_0_acquire_bits_union;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_acquire_bits_data = tileList_0_io_cached_0_acquire_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_probe_ready = tileList_0_io_cached_0_probe_ready;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_valid = tileList_0_io_cached_0_release_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_beat = tileList_0_io_cached_0_release_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_addr_block = tileList_0_io_cached_0_release_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_client_xact_id = tileList_0_io_cached_0_release_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_voluntary = tileList_0_io_cached_0_release_bits_voluntary;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_r_type = tileList_0_io_cached_0_release_bits_r_type;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_release_bits_data = tileList_0_io_cached_0_release_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_grant_ready = tileList_0_io_cached_0_grant_ready;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_valid = tileList_0_io_cached_0_finish_valid;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_xact_id = tileList_0_io_cached_0_finish_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_cached_0_finish_bits_manager_id = tileList_0_io_cached_0_finish_bits_manager_id;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_valid = tileList_0_io_uncached_0_acquire_valid;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_block = tileList_0_io_uncached_0_acquire_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_client_xact_id = tileList_0_io_uncached_0_acquire_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_addr_beat = tileList_0_io_uncached_0_acquire_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_is_builtin_type = tileList_0_io_uncached_0_acquire_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_a_type = tileList_0_io_uncached_0_acquire_bits_a_type;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_union = tileList_0_io_uncached_0_acquire_bits_union;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_acquire_bits_data = tileList_0_io_uncached_0_acquire_bits_data;
  assign PortedTileLinkCrossbar_1_io_clients_uncached_0_grant_ready = tileList_0_io_uncached_0_grant_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_acquire_ready = L2BroadcastHub_1_io_inner_acquire_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_valid = L2BroadcastHub_1_io_inner_grant_valid;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_addr_beat = L2BroadcastHub_1_io_inner_grant_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_xact_id = L2BroadcastHub_1_io_inner_grant_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_manager_xact_id = L2BroadcastHub_1_io_inner_grant_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_is_builtin_type = L2BroadcastHub_1_io_inner_grant_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_g_type = L2BroadcastHub_1_io_inner_grant_bits_g_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_data = L2BroadcastHub_1_io_inner_grant_bits_data;
  assign PortedTileLinkCrossbar_1_io_managers_0_grant_bits_client_id = L2BroadcastHub_1_io_inner_grant_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_finish_ready = L2BroadcastHub_1_io_inner_finish_ready;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_valid = L2BroadcastHub_1_io_inner_probe_valid;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_addr_block = L2BroadcastHub_1_io_inner_probe_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_p_type = L2BroadcastHub_1_io_inner_probe_bits_p_type;
  assign PortedTileLinkCrossbar_1_io_managers_0_probe_bits_client_id = L2BroadcastHub_1_io_inner_probe_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_0_release_ready = L2BroadcastHub_1_io_inner_release_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_acquire_ready = MMIOTileLinkManager_1_io_inner_acquire_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_valid = MMIOTileLinkManager_1_io_inner_grant_valid;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_addr_beat = MMIOTileLinkManager_1_io_inner_grant_bits_addr_beat;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_xact_id = MMIOTileLinkManager_1_io_inner_grant_bits_client_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_manager_xact_id = MMIOTileLinkManager_1_io_inner_grant_bits_manager_xact_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_is_builtin_type = MMIOTileLinkManager_1_io_inner_grant_bits_is_builtin_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_g_type = MMIOTileLinkManager_1_io_inner_grant_bits_g_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_data = MMIOTileLinkManager_1_io_inner_grant_bits_data;
  assign PortedTileLinkCrossbar_1_io_managers_1_grant_bits_client_id = MMIOTileLinkManager_1_io_inner_grant_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_finish_ready = MMIOTileLinkManager_1_io_inner_finish_ready;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_valid = MMIOTileLinkManager_1_io_inner_probe_valid;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_addr_block = MMIOTileLinkManager_1_io_inner_probe_bits_addr_block;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_p_type = MMIOTileLinkManager_1_io_inner_probe_bits_p_type;
  assign PortedTileLinkCrossbar_1_io_managers_1_probe_bits_client_id = MMIOTileLinkManager_1_io_inner_probe_bits_client_id;
  assign PortedTileLinkCrossbar_1_io_managers_1_release_ready = MMIOTileLinkManager_1_io_inner_release_ready;
  assign L2BroadcastHub_1_clk = clk;
  assign L2BroadcastHub_1_reset = reset;
  assign L2BroadcastHub_1_io_inner_acquire_valid = PortedTileLinkCrossbar_1_io_managers_0_acquire_valid;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_acquire_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_acquire_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_a_type = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_a_type;
  assign L2BroadcastHub_1_io_inner_acquire_bits_union = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_union;
  assign L2BroadcastHub_1_io_inner_acquire_bits_data = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_data;
  assign L2BroadcastHub_1_io_inner_acquire_bits_client_id = PortedTileLinkCrossbar_1_io_managers_0_acquire_bits_client_id;
  assign L2BroadcastHub_1_io_inner_grant_ready = PortedTileLinkCrossbar_1_io_managers_0_grant_ready;
  assign L2BroadcastHub_1_io_inner_finish_valid = PortedTileLinkCrossbar_1_io_managers_0_finish_valid;
  assign L2BroadcastHub_1_io_inner_finish_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_managers_0_finish_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_inner_probe_ready = PortedTileLinkCrossbar_1_io_managers_0_probe_ready;
  assign L2BroadcastHub_1_io_inner_release_valid = PortedTileLinkCrossbar_1_io_managers_0_release_valid;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_beat;
  assign L2BroadcastHub_1_io_inner_release_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_0_release_bits_addr_block;
  assign L2BroadcastHub_1_io_inner_release_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_xact_id;
  assign L2BroadcastHub_1_io_inner_release_bits_voluntary = PortedTileLinkCrossbar_1_io_managers_0_release_bits_voluntary;
  assign L2BroadcastHub_1_io_inner_release_bits_r_type = PortedTileLinkCrossbar_1_io_managers_0_release_bits_r_type;
  assign L2BroadcastHub_1_io_inner_release_bits_data = PortedTileLinkCrossbar_1_io_managers_0_release_bits_data;
  assign L2BroadcastHub_1_io_inner_release_bits_client_id = PortedTileLinkCrossbar_1_io_managers_0_release_bits_client_id;
  assign L2BroadcastHub_1_io_incoherent_0 = 1'h0;
  assign L2BroadcastHub_1_io_outer_acquire_ready = ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign L2BroadcastHub_1_io_outer_probe_valid = ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  assign L2BroadcastHub_1_io_outer_probe_bits_addr_block = ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  assign L2BroadcastHub_1_io_outer_probe_bits_p_type = ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  assign L2BroadcastHub_1_io_outer_release_ready = ClientTileLinkEnqueuer_1_io_inner_release_ready;
  assign L2BroadcastHub_1_io_outer_grant_valid = ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  assign L2BroadcastHub_1_io_outer_grant_bits_addr_beat = ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign L2BroadcastHub_1_io_outer_grant_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  assign L2BroadcastHub_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_g_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign L2BroadcastHub_1_io_outer_grant_bits_data = ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign L2BroadcastHub_1_io_outer_grant_bits_manager_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  assign L2BroadcastHub_1_io_outer_finish_ready = ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  assign MMIOTileLinkManager_1_clk = clk;
  assign MMIOTileLinkManager_1_reset = reset;
  assign MMIOTileLinkManager_1_io_inner_acquire_valid = PortedTileLinkCrossbar_1_io_managers_1_acquire_valid;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_block;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_xact_id;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_is_builtin_type = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_is_builtin_type;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_a_type = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_a_type;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_union = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_union;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_data = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_data;
  assign MMIOTileLinkManager_1_io_inner_acquire_bits_client_id = PortedTileLinkCrossbar_1_io_managers_1_acquire_bits_client_id;
  assign MMIOTileLinkManager_1_io_inner_grant_ready = PortedTileLinkCrossbar_1_io_managers_1_grant_ready;
  assign MMIOTileLinkManager_1_io_inner_finish_valid = PortedTileLinkCrossbar_1_io_managers_1_finish_valid;
  assign MMIOTileLinkManager_1_io_inner_finish_bits_manager_xact_id = PortedTileLinkCrossbar_1_io_managers_1_finish_bits_manager_xact_id;
  assign MMIOTileLinkManager_1_io_inner_probe_ready = PortedTileLinkCrossbar_1_io_managers_1_probe_ready;
  assign MMIOTileLinkManager_1_io_inner_release_valid = PortedTileLinkCrossbar_1_io_managers_1_release_valid;
  assign MMIOTileLinkManager_1_io_inner_release_bits_addr_beat = PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_inner_release_bits_addr_block = PortedTileLinkCrossbar_1_io_managers_1_release_bits_addr_block;
  assign MMIOTileLinkManager_1_io_inner_release_bits_client_xact_id = PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_xact_id;
  assign MMIOTileLinkManager_1_io_inner_release_bits_voluntary = PortedTileLinkCrossbar_1_io_managers_1_release_bits_voluntary;
  assign MMIOTileLinkManager_1_io_inner_release_bits_r_type = PortedTileLinkCrossbar_1_io_managers_1_release_bits_r_type;
  assign MMIOTileLinkManager_1_io_inner_release_bits_data = PortedTileLinkCrossbar_1_io_managers_1_release_bits_data;
  assign MMIOTileLinkManager_1_io_inner_release_bits_client_id = PortedTileLinkCrossbar_1_io_managers_1_release_bits_client_id;
  assign MMIOTileLinkManager_1_io_incoherent_0 = GEN_0;
  assign MMIOTileLinkManager_1_io_outer_acquire_ready = ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign MMIOTileLinkManager_1_io_outer_grant_valid = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_valid;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_addr_beat = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_client_xact_id = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_manager_xact_id = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id[0];
  assign MMIOTileLinkManager_1_io_outer_grant_bits_is_builtin_type = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_g_type = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign MMIOTileLinkManager_1_io_outer_grant_bits_data = ClientUncachedTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign TileLinkMemoryInterconnect_1_clk = clk;
  assign TileLinkMemoryInterconnect_1_reset = reset;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_valid = ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_a_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_union = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  assign TileLinkMemoryInterconnect_1_io_in_0_acquire_bits_data = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  assign TileLinkMemoryInterconnect_1_io_in_0_grant_ready = ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  assign TileLinkMemoryInterconnect_1_io_out_0_acquire_ready = io_mem_0_acquire_ready;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_valid = io_mem_0_grant_valid;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_addr_beat = io_mem_0_grant_bits_addr_beat;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_client_xact_id = io_mem_0_grant_bits_client_xact_id;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_manager_xact_id = io_mem_0_grant_bits_manager_xact_id;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_is_builtin_type = io_mem_0_grant_bits_is_builtin_type;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_g_type = io_mem_0_grant_bits_g_type;
  assign TileLinkMemoryInterconnect_1_io_out_0_grant_bits_data = io_mem_0_grant_bits_data;
  assign ClientTileLinkIOUnwrapper_1_clk = clk;
  assign ClientTileLinkIOUnwrapper_1_reset = reset;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_valid = ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_probe_ready = ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_valid = ClientTileLinkEnqueuer_1_io_outer_release_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary = ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type = ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_data = ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_grant_ready = ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_valid = ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_acquire_ready = TileLinkMemoryInterconnect_1_io_in_0_acquire_ready;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_valid = TileLinkMemoryInterconnect_1_io_in_0_grant_valid;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_g_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data = TileLinkMemoryInterconnect_1_io_in_0_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_clk = clk;
  assign ClientTileLinkEnqueuer_1_reset = reset;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_valid = L2BroadcastHub_1_io_outer_acquire_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = L2BroadcastHub_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = L2BroadcastHub_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = L2BroadcastHub_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = L2BroadcastHub_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = L2BroadcastHub_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union = L2BroadcastHub_1_io_outer_acquire_bits_union;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data = L2BroadcastHub_1_io_outer_acquire_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_probe_ready = L2BroadcastHub_1_io_outer_probe_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_release_valid = L2BroadcastHub_1_io_outer_release_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat = L2BroadcastHub_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block = L2BroadcastHub_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id = L2BroadcastHub_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary = L2BroadcastHub_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type = L2BroadcastHub_1_io_outer_release_bits_r_type;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_data = L2BroadcastHub_1_io_outer_release_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_grant_ready = L2BroadcastHub_1_io_outer_grant_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_valid = L2BroadcastHub_1_io_outer_finish_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id = L2BroadcastHub_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id = L2BroadcastHub_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_acquire_ready = ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_valid = ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  assign ClientTileLinkEnqueuer_1_io_outer_release_ready = ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_valid = ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_data = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_finish_ready = ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  assign ClientUncachedTileLinkEnqueuer_1_clk = clk;
  assign ClientUncachedTileLinkEnqueuer_1_reset = reset;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_valid = MMIOTileLinkManager_1_io_outer_acquire_valid;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = MMIOTileLinkManager_1_io_outer_acquire_bits_addr_block;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = MMIOTileLinkManager_1_io_outer_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = MMIOTileLinkManager_1_io_outer_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = MMIOTileLinkManager_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = MMIOTileLinkManager_1_io_outer_acquire_bits_a_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_union = MMIOTileLinkManager_1_io_outer_acquire_bits_union;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_acquire_bits_data = MMIOTileLinkManager_1_io_outer_acquire_bits_data;
  assign ClientUncachedTileLinkEnqueuer_1_io_inner_grant_ready = MMIOTileLinkManager_1_io_outer_grant_ready;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_ready = TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_valid = TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = {{2'd0}, TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id};
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_g_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  assign ClientUncachedTileLinkEnqueuer_1_io_outer_grant_bits_data = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_clk = clk;
  assign TileLinkRecursiveInterconnect_2_reset = reset;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data = ClientUncachedTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_in_0_grant_ready = ClientUncachedTileLinkEnqueuer_1_io_outer_grant_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready = DebugModule_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_valid = DebugModule_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat = DebugModule_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id = DebugModule_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id = DebugModule_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type = DebugModule_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type = DebugModule_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data = DebugModule_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready = ROMSlave_1_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_valid = ROMSlave_1_io_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat = ROMSlave_1_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id = ROMSlave_1_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id = ROMSlave_1_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type = ROMSlave_1_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type = ROMSlave_1_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data = ROMSlave_1_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready = PLIC_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_valid = PLIC_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat = PLIC_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id = PLIC_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id = PLIC_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type = PLIC_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type = PLIC_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data = PLIC_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready = PRCI_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_valid = PRCI_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat = PRCI_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id = PRCI_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id = PRCI_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type = PRCI_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type = PRCI_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data = PRCI_1_io_tl_grant_bits_data;
  assign PLIC_1_clk = clk;
  assign PLIC_1_reset = reset;
  assign PLIC_1_io_devices_0_valid = LevelGateway_2_io_plic_valid;
  assign PLIC_1_io_devices_1_valid = LevelGateway_1_1_io_plic_valid;
  assign PLIC_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  assign PLIC_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  assign PLIC_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  assign PLIC_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  assign PLIC_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  assign PLIC_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  assign PLIC_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  assign PLIC_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  assign PLIC_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  assign LevelGateway_2_clk = clk;
  assign LevelGateway_2_reset = reset;
  assign LevelGateway_2_io_interrupt = io_interrupts_0;
  assign LevelGateway_2_io_plic_ready = PLIC_1_io_devices_0_ready;
  assign LevelGateway_2_io_plic_complete = PLIC_1_io_devices_0_complete;
  assign LevelGateway_1_1_clk = clk;
  assign LevelGateway_1_1_reset = reset;
  assign LevelGateway_1_1_io_interrupt = io_interrupts_1;
  assign LevelGateway_1_1_io_plic_ready = PLIC_1_io_devices_1_ready;
  assign LevelGateway_1_1_io_plic_complete = PLIC_1_io_devices_1_complete;
  assign DebugModule_1_clk = clk;
  assign DebugModule_1_reset = reset;
  assign DebugModule_1_io_db_req_valid = io_debug_req_valid;
  assign DebugModule_1_io_db_req_bits_addr = io_debug_req_bits_addr;
  assign DebugModule_1_io_db_req_bits_data = io_debug_req_bits_data;
  assign DebugModule_1_io_db_req_bits_op = io_debug_req_bits_op;
  assign DebugModule_1_io_db_resp_ready = io_debug_resp_ready;
  assign DebugModule_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  assign DebugModule_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  assign DebugModule_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  assign DebugModule_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  assign DebugModule_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  assign DebugModule_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  assign DebugModule_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  assign DebugModule_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  assign DebugModule_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  assign PRCI_1_clk = clk;
  assign PRCI_1_reset = reset;
  assign PRCI_1_io_interrupts_0_meip = PLIC_1_io_harts_0;
  assign PRCI_1_io_interrupts_0_seip = PLIC_1_io_harts_1;
  assign PRCI_1_io_interrupts_0_debug = DebugModule_1_io_debugInterrupts_0;
  assign PRCI_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  assign PRCI_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  assign PRCI_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  assign PRCI_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  assign PRCI_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  assign PRCI_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  assign PRCI_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  assign PRCI_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  assign PRCI_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  assign PRCI_1_io_rtcTick = io_rtcTick;
  assign ROMSlave_1_clk = clk;
  assign ROMSlave_1_reset = reset;
  assign ROMSlave_1_io_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  assign ROMSlave_1_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  assign ROMSlave_1_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  assign ROMSlave_1_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  assign ROMSlave_1_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  assign ROMSlave_1_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  assign ROMSlave_1_io_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  assign ROMSlave_1_io_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  assign ROMSlave_1_io_grant_ready = TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_0 = GEN_1[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_1 = {1{$random}};
  end
`endif
endmodule
module ReorderQueue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [2:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [2:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] T_229_addr_beat [0:7];
  reg [31:0] GEN_26;
  wire [2:0] T_229_addr_beat_T_249_data;
  wire [2:0] T_229_addr_beat_T_249_addr;
  wire  T_229_addr_beat_T_249_en;
  wire [2:0] T_229_addr_beat_T_275_data;
  wire [2:0] T_229_addr_beat_T_275_addr;
  wire  T_229_addr_beat_T_275_mask;
  wire  T_229_addr_beat_T_275_en;
  reg  T_229_subblock [0:7];
  reg [31:0] GEN_27;
  wire  T_229_subblock_T_249_data;
  wire [2:0] T_229_subblock_T_249_addr;
  wire  T_229_subblock_T_249_en;
  wire  T_229_subblock_T_275_data;
  wire [2:0] T_229_subblock_T_275_addr;
  wire  T_229_subblock_T_275_mask;
  wire  T_229_subblock_T_275_en;
  wire  T_243_0;
  wire  T_243_1;
  wire  T_243_2;
  wire  T_243_3;
  wire  T_243_4;
  wire  T_243_5;
  wire  T_243_6;
  wire  T_243_7;
  reg  T_247_0;
  reg [31:0] GEN_28;
  reg  T_247_1;
  reg [31:0] GEN_29;
  reg  T_247_2;
  reg [31:0] GEN_30;
  reg  T_247_3;
  reg [31:0] GEN_31;
  reg  T_247_4;
  reg [31:0] GEN_32;
  reg  T_247_5;
  reg [31:0] GEN_33;
  reg  T_247_6;
  reg [31:0] GEN_50;
  reg  T_247_7;
  reg [31:0] GEN_59;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_1;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  T_273;
  wire  T_274;
  wire  GEN_2;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_3;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  assign io_enq_ready = GEN_0;
  assign io_deq_data_addr_beat = T_229_addr_beat_T_249_data;
  assign io_deq_data_subblock = T_229_subblock_T_249_data;
  assign io_deq_matches = T_273;
  assign T_229_addr_beat_T_249_addr = io_deq_tag;
  assign T_229_addr_beat_T_249_en = 1'h1;
  assign T_229_addr_beat_T_249_data = T_229_addr_beat[T_229_addr_beat_T_249_addr];
  assign T_229_addr_beat_T_275_data = io_enq_bits_data_addr_beat;
  assign T_229_addr_beat_T_275_addr = io_enq_bits_tag;
  assign T_229_addr_beat_T_275_mask = T_274;
  assign T_229_addr_beat_T_275_en = T_274;
  assign T_229_subblock_T_249_addr = io_deq_tag;
  assign T_229_subblock_T_249_en = 1'h1;
  assign T_229_subblock_T_249_data = T_229_subblock[T_229_subblock_T_249_addr];
  assign T_229_subblock_T_275_data = io_enq_bits_data_subblock;
  assign T_229_subblock_T_275_addr = io_enq_bits_tag;
  assign T_229_subblock_T_275_mask = T_274;
  assign T_229_subblock_T_275_en = T_274;
  assign T_243_0 = 1'h1;
  assign T_243_1 = 1'h1;
  assign T_243_2 = 1'h1;
  assign T_243_3 = 1'h1;
  assign T_243_4 = 1'h1;
  assign T_243_5 = 1'h1;
  assign T_243_6 = 1'h1;
  assign T_243_7 = 1'h1;
  assign GEN_0 = GEN_10;
  assign GEN_4 = 3'h1 == io_enq_bits_tag ? T_247_1 : T_247_0;
  assign GEN_5 = 3'h2 == io_enq_bits_tag ? T_247_2 : GEN_4;
  assign GEN_6 = 3'h3 == io_enq_bits_tag ? T_247_3 : GEN_5;
  assign GEN_7 = 3'h4 == io_enq_bits_tag ? T_247_4 : GEN_6;
  assign GEN_8 = 3'h5 == io_enq_bits_tag ? T_247_5 : GEN_7;
  assign GEN_9 = 3'h6 == io_enq_bits_tag ? T_247_6 : GEN_8;
  assign GEN_10 = 3'h7 == io_enq_bits_tag ? T_247_7 : GEN_9;
  assign GEN_1 = GEN_17;
  assign GEN_11 = 3'h1 == io_deq_tag ? T_247_1 : T_247_0;
  assign GEN_12 = 3'h2 == io_deq_tag ? T_247_2 : GEN_11;
  assign GEN_13 = 3'h3 == io_deq_tag ? T_247_3 : GEN_12;
  assign GEN_14 = 3'h4 == io_deq_tag ? T_247_4 : GEN_13;
  assign GEN_15 = 3'h5 == io_deq_tag ? T_247_5 : GEN_14;
  assign GEN_16 = 3'h6 == io_deq_tag ? T_247_6 : GEN_15;
  assign GEN_17 = 3'h7 == io_deq_tag ? T_247_7 : GEN_16;
  assign T_273 = GEN_1 == 1'h0;
  assign T_274 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_18 = 3'h0 == io_enq_bits_tag ? GEN_2 : T_247_0;
  assign GEN_19 = 3'h1 == io_enq_bits_tag ? GEN_2 : T_247_1;
  assign GEN_20 = 3'h2 == io_enq_bits_tag ? GEN_2 : T_247_2;
  assign GEN_21 = 3'h3 == io_enq_bits_tag ? GEN_2 : T_247_3;
  assign GEN_22 = 3'h4 == io_enq_bits_tag ? GEN_2 : T_247_4;
  assign GEN_23 = 3'h5 == io_enq_bits_tag ? GEN_2 : T_247_5;
  assign GEN_24 = 3'h6 == io_enq_bits_tag ? GEN_2 : T_247_6;
  assign GEN_25 = 3'h7 == io_enq_bits_tag ? GEN_2 : T_247_7;
  assign GEN_34 = T_274 ? GEN_18 : T_247_0;
  assign GEN_35 = T_274 ? GEN_19 : T_247_1;
  assign GEN_36 = T_274 ? GEN_20 : T_247_2;
  assign GEN_37 = T_274 ? GEN_21 : T_247_3;
  assign GEN_38 = T_274 ? GEN_22 : T_247_4;
  assign GEN_39 = T_274 ? GEN_23 : T_247_5;
  assign GEN_40 = T_274 ? GEN_24 : T_247_6;
  assign GEN_41 = T_274 ? GEN_25 : T_247_7;
  assign GEN_3 = 1'h1;
  assign GEN_42 = 3'h0 == io_deq_tag ? GEN_3 : GEN_34;
  assign GEN_43 = 3'h1 == io_deq_tag ? GEN_3 : GEN_35;
  assign GEN_44 = 3'h2 == io_deq_tag ? GEN_3 : GEN_36;
  assign GEN_45 = 3'h3 == io_deq_tag ? GEN_3 : GEN_37;
  assign GEN_46 = 3'h4 == io_deq_tag ? GEN_3 : GEN_38;
  assign GEN_47 = 3'h5 == io_deq_tag ? GEN_3 : GEN_39;
  assign GEN_48 = 3'h6 == io_deq_tag ? GEN_3 : GEN_40;
  assign GEN_49 = 3'h7 == io_deq_tag ? GEN_3 : GEN_41;
  assign GEN_51 = io_deq_valid ? GEN_42 : GEN_34;
  assign GEN_52 = io_deq_valid ? GEN_43 : GEN_35;
  assign GEN_53 = io_deq_valid ? GEN_44 : GEN_36;
  assign GEN_54 = io_deq_valid ? GEN_45 : GEN_37;
  assign GEN_55 = io_deq_valid ? GEN_46 : GEN_38;
  assign GEN_56 = io_deq_valid ? GEN_47 : GEN_39;
  assign GEN_57 = io_deq_valid ? GEN_48 : GEN_40;
  assign GEN_58 = io_deq_valid ? GEN_49 : GEN_41;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_26 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    T_229_addr_beat[initvar] = GEN_26[2:0];
  `endif
  GEN_27 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    T_229_subblock[initvar] = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_28 = {1{$random}};
  T_247_0 = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_29 = {1{$random}};
  T_247_1 = GEN_29[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_30 = {1{$random}};
  T_247_2 = GEN_30[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_31 = {1{$random}};
  T_247_3 = GEN_31[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_32 = {1{$random}};
  T_247_4 = GEN_32[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_33 = {1{$random}};
  T_247_5 = GEN_33[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_50 = {1{$random}};
  T_247_6 = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_59 = {1{$random}};
  T_247_7 = GEN_59[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_229_addr_beat_T_275_en & T_229_addr_beat_T_275_mask) begin
      T_229_addr_beat[T_229_addr_beat_T_275_addr] <= T_229_addr_beat_T_275_data;
    end
    if(T_229_subblock_T_275_en & T_229_subblock_T_275_mask) begin
      T_229_subblock[T_229_subblock_T_275_addr] <= T_229_subblock_T_275_data;
    end
    if(reset) begin
      T_247_0 <= T_243_0;
    end else begin
      if(io_deq_valid) begin
        if(3'h0 == io_deq_tag) begin
          T_247_0 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h0 == io_enq_bits_tag) begin
              T_247_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h0 == io_enq_bits_tag) begin
            T_247_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_1 <= T_243_1;
    end else begin
      if(io_deq_valid) begin
        if(3'h1 == io_deq_tag) begin
          T_247_1 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h1 == io_enq_bits_tag) begin
              T_247_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h1 == io_enq_bits_tag) begin
            T_247_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_2 <= T_243_2;
    end else begin
      if(io_deq_valid) begin
        if(3'h2 == io_deq_tag) begin
          T_247_2 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h2 == io_enq_bits_tag) begin
              T_247_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h2 == io_enq_bits_tag) begin
            T_247_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_3 <= T_243_3;
    end else begin
      if(io_deq_valid) begin
        if(3'h3 == io_deq_tag) begin
          T_247_3 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h3 == io_enq_bits_tag) begin
              T_247_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h3 == io_enq_bits_tag) begin
            T_247_3 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_4 <= T_243_4;
    end else begin
      if(io_deq_valid) begin
        if(3'h4 == io_deq_tag) begin
          T_247_4 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h4 == io_enq_bits_tag) begin
              T_247_4 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h4 == io_enq_bits_tag) begin
            T_247_4 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_5 <= T_243_5;
    end else begin
      if(io_deq_valid) begin
        if(3'h5 == io_deq_tag) begin
          T_247_5 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h5 == io_enq_bits_tag) begin
              T_247_5 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h5 == io_enq_bits_tag) begin
            T_247_5 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_6 <= T_243_6;
    end else begin
      if(io_deq_valid) begin
        if(3'h6 == io_deq_tag) begin
          T_247_6 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h6 == io_enq_bits_tag) begin
              T_247_6 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h6 == io_enq_bits_tag) begin
            T_247_6 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_247_7 <= T_243_7;
    end else begin
      if(io_deq_valid) begin
        if(3'h7 == io_deq_tag) begin
          T_247_7 <= GEN_3;
        end else begin
          if(T_274) begin
            if(3'h7 == io_enq_bits_tag) begin
              T_247_7 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_274) begin
          if(3'h7 == io_enq_bits_tag) begin
            T_247_7 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module IdMapper(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [2:0] io_req_in_id,
  output [4:0] io_req_out_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_out_id,
  output [2:0] io_resp_in_id
);
  assign io_req_ready = 1'h1;
  assign io_req_out_id = {{2'd0}, io_req_in_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_in_id = io_resp_out_id[2:0];
endmodule
module LockingArbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [2:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [2:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [2:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0_ready;
  wire  GEN_0_valid;
  wire [2:0] GEN_0_bits_addr_beat;
  wire [2:0] GEN_0_bits_client_xact_id;
  wire  GEN_0_bits_manager_xact_id;
  wire  GEN_0_bits_is_builtin_type;
  wire [3:0] GEN_0_bits_g_type;
  wire [63:0] GEN_0_bits_data;
  wire  GEN_0_bits_client_id;
  wire  GEN_8;
  wire  GEN_9;
  wire [2:0] GEN_10;
  wire [2:0] GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire [3:0] GEN_14;
  wire [63:0] GEN_15;
  wire  GEN_16;
  wire  GEN_1_ready;
  wire  GEN_1_valid;
  wire [2:0] GEN_1_bits_addr_beat;
  wire [2:0] GEN_1_bits_client_xact_id;
  wire  GEN_1_bits_manager_xact_id;
  wire  GEN_1_bits_is_builtin_type;
  wire [3:0] GEN_1_bits_g_type;
  wire [63:0] GEN_1_bits_data;
  wire  GEN_1_bits_client_id;
  wire  GEN_2_ready;
  wire  GEN_2_valid;
  wire [2:0] GEN_2_bits_addr_beat;
  wire [2:0] GEN_2_bits_client_xact_id;
  wire  GEN_2_bits_manager_xact_id;
  wire  GEN_2_bits_is_builtin_type;
  wire [3:0] GEN_2_bits_g_type;
  wire [63:0] GEN_2_bits_data;
  wire  GEN_2_bits_client_id;
  wire  GEN_3_ready;
  wire  GEN_3_valid;
  wire [2:0] GEN_3_bits_addr_beat;
  wire [2:0] GEN_3_bits_client_xact_id;
  wire  GEN_3_bits_manager_xact_id;
  wire  GEN_3_bits_is_builtin_type;
  wire [3:0] GEN_3_bits_g_type;
  wire [63:0] GEN_3_bits_data;
  wire  GEN_3_bits_client_id;
  wire  GEN_4_ready;
  wire  GEN_4_valid;
  wire [2:0] GEN_4_bits_addr_beat;
  wire [2:0] GEN_4_bits_client_xact_id;
  wire  GEN_4_bits_manager_xact_id;
  wire  GEN_4_bits_is_builtin_type;
  wire [3:0] GEN_4_bits_g_type;
  wire [63:0] GEN_4_bits_data;
  wire  GEN_4_bits_client_id;
  wire  GEN_5_ready;
  wire  GEN_5_valid;
  wire [2:0] GEN_5_bits_addr_beat;
  wire [2:0] GEN_5_bits_client_xact_id;
  wire  GEN_5_bits_manager_xact_id;
  wire  GEN_5_bits_is_builtin_type;
  wire [3:0] GEN_5_bits_g_type;
  wire [63:0] GEN_5_bits_data;
  wire  GEN_5_bits_client_id;
  wire  GEN_6_ready;
  wire  GEN_6_valid;
  wire [2:0] GEN_6_bits_addr_beat;
  wire [2:0] GEN_6_bits_client_xact_id;
  wire  GEN_6_bits_manager_xact_id;
  wire  GEN_6_bits_is_builtin_type;
  wire [3:0] GEN_6_bits_g_type;
  wire [63:0] GEN_6_bits_data;
  wire  GEN_6_bits_client_id;
  wire  GEN_7_ready;
  wire  GEN_7_valid;
  wire [2:0] GEN_7_bits_addr_beat;
  wire [2:0] GEN_7_bits_client_xact_id;
  wire  GEN_7_bits_manager_xact_id;
  wire  GEN_7_bits_is_builtin_type;
  wire [3:0] GEN_7_bits_g_type;
  wire [63:0] GEN_7_bits_data;
  wire  GEN_7_bits_client_id;
  reg [2:0] T_766;
  reg [31:0] GEN_1;
  reg  T_768;
  reg [31:0] GEN_2;
  wire  T_770;
  wire [2:0] T_778_0;
  wire [3:0] GEN_0;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire  T_785;
  wire [3:0] T_789;
  wire [2:0] T_790;
  wire  GEN_80;
  wire [2:0] GEN_81;
  wire  GEN_82;
  wire  T_793;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire  T_800;
  wire  T_801;
  wire  GEN_83;
  assign io_in_0_ready = T_797;
  assign io_in_1_ready = T_801;
  assign io_out_valid = GEN_0_valid;
  assign io_out_bits_addr_beat = GEN_1_bits_addr_beat;
  assign io_out_bits_client_xact_id = GEN_2_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = GEN_3_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = GEN_4_bits_is_builtin_type;
  assign io_out_bits_g_type = GEN_5_bits_g_type;
  assign io_out_bits_data = GEN_6_bits_data;
  assign io_out_bits_client_id = GEN_7_bits_client_id;
  assign io_chosen = GEN_82;
  assign choice = GEN_83;
  assign GEN_0_ready = GEN_8;
  assign GEN_0_valid = GEN_9;
  assign GEN_0_bits_addr_beat = GEN_10;
  assign GEN_0_bits_client_xact_id = GEN_11;
  assign GEN_0_bits_manager_xact_id = GEN_12;
  assign GEN_0_bits_is_builtin_type = GEN_13;
  assign GEN_0_bits_g_type = GEN_14;
  assign GEN_0_bits_data = GEN_15;
  assign GEN_0_bits_client_id = GEN_16;
  assign GEN_8 = io_chosen ? io_in_1_ready : io_in_0_ready;
  assign GEN_9 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_11 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_12 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_13 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_14 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_15 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_16 = io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_1_ready = GEN_8;
  assign GEN_1_valid = GEN_9;
  assign GEN_1_bits_addr_beat = GEN_10;
  assign GEN_1_bits_client_xact_id = GEN_11;
  assign GEN_1_bits_manager_xact_id = GEN_12;
  assign GEN_1_bits_is_builtin_type = GEN_13;
  assign GEN_1_bits_g_type = GEN_14;
  assign GEN_1_bits_data = GEN_15;
  assign GEN_1_bits_client_id = GEN_16;
  assign GEN_2_ready = GEN_8;
  assign GEN_2_valid = GEN_9;
  assign GEN_2_bits_addr_beat = GEN_10;
  assign GEN_2_bits_client_xact_id = GEN_11;
  assign GEN_2_bits_manager_xact_id = GEN_12;
  assign GEN_2_bits_is_builtin_type = GEN_13;
  assign GEN_2_bits_g_type = GEN_14;
  assign GEN_2_bits_data = GEN_15;
  assign GEN_2_bits_client_id = GEN_16;
  assign GEN_3_ready = GEN_8;
  assign GEN_3_valid = GEN_9;
  assign GEN_3_bits_addr_beat = GEN_10;
  assign GEN_3_bits_client_xact_id = GEN_11;
  assign GEN_3_bits_manager_xact_id = GEN_12;
  assign GEN_3_bits_is_builtin_type = GEN_13;
  assign GEN_3_bits_g_type = GEN_14;
  assign GEN_3_bits_data = GEN_15;
  assign GEN_3_bits_client_id = GEN_16;
  assign GEN_4_ready = GEN_8;
  assign GEN_4_valid = GEN_9;
  assign GEN_4_bits_addr_beat = GEN_10;
  assign GEN_4_bits_client_xact_id = GEN_11;
  assign GEN_4_bits_manager_xact_id = GEN_12;
  assign GEN_4_bits_is_builtin_type = GEN_13;
  assign GEN_4_bits_g_type = GEN_14;
  assign GEN_4_bits_data = GEN_15;
  assign GEN_4_bits_client_id = GEN_16;
  assign GEN_5_ready = GEN_8;
  assign GEN_5_valid = GEN_9;
  assign GEN_5_bits_addr_beat = GEN_10;
  assign GEN_5_bits_client_xact_id = GEN_11;
  assign GEN_5_bits_manager_xact_id = GEN_12;
  assign GEN_5_bits_is_builtin_type = GEN_13;
  assign GEN_5_bits_g_type = GEN_14;
  assign GEN_5_bits_data = GEN_15;
  assign GEN_5_bits_client_id = GEN_16;
  assign GEN_6_ready = GEN_8;
  assign GEN_6_valid = GEN_9;
  assign GEN_6_bits_addr_beat = GEN_10;
  assign GEN_6_bits_client_xact_id = GEN_11;
  assign GEN_6_bits_manager_xact_id = GEN_12;
  assign GEN_6_bits_is_builtin_type = GEN_13;
  assign GEN_6_bits_g_type = GEN_14;
  assign GEN_6_bits_data = GEN_15;
  assign GEN_6_bits_client_id = GEN_16;
  assign GEN_7_ready = GEN_8;
  assign GEN_7_valid = GEN_9;
  assign GEN_7_bits_addr_beat = GEN_10;
  assign GEN_7_bits_client_xact_id = GEN_11;
  assign GEN_7_bits_manager_xact_id = GEN_12;
  assign GEN_7_bits_is_builtin_type = GEN_13;
  assign GEN_7_bits_g_type = GEN_14;
  assign GEN_7_bits_data = GEN_15;
  assign GEN_7_bits_client_id = GEN_16;
  assign T_770 = T_766 != 3'h0;
  assign T_778_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_778_0};
  assign T_780 = io_out_bits_g_type == GEN_0;
  assign T_781 = io_out_bits_g_type == 4'h0;
  assign T_782 = io_out_bits_is_builtin_type ? T_780 : T_781;
  assign T_784 = io_out_ready & io_out_valid;
  assign T_785 = T_784 & T_782;
  assign T_789 = T_766 + 3'h1;
  assign T_790 = T_789[2:0];
  assign GEN_80 = T_785 ? io_chosen : T_768;
  assign GEN_81 = T_785 ? T_790 : T_766;
  assign GEN_82 = T_770 ? T_768 : choice;
  assign T_793 = io_in_0_valid == 1'h0;
  assign T_795 = T_768 == 1'h0;
  assign T_796 = T_770 ? T_795 : 1'h1;
  assign T_797 = T_796 & io_out_ready;
  assign T_800 = T_770 ? T_768 : T_793;
  assign T_801 = T_800 & io_out_ready;
  assign GEN_83 = io_in_0_valid ? 1'h0 : 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_766 = GEN_1[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_2 = {1{$random}};
  T_768 = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_785) begin
        T_766 <= T_790;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_785) begin
        T_768 <= io_chosen;
      end
    end
  end
endmodule
module NastiIOTileLinkIOConverter(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [2:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [10:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [2:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_688_0;
  wire [2:0] T_688_1;
  wire [2:0] T_688_2;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire  T_694;
  wire  has_data;
  wire [2:0] T_703_0;
  wire [2:0] T_703_1;
  wire [2:0] T_703_2;
  wire  T_705;
  wire  T_706;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  is_subblock;
  wire [2:0] T_718_0;
  wire  T_720;
  wire  is_multibeat;
  wire  T_721;
  wire  T_722;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_11;
  wire  T_725;
  wire [3:0] T_727;
  wire [2:0] T_728;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_730;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [2:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [2:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [2:0] get_id_mapper_io_req_in_id;
  wire [4:0] get_id_mapper_io_req_out_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_out_id;
  wire [2:0] get_id_mapper_io_resp_in_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [2:0] put_id_mapper_io_req_in_id;
  wire [4:0] put_id_mapper_io_req_out_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_out_id;
  wire [2:0] put_id_mapper_io_resp_in_id;
  wire  T_755;
  wire  put_id_mask;
  wire  T_757;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_12;
  reg [4:0] w_id_reg;
  reg [31:0] GEN_13;
  wire [4:0] w_id;
  wire  aw_ready;
  wire  T_760;
  wire  T_762;
  wire  T_763;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_14;
  wire  T_766;
  wire [3:0] T_768;
  wire [2:0] T_769;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_770;
  wire  T_771;
  wire  T_773;
  wire  T_774;
  wire  T_775;
  wire  T_776;
  wire  T_778;
  wire  T_779;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire [2:0] T_792_0;
  wire [2:0] T_792_1;
  wire  T_794;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire [2:0] T_798;
  wire [2:0] T_800;
  wire [28:0] T_801;
  wire [31:0] T_802;
  wire [1:0] T_803;
  wire [1:0] T_805;
  wire [2:0] T_808;
  wire [31:0] T_821_addr;
  wire [7:0] T_821_len;
  wire [2:0] T_821_size;
  wire [1:0] T_821_burst;
  wire  T_821_lock;
  wire [3:0] T_821_cache;
  wire [2:0] T_821_prot;
  wire [3:0] T_821_qos;
  wire [3:0] T_821_region;
  wire [4:0] T_821_id;
  wire  T_821_user;
  wire  T_840;
  wire  T_841;
  wire  T_865;
  wire  T_866;
  wire  T_868;
  wire  T_869;
  wire  T_870;
  wire [7:0] T_871;
  wire [7:0] T_873;
  wire [7:0] T_874;
  wire [7:0] T_875;
  wire  all_inside_0_0;
  wire  all_inside_0_1;
  wire  all_inside_0_2;
  wire  all_inside_0_3;
  wire  all_inside_0_4;
  wire  all_inside_0_5;
  wire  all_inside_0_6;
  wire  all_inside_0_7;
  wire  T_876;
  wire  T_877;
  wire  T_878;
  wire  T_879;
  wire  T_880;
  wire  T_881;
  wire  T_888;
  wire [1:0] T_889;
  wire [1:0] T_891;
  wire  T_892;
  wire  T_893;
  wire  T_894;
  wire  T_895;
  wire  T_896;
  wire  T_897;
  wire  T_898;
  wire  T_899;
  wire [2:0] T_900;
  wire [1:0] T_902;
  wire  T_903;
  wire  T_904;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_908;
  wire  T_909;
  wire  T_910;
  wire  T_911;
  wire  T_912;
  wire  T_913;
  wire  T_914;
  wire  T_915;
  wire  T_916;
  wire  T_917;
  wire  T_918;
  wire  T_919;
  wire  T_920;
  wire [3:0] put_offset;
  wire [1:0] put_size;
  wire  T_923;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire [2:0] T_934_0;
  wire [2:0] T_934_1;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire [2:0] T_942;
  wire [31:0] T_944;
  wire [3:0] T_946;
  wire [31:0] GEN_7;
  wire [31:0] T_947;
  wire [1:0] T_949;
  wire [2:0] T_952;
  wire [31:0] T_965_addr;
  wire [7:0] T_965_len;
  wire [2:0] T_965_size;
  wire [1:0] T_965_burst;
  wire  T_965_lock;
  wire [3:0] T_965_cache;
  wire [2:0] T_965_prot;
  wire [3:0] T_965_qos;
  wire [3:0] T_965_region;
  wire [4:0] T_965_id;
  wire  T_965_user;
  wire  T_984;
  wire  T_1024;
  wire  T_1025;
  wire [63:0] T_1032_data;
  wire  T_1032_last;
  wire [4:0] T_1032_id;
  wire [7:0] T_1032_strb;
  wire  T_1032_user;
  wire  T_1039;
  wire  T_1040;
  wire  T_1041;
  wire  T_1042;
  wire  T_1043;
  wire  T_1047;
  wire  T_1048;
  wire  GEN_2;
  wire [4:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_1051;
  wire [2:0] T_1059_0;
  wire [3:0] GEN_8;
  wire  T_1061;
  wire  T_1062;
  wire  T_1063;
  wire  T_1065;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_15;
  wire [3:0] T_1070;
  wire [2:0] T_1071;
  wire [2:0] GEN_6;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [2:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1133_addr_beat;
  wire [2:0] T_1133_client_xact_id;
  wire  T_1133_manager_xact_id;
  wire  T_1133_is_builtin_type;
  wire [3:0] T_1133_g_type;
  wire [63:0] T_1133_data;
  wire  T_1161;
  wire  T_1162;
  wire  T_1163;
  wire  T_1165;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1171;
  wire [2:0] T_1204_addr_beat;
  wire [2:0] T_1204_client_xact_id;
  wire  T_1204_manager_xact_id;
  wire  T_1204_is_builtin_type;
  wire [3:0] T_1204_g_type;
  wire [63:0] T_1204_data;
  wire  T_1232;
  wire  T_1233;
  wire  T_1234;
  wire  T_1236;
  wire  T_1238;
  wire  T_1240;
  wire  T_1241;
  wire  T_1242;
  wire  T_1244;
  wire  T_1246;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1252;
  wire  GEN_9;
  reg [31:0] GEN_16;
  wire  GEN_10;
  reg [31:0] GEN_17;
  ReorderQueue_2 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  IdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_in_id(get_id_mapper_io_req_in_id),
    .io_req_out_id(get_id_mapper_io_req_out_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_out_id(get_id_mapper_io_resp_out_id),
    .io_resp_in_id(get_id_mapper_io_resp_in_id)
  );
  IdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_in_id(put_id_mapper_io_req_in_id),
    .io_req_out_id(put_id_mapper_io_req_out_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_out_id(put_id_mapper_io_resp_out_id),
    .io_resp_in_id(put_id_mapper_io_resp_in_id)
  );
  LockingArbiter_2 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_1043;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_926;
  assign io_nasti_aw_bits_addr = T_965_addr;
  assign io_nasti_aw_bits_len = T_965_len;
  assign io_nasti_aw_bits_size = T_965_size;
  assign io_nasti_aw_bits_burst = T_965_burst;
  assign io_nasti_aw_bits_lock = T_965_lock;
  assign io_nasti_aw_bits_cache = T_965_cache;
  assign io_nasti_aw_bits_prot = T_965_prot;
  assign io_nasti_aw_bits_qos = T_965_qos;
  assign io_nasti_aw_bits_region = T_965_region;
  assign io_nasti_aw_bits_id = T_965_id;
  assign io_nasti_aw_bits_user = T_965_user;
  assign io_nasti_w_valid = T_984;
  assign io_nasti_w_bits_data = T_1032_data;
  assign io_nasti_w_bits_last = T_1032_last;
  assign io_nasti_w_bits_id = T_1032_id;
  assign io_nasti_w_bits_strb = T_1032_strb;
  assign io_nasti_w_bits_user = T_1032_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_784;
  assign io_nasti_ar_bits_addr = T_821_addr;
  assign io_nasti_ar_bits_len = T_821_len;
  assign io_nasti_ar_bits_size = T_821_size;
  assign io_nasti_ar_bits_burst = T_821_burst;
  assign io_nasti_ar_bits_lock = T_821_lock;
  assign io_nasti_ar_bits_cache = T_821_cache;
  assign io_nasti_ar_bits_prot = T_821_prot;
  assign io_nasti_ar_bits_qos = T_821_qos;
  assign io_nasti_ar_bits_region = T_821_region;
  assign io_nasti_ar_bits_id = T_821_id;
  assign io_nasti_ar_bits_user = T_821_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_688_0 = 3'h2;
  assign T_688_1 = 3'h3;
  assign T_688_2 = 3'h4;
  assign T_690 = io_tl_acquire_bits_a_type == T_688_0;
  assign T_691 = io_tl_acquire_bits_a_type == T_688_1;
  assign T_692 = io_tl_acquire_bits_a_type == T_688_2;
  assign T_693 = T_690 | T_691;
  assign T_694 = T_693 | T_692;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_694;
  assign T_703_0 = 3'h2;
  assign T_703_1 = 3'h0;
  assign T_703_2 = 3'h4;
  assign T_705 = io_tl_acquire_bits_a_type == T_703_0;
  assign T_706 = io_tl_acquire_bits_a_type == T_703_1;
  assign T_707 = io_tl_acquire_bits_a_type == T_703_2;
  assign T_708 = T_705 | T_706;
  assign T_709 = T_708 | T_707;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_709;
  assign T_718_0 = 3'h3;
  assign T_720 = io_tl_acquire_bits_a_type == T_718_0;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_720;
  assign T_721 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_722 = T_721 & is_multibeat;
  assign T_725 = tl_cnt_out == 3'h7;
  assign T_727 = tl_cnt_out + 3'h1;
  assign T_728 = T_727[2:0];
  assign GEN_0 = T_722 ? T_728 : tl_cnt_out;
  assign tl_wrap_out = T_722 & T_725;
  assign T_730 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_730;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_771;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id[2:0];
  assign roq_io_deq_valid = T_774;
  assign roq_io_deq_tag = io_nasti_r_bits_id[2:0];
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_776;
  assign get_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_778;
  assign get_id_mapper_io_resp_out_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_781;
  assign put_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_782;
  assign put_id_mapper_io_resp_out_id = io_nasti_b_bits_id;
  assign T_755 = io_tl_acquire_bits_addr_beat == 3'h0;
  assign put_id_mask = is_subblock | T_755;
  assign T_757 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_757;
  assign w_id = w_inflight ? w_id_reg : put_id_mapper_io_req_out_id;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_760 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_762 = roq_io_deq_data_subblock == 1'h0;
  assign T_763 = T_760 & T_762;
  assign T_766 = nasti_cnt_out == 3'h7;
  assign T_768 = nasti_cnt_out + 3'h1;
  assign T_769 = T_768[2:0];
  assign GEN_1 = T_763 ? T_769 : nasti_cnt_out;
  assign nasti_wrap_out = T_763 & T_766;
  assign T_770 = get_valid & io_nasti_ar_ready;
  assign T_771 = T_770 & get_id_mapper_io_req_ready;
  assign T_773 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_774 = T_760 & T_773;
  assign T_775 = get_valid & roq_io_enq_ready;
  assign T_776 = T_775 & io_nasti_ar_ready;
  assign T_778 = T_760 & io_nasti_r_bits_last;
  assign T_779 = put_valid & aw_ready;
  assign T_780 = T_779 & io_nasti_w_ready;
  assign T_781 = T_780 & put_id_mask;
  assign T_782 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_784 = T_775 & get_id_mapper_io_req_ready;
  assign T_792_0 = 3'h0;
  assign T_792_1 = 3'h4;
  assign T_794 = io_tl_acquire_bits_a_type == T_792_0;
  assign T_795 = io_tl_acquire_bits_a_type == T_792_1;
  assign T_796 = T_794 | T_795;
  assign T_797 = io_tl_acquire_bits_is_builtin_type & T_796;
  assign T_798 = io_tl_acquire_bits_union[10:8];
  assign T_800 = T_797 ? T_798 : 3'h0;
  assign T_801 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_802 = {T_801,T_800};
  assign T_803 = io_tl_acquire_bits_union[7:6];
  assign T_805 = is_subblock ? T_803 : 2'h3;
  assign T_808 = is_subblock ? 3'h0 : 3'h7;
  assign T_821_addr = T_802;
  assign T_821_len = {{5'd0}, T_808};
  assign T_821_size = {{1'd0}, T_805};
  assign T_821_burst = 2'h1;
  assign T_821_lock = 1'h0;
  assign T_821_cache = 4'h0;
  assign T_821_prot = 3'h0;
  assign T_821_qos = 4'h0;
  assign T_821_region = 4'h0;
  assign T_821_id = get_id_mapper_io_req_out_id;
  assign T_821_user = 1'h0;
  assign T_840 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_841 = io_tl_acquire_bits_is_builtin_type & T_840;
  assign T_865 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_866 = io_tl_acquire_bits_is_builtin_type & T_865;
  assign T_868 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_869 = io_tl_acquire_bits_is_builtin_type & T_868;
  assign T_870 = T_866 | T_869;
  assign T_871 = io_tl_acquire_bits_union[8:1];
  assign T_873 = T_870 ? T_871 : 8'h0;
  assign T_874 = T_841 ? 8'hff : T_873;
  assign T_875 = ~ T_874;
  assign all_inside_0_0 = T_875[0];
  assign all_inside_0_1 = T_875[1];
  assign all_inside_0_2 = T_875[2];
  assign all_inside_0_3 = T_875[3];
  assign all_inside_0_4 = T_875[4];
  assign all_inside_0_5 = T_875[5];
  assign all_inside_0_6 = T_875[6];
  assign all_inside_0_7 = T_875[7];
  assign T_876 = all_inside_0_0 & all_inside_0_1;
  assign T_877 = all_inside_0_2 & all_inside_0_3;
  assign T_878 = all_inside_0_4 & all_inside_0_5;
  assign T_879 = all_inside_0_6 & all_inside_0_7;
  assign T_880 = T_876 & T_877;
  assign T_881 = T_878 & T_879;
  assign T_888 = T_881 | T_880;
  assign T_889 = {1'h0,T_880};
  assign T_891 = T_888 ? 2'h2 : 2'h3;
  assign T_892 = T_881 & T_877;
  assign T_893 = T_881 & T_876;
  assign T_894 = T_880 & T_879;
  assign T_895 = T_880 & T_878;
  assign T_896 = T_893 | T_895;
  assign T_897 = T_892 | T_893;
  assign T_898 = T_897 | T_894;
  assign T_899 = T_898 | T_895;
  assign T_900 = {T_889,T_896};
  assign T_902 = T_899 ? 2'h1 : T_891;
  assign T_903 = T_892 & all_inside_0_1;
  assign T_904 = T_892 & all_inside_0_0;
  assign T_905 = T_893 & all_inside_0_3;
  assign T_906 = T_893 & all_inside_0_2;
  assign T_907 = T_894 & all_inside_0_5;
  assign T_908 = T_894 & all_inside_0_4;
  assign T_909 = T_895 & all_inside_0_7;
  assign T_910 = T_895 & all_inside_0_6;
  assign T_911 = T_904 | T_906;
  assign T_912 = T_911 | T_908;
  assign T_913 = T_912 | T_910;
  assign T_914 = T_903 | T_904;
  assign T_915 = T_914 | T_905;
  assign T_916 = T_915 | T_906;
  assign T_917 = T_916 | T_907;
  assign T_918 = T_917 | T_908;
  assign T_919 = T_918 | T_909;
  assign T_920 = T_919 | T_910;
  assign put_offset = {T_900,T_913};
  assign put_size = T_920 ? 2'h0 : T_902;
  assign T_923 = w_inflight == 1'h0;
  assign T_924 = put_valid & io_nasti_w_ready;
  assign T_925 = T_924 & put_id_ready;
  assign T_926 = T_925 & T_923;
  assign T_934_0 = 3'h0;
  assign T_934_1 = 3'h4;
  assign T_936 = io_tl_acquire_bits_a_type == T_934_0;
  assign T_937 = io_tl_acquire_bits_a_type == T_934_1;
  assign T_938 = T_936 | T_937;
  assign T_939 = io_tl_acquire_bits_is_builtin_type & T_938;
  assign T_942 = T_939 ? T_798 : 3'h0;
  assign T_944 = {T_801,T_942};
  assign T_946 = is_multibeat ? 4'h0 : put_offset;
  assign GEN_7 = {{28'd0}, T_946};
  assign T_947 = T_944 | GEN_7;
  assign T_949 = is_multibeat ? 2'h3 : put_size;
  assign T_952 = is_multibeat ? 3'h7 : 3'h0;
  assign T_965_addr = T_947;
  assign T_965_len = {{5'd0}, T_952};
  assign T_965_size = {{1'd0}, T_949};
  assign T_965_burst = 2'h1;
  assign T_965_lock = 1'h0;
  assign T_965_cache = 4'h0;
  assign T_965_prot = 3'h0;
  assign T_965_qos = 4'h0;
  assign T_965_region = 4'h0;
  assign T_965_id = put_id_mapper_io_req_out_id;
  assign T_965_user = 1'h0;
  assign T_984 = T_779 & put_id_ready;
  assign T_1024 = is_multibeat == 1'h0;
  assign T_1025 = w_inflight ? T_725 : T_1024;
  assign T_1032_data = io_tl_acquire_bits_data;
  assign T_1032_last = T_1025;
  assign T_1032_id = w_id;
  assign T_1032_strb = T_874;
  assign T_1032_user = 1'h0;
  assign T_1039 = aw_ready & io_nasti_w_ready;
  assign T_1040 = T_1039 & put_id_ready;
  assign T_1041 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_1042 = T_1041 & get_id_mapper_io_req_ready;
  assign T_1043 = has_data ? T_1040 : T_1042;
  assign T_1047 = T_923 & T_721;
  assign T_1048 = T_1047 & is_multibeat;
  assign GEN_2 = T_1048 ? 1'h1 : w_inflight;
  assign GEN_3 = T_1048 ? w_id : w_id_reg;
  assign GEN_4 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_5 = w_inflight ? GEN_4 : GEN_2;
  assign T_1051 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1059_0 = 3'h5;
  assign GEN_8 = {{1'd0}, T_1059_0};
  assign T_1061 = io_tl_grant_bits_g_type == GEN_8;
  assign T_1062 = io_tl_grant_bits_g_type == 4'h0;
  assign T_1063 = io_tl_grant_bits_is_builtin_type ? T_1061 : T_1062;
  assign T_1065 = T_1051 & T_1063;
  assign T_1070 = tl_cnt_in + 3'h1;
  assign T_1071 = T_1070[2:0];
  assign GEN_6 = T_1065 ? T_1071 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1133_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1133_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1133_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1133_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1133_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1133_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_9;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1204_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1204_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1204_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1204_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1204_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1204_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_10;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1103 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1105 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1133_addr_beat = T_1105;
  assign T_1133_client_xact_id = get_id_mapper_io_resp_in_id;
  assign T_1133_manager_xact_id = 1'h0;
  assign T_1133_is_builtin_type = 1'h1;
  assign T_1133_g_type = {{1'd0}, T_1103};
  assign T_1133_data = io_nasti_r_bits_data;
  assign T_1161 = roq_io_deq_valid == 1'h0;
  assign T_1162 = T_1161 | roq_io_deq_matches;
  assign T_1163 = T_1162 | reset;
  assign T_1165 = T_1163 == 1'h0;
  assign T_1167 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1168 = T_1167 | get_id_mapper_io_resp_matches;
  assign T_1169 = T_1168 | reset;
  assign T_1171 = T_1169 == 1'h0;
  assign T_1204_addr_beat = 3'h0;
  assign T_1204_client_xact_id = put_id_mapper_io_resp_in_id;
  assign T_1204_manager_xact_id = 1'h0;
  assign T_1204_is_builtin_type = 1'h1;
  assign T_1204_g_type = 4'h3;
  assign T_1204_data = 64'h0;
  assign T_1232 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1233 = T_1232 | put_id_mapper_io_resp_matches;
  assign T_1234 = T_1233 | reset;
  assign T_1236 = T_1234 == 1'h0;
  assign T_1238 = io_nasti_r_valid == 1'h0;
  assign T_1240 = io_nasti_r_bits_resp == 2'h0;
  assign T_1241 = T_1238 | T_1240;
  assign T_1242 = T_1241 | reset;
  assign T_1244 = T_1242 == 1'h0;
  assign T_1246 = io_nasti_b_valid == 1'h0;
  assign T_1248 = io_nasti_b_bits_resp == 2'h0;
  assign T_1249 = T_1246 | T_1248;
  assign T_1250 = T_1249 | reset;
  assign T_1252 = T_1250 == 1'h0;
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_9 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE_INVALID_ASSIGN
  assign GEN_10 = GEN_17[0:0];
  `endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  tl_cnt_out = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_12 = {1{$random}};
  w_inflight = GEN_12[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_13 = {1{$random}};
  w_id_reg = GEN_13[4:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_14 = {1{$random}};
  nasti_cnt_out = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_15 = {1{$random}};
  tl_cnt_in = GEN_15[2:0];
  `endif
  GEN_16 = {1{$random}};
  GEN_17 = {1{$random}};
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_722) begin
        tl_cnt_out <= T_728;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_1048) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_1048) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      w_id_reg <= 5'h0;
    end else begin
      if(T_1048) begin
        if(w_inflight) begin
        end else begin
          w_id_reg <= put_id_mapper_io_req_out_id;
        end
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_763) begin
        nasti_cnt_out <= T_769;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_1065) begin
        tl_cnt_in <= T_1071;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1165) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:220 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1171) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:222 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1236) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:234 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1244) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:236 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1252) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:237 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_19(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0] io_enq_bits_len,
  input  [2:0] io_enq_bits_size,
  input  [1:0] io_enq_bits_burst,
  input   io_enq_bits_lock,
  input  [3:0] io_enq_bits_cache,
  input  [2:0] io_enq_bits_prot,
  input  [3:0] io_enq_bits_qos,
  input  [3:0] io_enq_bits_region,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output  io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos,
  output [3:0] io_deq_bits_region,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [31:0] ram_addr [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_addr_T_144_data;
  wire  ram_addr_T_144_addr;
  wire  ram_addr_T_144_en;
  wire [31:0] ram_addr_T_125_data;
  wire  ram_addr_T_125_addr;
  wire  ram_addr_T_125_mask;
  wire  ram_addr_T_125_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] GEN_1;
  wire [7:0] ram_len_T_144_data;
  wire  ram_len_T_144_addr;
  wire  ram_len_T_144_en;
  wire [7:0] ram_len_T_125_data;
  wire  ram_len_T_125_addr;
  wire  ram_len_T_125_mask;
  wire  ram_len_T_125_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_size_T_144_data;
  wire  ram_size_T_144_addr;
  wire  ram_size_T_144_en;
  wire [2:0] ram_size_T_125_data;
  wire  ram_size_T_125_addr;
  wire  ram_size_T_125_mask;
  wire  ram_size_T_125_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_burst_T_144_data;
  wire  ram_burst_T_144_addr;
  wire  ram_burst_T_144_en;
  wire [1:0] ram_burst_T_125_data;
  wire  ram_burst_T_125_addr;
  wire  ram_burst_T_125_mask;
  wire  ram_burst_T_125_en;
  reg  ram_lock [0:0];
  reg [31:0] GEN_4;
  wire  ram_lock_T_144_data;
  wire  ram_lock_T_144_addr;
  wire  ram_lock_T_144_en;
  wire  ram_lock_T_125_data;
  wire  ram_lock_T_125_addr;
  wire  ram_lock_T_125_mask;
  wire  ram_lock_T_125_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] GEN_5;
  wire [3:0] ram_cache_T_144_data;
  wire  ram_cache_T_144_addr;
  wire  ram_cache_T_144_en;
  wire [3:0] ram_cache_T_125_data;
  wire  ram_cache_T_125_addr;
  wire  ram_cache_T_125_mask;
  wire  ram_cache_T_125_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_prot_T_144_data;
  wire  ram_prot_T_144_addr;
  wire  ram_prot_T_144_en;
  wire [2:0] ram_prot_T_125_data;
  wire  ram_prot_T_125_addr;
  wire  ram_prot_T_125_mask;
  wire  ram_prot_T_125_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] GEN_7;
  wire [3:0] ram_qos_T_144_data;
  wire  ram_qos_T_144_addr;
  wire  ram_qos_T_144_en;
  wire [3:0] ram_qos_T_125_data;
  wire  ram_qos_T_125_addr;
  wire  ram_qos_T_125_mask;
  wire  ram_qos_T_125_en;
  reg [3:0] ram_region [0:0];
  reg [31:0] GEN_8;
  wire [3:0] ram_region_T_144_data;
  wire  ram_region_T_144_addr;
  wire  ram_region_T_144_en;
  wire [3:0] ram_region_T_125_data;
  wire  ram_region_T_125_addr;
  wire  ram_region_T_125_mask;
  wire  ram_region_T_125_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_9;
  wire [4:0] ram_id_T_144_data;
  wire  ram_id_T_144_addr;
  wire  ram_id_T_144_en;
  wire [4:0] ram_id_T_125_data;
  wire  ram_id_T_125_addr;
  wire  ram_id_T_125_mask;
  wire  ram_id_T_125_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_10;
  wire  ram_user_T_144_data;
  wire  ram_user_T_144_addr;
  wire  ram_user_T_144_en;
  wire  ram_user_T_125_data;
  wire  ram_user_T_125_addr;
  wire  ram_user_T_125_mask;
  wire  ram_user_T_125_en;
  reg  maybe_full;
  reg [31:0] GEN_11;
  wire  T_122;
  wire  T_123;
  wire  do_enq;
  wire  T_124;
  wire  do_deq;
  wire  T_139;
  wire  GEN_25;
  wire  T_141;
  wire [1:0] T_156;
  wire  ptr_diff;
  wire [1:0] T_158;
  assign io_enq_ready = T_122;
  assign io_deq_valid = T_141;
  assign io_deq_bits_addr = ram_addr_T_144_data;
  assign io_deq_bits_len = ram_len_T_144_data;
  assign io_deq_bits_size = ram_size_T_144_data;
  assign io_deq_bits_burst = ram_burst_T_144_data;
  assign io_deq_bits_lock = ram_lock_T_144_data;
  assign io_deq_bits_cache = ram_cache_T_144_data;
  assign io_deq_bits_prot = ram_prot_T_144_data;
  assign io_deq_bits_qos = ram_qos_T_144_data;
  assign io_deq_bits_region = ram_region_T_144_data;
  assign io_deq_bits_id = ram_id_T_144_data;
  assign io_deq_bits_user = ram_user_T_144_data;
  assign io_count = T_158[0];
  assign ram_addr_T_144_addr = 1'h0;
  assign ram_addr_T_144_en = 1'h1;
  assign ram_addr_T_144_data = ram_addr[ram_addr_T_144_addr];
  assign ram_addr_T_125_data = io_enq_bits_addr;
  assign ram_addr_T_125_addr = 1'h0;
  assign ram_addr_T_125_mask = do_enq;
  assign ram_addr_T_125_en = do_enq;
  assign ram_len_T_144_addr = 1'h0;
  assign ram_len_T_144_en = 1'h1;
  assign ram_len_T_144_data = ram_len[ram_len_T_144_addr];
  assign ram_len_T_125_data = io_enq_bits_len;
  assign ram_len_T_125_addr = 1'h0;
  assign ram_len_T_125_mask = do_enq;
  assign ram_len_T_125_en = do_enq;
  assign ram_size_T_144_addr = 1'h0;
  assign ram_size_T_144_en = 1'h1;
  assign ram_size_T_144_data = ram_size[ram_size_T_144_addr];
  assign ram_size_T_125_data = io_enq_bits_size;
  assign ram_size_T_125_addr = 1'h0;
  assign ram_size_T_125_mask = do_enq;
  assign ram_size_T_125_en = do_enq;
  assign ram_burst_T_144_addr = 1'h0;
  assign ram_burst_T_144_en = 1'h1;
  assign ram_burst_T_144_data = ram_burst[ram_burst_T_144_addr];
  assign ram_burst_T_125_data = io_enq_bits_burst;
  assign ram_burst_T_125_addr = 1'h0;
  assign ram_burst_T_125_mask = do_enq;
  assign ram_burst_T_125_en = do_enq;
  assign ram_lock_T_144_addr = 1'h0;
  assign ram_lock_T_144_en = 1'h1;
  assign ram_lock_T_144_data = ram_lock[ram_lock_T_144_addr];
  assign ram_lock_T_125_data = io_enq_bits_lock;
  assign ram_lock_T_125_addr = 1'h0;
  assign ram_lock_T_125_mask = do_enq;
  assign ram_lock_T_125_en = do_enq;
  assign ram_cache_T_144_addr = 1'h0;
  assign ram_cache_T_144_en = 1'h1;
  assign ram_cache_T_144_data = ram_cache[ram_cache_T_144_addr];
  assign ram_cache_T_125_data = io_enq_bits_cache;
  assign ram_cache_T_125_addr = 1'h0;
  assign ram_cache_T_125_mask = do_enq;
  assign ram_cache_T_125_en = do_enq;
  assign ram_prot_T_144_addr = 1'h0;
  assign ram_prot_T_144_en = 1'h1;
  assign ram_prot_T_144_data = ram_prot[ram_prot_T_144_addr];
  assign ram_prot_T_125_data = io_enq_bits_prot;
  assign ram_prot_T_125_addr = 1'h0;
  assign ram_prot_T_125_mask = do_enq;
  assign ram_prot_T_125_en = do_enq;
  assign ram_qos_T_144_addr = 1'h0;
  assign ram_qos_T_144_en = 1'h1;
  assign ram_qos_T_144_data = ram_qos[ram_qos_T_144_addr];
  assign ram_qos_T_125_data = io_enq_bits_qos;
  assign ram_qos_T_125_addr = 1'h0;
  assign ram_qos_T_125_mask = do_enq;
  assign ram_qos_T_125_en = do_enq;
  assign ram_region_T_144_addr = 1'h0;
  assign ram_region_T_144_en = 1'h1;
  assign ram_region_T_144_data = ram_region[ram_region_T_144_addr];
  assign ram_region_T_125_data = io_enq_bits_region;
  assign ram_region_T_125_addr = 1'h0;
  assign ram_region_T_125_mask = do_enq;
  assign ram_region_T_125_en = do_enq;
  assign ram_id_T_144_addr = 1'h0;
  assign ram_id_T_144_en = 1'h1;
  assign ram_id_T_144_data = ram_id[ram_id_T_144_addr];
  assign ram_id_T_125_data = io_enq_bits_id;
  assign ram_id_T_125_addr = 1'h0;
  assign ram_id_T_125_mask = do_enq;
  assign ram_id_T_125_en = do_enq;
  assign ram_user_T_144_addr = 1'h0;
  assign ram_user_T_144_en = 1'h1;
  assign ram_user_T_144_data = ram_user[ram_user_T_144_addr];
  assign ram_user_T_125_data = io_enq_bits_user;
  assign ram_user_T_125_addr = 1'h0;
  assign ram_user_T_125_mask = do_enq;
  assign ram_user_T_125_en = do_enq;
  assign T_122 = maybe_full == 1'h0;
  assign T_123 = io_enq_ready & io_enq_valid;
  assign do_enq = T_123;
  assign T_124 = io_deq_ready & io_deq_valid;
  assign do_deq = T_124;
  assign T_139 = do_enq != do_deq;
  assign GEN_25 = T_139 ? do_enq : maybe_full;
  assign T_141 = T_122 == 1'h0;
  assign T_156 = 1'h0 - 1'h0;
  assign ptr_diff = T_156[0:0];
  assign T_158 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[31:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = GEN_1[7:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = GEN_3[1:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = GEN_5[3:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = GEN_7[3:0];
  `endif
  GEN_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_region[initvar] = GEN_8[3:0];
  `endif
  GEN_9 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_9[4:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_10[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_11 = {1{$random}};
  maybe_full = GEN_11[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_125_en & ram_addr_T_125_mask) begin
      ram_addr[ram_addr_T_125_addr] <= ram_addr_T_125_data;
    end
    if(ram_len_T_125_en & ram_len_T_125_mask) begin
      ram_len[ram_len_T_125_addr] <= ram_len_T_125_data;
    end
    if(ram_size_T_125_en & ram_size_T_125_mask) begin
      ram_size[ram_size_T_125_addr] <= ram_size_T_125_data;
    end
    if(ram_burst_T_125_en & ram_burst_T_125_mask) begin
      ram_burst[ram_burst_T_125_addr] <= ram_burst_T_125_data;
    end
    if(ram_lock_T_125_en & ram_lock_T_125_mask) begin
      ram_lock[ram_lock_T_125_addr] <= ram_lock_T_125_data;
    end
    if(ram_cache_T_125_en & ram_cache_T_125_mask) begin
      ram_cache[ram_cache_T_125_addr] <= ram_cache_T_125_data;
    end
    if(ram_prot_T_125_en & ram_prot_T_125_mask) begin
      ram_prot[ram_prot_T_125_addr] <= ram_prot_T_125_data;
    end
    if(ram_qos_T_125_en & ram_qos_T_125_mask) begin
      ram_qos[ram_qos_T_125_addr] <= ram_qos_T_125_data;
    end
    if(ram_region_T_125_en & ram_region_T_125_mask) begin
      ram_region[ram_region_T_125_addr] <= ram_region_T_125_data;
    end
    if(ram_id_T_125_en & ram_id_T_125_mask) begin
      ram_id[ram_id_T_125_addr] <= ram_id_T_125_data;
    end
    if(ram_user_T_125_en & ram_user_T_125_mask) begin
      ram_user[ram_user_T_125_addr] <= ram_user_T_125_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_21(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input  [7:0] io_enq_bits_strb,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output [7:0] io_deq_bits_strb,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_0;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_1;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_2;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] GEN_3;
  wire [7:0] ram_strb_T_94_data;
  wire  ram_strb_T_94_addr;
  wire  ram_strb_T_94_en;
  wire [7:0] ram_strb_T_73_data;
  wire  ram_strb_T_73_addr;
  wire  ram_strb_T_73_mask;
  wire  ram_strb_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_strb = ram_strb_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_strb_T_94_addr = T_67;
  assign ram_strb_T_94_en = 1'h1;
  assign ram_strb_T_94_data = ram_strb[ram_strb_T_94_addr];
  assign ram_strb_T_73_data = io_enq_bits_strb;
  assign ram_strb_T_73_addr = T_65;
  assign ram_strb_T_73_mask = do_enq;
  assign ram_strb_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_0[63:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_1[0:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_2[4:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = GEN_3[7:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_strb_T_73_en & ram_strb_T_73_mask) begin
      ram_strb[ram_strb_T_73_addr] <= ram_strb_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_22(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [1:0] ram_resp [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_94_data;
  wire  ram_resp_T_94_addr;
  wire  ram_resp_T_94_en;
  wire [1:0] ram_resp_T_73_data;
  wire  ram_resp_T_73_addr;
  wire  ram_resp_T_73_mask;
  wire  ram_resp_T_73_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_1;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_2;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_3;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_resp = ram_resp_T_94_data;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_resp_T_94_addr = T_67;
  assign ram_resp_T_94_en = 1'h1;
  assign ram_resp_T_94_data = ram_resp[ram_resp_T_94_addr];
  assign ram_resp_T_73_data = io_enq_bits_resp;
  assign ram_resp_T_73_addr = T_65;
  assign ram_resp_T_73_mask = do_enq;
  assign ram_resp_T_73_en = do_enq;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_1[63:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_3[4:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_73_en & ram_resp_T_73_mask) begin
      ram_resp[ram_resp_T_73_addr] <= ram_resp_T_73_data;
    end
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_23(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [1:0] ram_resp [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_64_data;
  wire  ram_resp_T_64_addr;
  wire  ram_resp_T_64_en;
  wire [1:0] ram_resp_T_53_data;
  wire  ram_resp_T_53_addr;
  wire  ram_resp_T_53_mask;
  wire  ram_resp_T_53_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_1;
  wire [4:0] ram_id_T_64_data;
  wire  ram_id_T_64_addr;
  wire  ram_id_T_64_en;
  wire [4:0] ram_id_T_53_data;
  wire  ram_id_T_53_addr;
  wire  ram_id_T_53_mask;
  wire  ram_id_T_53_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_2;
  wire  ram_user_T_64_data;
  wire  ram_user_T_64_addr;
  wire  ram_user_T_64_en;
  wire  ram_user_T_53_data;
  wire  ram_user_T_53_addr;
  wire  ram_user_T_53_mask;
  wire  ram_user_T_53_en;
  reg  maybe_full;
  reg [31:0] GEN_3;
  wire  T_50;
  wire  T_51;
  wire  do_enq;
  wire  T_52;
  wire  do_deq;
  wire  T_59;
  wire  GEN_9;
  wire  T_61;
  wire [1:0] T_68;
  wire  ptr_diff;
  wire [1:0] T_70;
  assign io_enq_ready = T_50;
  assign io_deq_valid = T_61;
  assign io_deq_bits_resp = ram_resp_T_64_data;
  assign io_deq_bits_id = ram_id_T_64_data;
  assign io_deq_bits_user = ram_user_T_64_data;
  assign io_count = T_70[0];
  assign ram_resp_T_64_addr = 1'h0;
  assign ram_resp_T_64_en = 1'h1;
  assign ram_resp_T_64_data = ram_resp[ram_resp_T_64_addr];
  assign ram_resp_T_53_data = io_enq_bits_resp;
  assign ram_resp_T_53_addr = 1'h0;
  assign ram_resp_T_53_mask = do_enq;
  assign ram_resp_T_53_en = do_enq;
  assign ram_id_T_64_addr = 1'h0;
  assign ram_id_T_64_en = 1'h1;
  assign ram_id_T_64_data = ram_id[ram_id_T_64_addr];
  assign ram_id_T_53_data = io_enq_bits_id;
  assign ram_id_T_53_addr = 1'h0;
  assign ram_id_T_53_mask = do_enq;
  assign ram_id_T_53_en = do_enq;
  assign ram_user_T_64_addr = 1'h0;
  assign ram_user_T_64_en = 1'h1;
  assign ram_user_T_64_data = ram_user[ram_user_T_64_addr];
  assign ram_user_T_53_data = io_enq_bits_user;
  assign ram_user_T_53_addr = 1'h0;
  assign ram_user_T_53_mask = do_enq;
  assign ram_user_T_53_en = do_enq;
  assign T_50 = maybe_full == 1'h0;
  assign T_51 = io_enq_ready & io_enq_valid;
  assign do_enq = T_51;
  assign T_52 = io_deq_ready & io_deq_valid;
  assign do_deq = T_52;
  assign T_59 = do_enq != do_deq;
  assign GEN_9 = T_59 ? do_enq : maybe_full;
  assign T_61 = T_50 == 1'h0;
  assign T_68 = 1'h0 - 1'h0;
  assign ptr_diff = T_68[0:0];
  assign T_70 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_1[4:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_3 = {1{$random}};
  maybe_full = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_53_en & ram_resp_T_53_mask) begin
      ram_resp[ram_resp_T_53_addr] <= ram_resp_T_53_data;
    end
    if(ram_id_T_53_en & ram_id_T_53_mask) begin
      ram_id[ram_id_T_53_addr] <= ram_id_T_53_data;
    end
    if(ram_user_T_53_en & ram_user_T_53_mask) begin
      ram_user[ram_user_T_53_addr] <= ram_user_T_53_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_59) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Periphery(
  input   clk,
  input   reset,
  output  io_mem_in_0_acquire_ready,
  input   io_mem_in_0_acquire_valid,
  input  [25:0] io_mem_in_0_acquire_bits_addr_block,
  input  [2:0] io_mem_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_mem_in_0_acquire_bits_addr_beat,
  input   io_mem_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_mem_in_0_acquire_bits_a_type,
  input  [10:0] io_mem_in_0_acquire_bits_union,
  input  [63:0] io_mem_in_0_acquire_bits_data,
  input   io_mem_in_0_grant_ready,
  output  io_mem_in_0_grant_valid,
  output [2:0] io_mem_in_0_grant_bits_addr_beat,
  output [2:0] io_mem_in_0_grant_bits_client_xact_id,
  output  io_mem_in_0_grant_bits_manager_xact_id,
  output  io_mem_in_0_grant_bits_is_builtin_type,
  output [3:0] io_mem_in_0_grant_bits_g_type,
  output [63:0] io_mem_in_0_grant_bits_data,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user
);
  wire  NastiIOTileLinkIOConverter_1_clk;
  wire  NastiIOTileLinkIOConverter_1_reset;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type;
  wire [10:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user;
  wire  Queue_19_1_clk;
  wire  Queue_19_1_reset;
  wire  Queue_19_1_io_enq_ready;
  wire  Queue_19_1_io_enq_valid;
  wire [31:0] Queue_19_1_io_enq_bits_addr;
  wire [7:0] Queue_19_1_io_enq_bits_len;
  wire [2:0] Queue_19_1_io_enq_bits_size;
  wire [1:0] Queue_19_1_io_enq_bits_burst;
  wire  Queue_19_1_io_enq_bits_lock;
  wire [3:0] Queue_19_1_io_enq_bits_cache;
  wire [2:0] Queue_19_1_io_enq_bits_prot;
  wire [3:0] Queue_19_1_io_enq_bits_qos;
  wire [3:0] Queue_19_1_io_enq_bits_region;
  wire [4:0] Queue_19_1_io_enq_bits_id;
  wire  Queue_19_1_io_enq_bits_user;
  wire  Queue_19_1_io_deq_ready;
  wire  Queue_19_1_io_deq_valid;
  wire [31:0] Queue_19_1_io_deq_bits_addr;
  wire [7:0] Queue_19_1_io_deq_bits_len;
  wire [2:0] Queue_19_1_io_deq_bits_size;
  wire [1:0] Queue_19_1_io_deq_bits_burst;
  wire  Queue_19_1_io_deq_bits_lock;
  wire [3:0] Queue_19_1_io_deq_bits_cache;
  wire [2:0] Queue_19_1_io_deq_bits_prot;
  wire [3:0] Queue_19_1_io_deq_bits_qos;
  wire [3:0] Queue_19_1_io_deq_bits_region;
  wire [4:0] Queue_19_1_io_deq_bits_id;
  wire  Queue_19_1_io_deq_bits_user;
  wire  Queue_19_1_io_count;
  wire  Queue_20_1_clk;
  wire  Queue_20_1_reset;
  wire  Queue_20_1_io_enq_ready;
  wire  Queue_20_1_io_enq_valid;
  wire [31:0] Queue_20_1_io_enq_bits_addr;
  wire [7:0] Queue_20_1_io_enq_bits_len;
  wire [2:0] Queue_20_1_io_enq_bits_size;
  wire [1:0] Queue_20_1_io_enq_bits_burst;
  wire  Queue_20_1_io_enq_bits_lock;
  wire [3:0] Queue_20_1_io_enq_bits_cache;
  wire [2:0] Queue_20_1_io_enq_bits_prot;
  wire [3:0] Queue_20_1_io_enq_bits_qos;
  wire [3:0] Queue_20_1_io_enq_bits_region;
  wire [4:0] Queue_20_1_io_enq_bits_id;
  wire  Queue_20_1_io_enq_bits_user;
  wire  Queue_20_1_io_deq_ready;
  wire  Queue_20_1_io_deq_valid;
  wire [31:0] Queue_20_1_io_deq_bits_addr;
  wire [7:0] Queue_20_1_io_deq_bits_len;
  wire [2:0] Queue_20_1_io_deq_bits_size;
  wire [1:0] Queue_20_1_io_deq_bits_burst;
  wire  Queue_20_1_io_deq_bits_lock;
  wire [3:0] Queue_20_1_io_deq_bits_cache;
  wire [2:0] Queue_20_1_io_deq_bits_prot;
  wire [3:0] Queue_20_1_io_deq_bits_qos;
  wire [3:0] Queue_20_1_io_deq_bits_region;
  wire [4:0] Queue_20_1_io_deq_bits_id;
  wire  Queue_20_1_io_deq_bits_user;
  wire  Queue_20_1_io_count;
  wire  Queue_21_1_clk;
  wire  Queue_21_1_reset;
  wire  Queue_21_1_io_enq_ready;
  wire  Queue_21_1_io_enq_valid;
  wire [63:0] Queue_21_1_io_enq_bits_data;
  wire  Queue_21_1_io_enq_bits_last;
  wire [4:0] Queue_21_1_io_enq_bits_id;
  wire [7:0] Queue_21_1_io_enq_bits_strb;
  wire  Queue_21_1_io_enq_bits_user;
  wire  Queue_21_1_io_deq_ready;
  wire  Queue_21_1_io_deq_valid;
  wire [63:0] Queue_21_1_io_deq_bits_data;
  wire  Queue_21_1_io_deq_bits_last;
  wire [4:0] Queue_21_1_io_deq_bits_id;
  wire [7:0] Queue_21_1_io_deq_bits_strb;
  wire  Queue_21_1_io_deq_bits_user;
  wire [1:0] Queue_21_1_io_count;
  wire  Queue_22_1_clk;
  wire  Queue_22_1_reset;
  wire  Queue_22_1_io_enq_ready;
  wire  Queue_22_1_io_enq_valid;
  wire [1:0] Queue_22_1_io_enq_bits_resp;
  wire [63:0] Queue_22_1_io_enq_bits_data;
  wire  Queue_22_1_io_enq_bits_last;
  wire [4:0] Queue_22_1_io_enq_bits_id;
  wire  Queue_22_1_io_enq_bits_user;
  wire  Queue_22_1_io_deq_ready;
  wire  Queue_22_1_io_deq_valid;
  wire [1:0] Queue_22_1_io_deq_bits_resp;
  wire [63:0] Queue_22_1_io_deq_bits_data;
  wire  Queue_22_1_io_deq_bits_last;
  wire [4:0] Queue_22_1_io_deq_bits_id;
  wire  Queue_22_1_io_deq_bits_user;
  wire [1:0] Queue_22_1_io_count;
  wire  Queue_23_1_clk;
  wire  Queue_23_1_reset;
  wire  Queue_23_1_io_enq_ready;
  wire  Queue_23_1_io_enq_valid;
  wire [1:0] Queue_23_1_io_enq_bits_resp;
  wire [4:0] Queue_23_1_io_enq_bits_id;
  wire  Queue_23_1_io_enq_bits_user;
  wire  Queue_23_1_io_deq_ready;
  wire  Queue_23_1_io_deq_valid;
  wire [1:0] Queue_23_1_io_deq_bits_resp;
  wire [4:0] Queue_23_1_io_deq_bits_id;
  wire  Queue_23_1_io_deq_bits_user;
  wire  Queue_23_1_io_count;
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter_1 (
    .clk(NastiIOTileLinkIOConverter_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user)
  );
  Queue_19 Queue_19_1 (
    .clk(Queue_19_1_clk),
    .reset(Queue_19_1_reset),
    .io_enq_ready(Queue_19_1_io_enq_ready),
    .io_enq_valid(Queue_19_1_io_enq_valid),
    .io_enq_bits_addr(Queue_19_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_19_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_19_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_19_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_19_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_19_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_19_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_19_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_19_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_19_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_19_1_io_enq_bits_user),
    .io_deq_ready(Queue_19_1_io_deq_ready),
    .io_deq_valid(Queue_19_1_io_deq_valid),
    .io_deq_bits_addr(Queue_19_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_19_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_19_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_19_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_19_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_19_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_19_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_19_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_19_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_19_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_19_1_io_deq_bits_user),
    .io_count(Queue_19_1_io_count)
  );
  Queue_19 Queue_20_1 (
    .clk(Queue_20_1_clk),
    .reset(Queue_20_1_reset),
    .io_enq_ready(Queue_20_1_io_enq_ready),
    .io_enq_valid(Queue_20_1_io_enq_valid),
    .io_enq_bits_addr(Queue_20_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_20_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_20_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_20_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_20_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_20_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_20_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_20_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_20_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_20_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_20_1_io_enq_bits_user),
    .io_deq_ready(Queue_20_1_io_deq_ready),
    .io_deq_valid(Queue_20_1_io_deq_valid),
    .io_deq_bits_addr(Queue_20_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_20_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_20_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_20_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_20_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_20_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_20_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_20_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_20_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_20_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_20_1_io_deq_bits_user),
    .io_count(Queue_20_1_io_count)
  );
  Queue_21 Queue_21_1 (
    .clk(Queue_21_1_clk),
    .reset(Queue_21_1_reset),
    .io_enq_ready(Queue_21_1_io_enq_ready),
    .io_enq_valid(Queue_21_1_io_enq_valid),
    .io_enq_bits_data(Queue_21_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_21_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_21_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_21_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_21_1_io_enq_bits_user),
    .io_deq_ready(Queue_21_1_io_deq_ready),
    .io_deq_valid(Queue_21_1_io_deq_valid),
    .io_deq_bits_data(Queue_21_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_21_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_21_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_21_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_21_1_io_deq_bits_user),
    .io_count(Queue_21_1_io_count)
  );
  Queue_22 Queue_22_1 (
    .clk(Queue_22_1_clk),
    .reset(Queue_22_1_reset),
    .io_enq_ready(Queue_22_1_io_enq_ready),
    .io_enq_valid(Queue_22_1_io_enq_valid),
    .io_enq_bits_resp(Queue_22_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_22_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_22_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_22_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_22_1_io_enq_bits_user),
    .io_deq_ready(Queue_22_1_io_deq_ready),
    .io_deq_valid(Queue_22_1_io_deq_valid),
    .io_deq_bits_resp(Queue_22_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_22_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_22_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_22_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_22_1_io_deq_bits_user),
    .io_count(Queue_22_1_io_count)
  );
  Queue_23 Queue_23_1 (
    .clk(Queue_23_1_clk),
    .reset(Queue_23_1_reset),
    .io_enq_ready(Queue_23_1_io_enq_ready),
    .io_enq_valid(Queue_23_1_io_enq_valid),
    .io_enq_bits_resp(Queue_23_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_23_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_23_1_io_enq_bits_user),
    .io_deq_ready(Queue_23_1_io_deq_ready),
    .io_deq_valid(Queue_23_1_io_deq_valid),
    .io_deq_bits_resp(Queue_23_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_23_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_23_1_io_deq_bits_user),
    .io_count(Queue_23_1_io_count)
  );
  assign io_mem_in_0_acquire_ready = NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  assign io_mem_in_0_grant_valid = NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  assign io_mem_in_0_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  assign io_mem_in_0_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  assign io_mem_in_0_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  assign io_mem_in_0_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  assign io_mem_in_0_grant_bits_g_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  assign io_mem_in_0_grant_bits_data = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  assign io_mem_axi_0_aw_valid = Queue_20_1_io_deq_valid;
  assign io_mem_axi_0_aw_bits_addr = Queue_20_1_io_deq_bits_addr;
  assign io_mem_axi_0_aw_bits_len = Queue_20_1_io_deq_bits_len;
  assign io_mem_axi_0_aw_bits_size = Queue_20_1_io_deq_bits_size;
  assign io_mem_axi_0_aw_bits_burst = Queue_20_1_io_deq_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = Queue_20_1_io_deq_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = 4'h3;
  assign io_mem_axi_0_aw_bits_prot = Queue_20_1_io_deq_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = Queue_20_1_io_deq_bits_qos;
  assign io_mem_axi_0_aw_bits_region = Queue_20_1_io_deq_bits_region;
  assign io_mem_axi_0_aw_bits_id = Queue_20_1_io_deq_bits_id;
  assign io_mem_axi_0_aw_bits_user = Queue_20_1_io_deq_bits_user;
  assign io_mem_axi_0_w_valid = Queue_21_1_io_deq_valid;
  assign io_mem_axi_0_w_bits_data = Queue_21_1_io_deq_bits_data;
  assign io_mem_axi_0_w_bits_last = Queue_21_1_io_deq_bits_last;
  assign io_mem_axi_0_w_bits_id = Queue_21_1_io_deq_bits_id;
  assign io_mem_axi_0_w_bits_strb = Queue_21_1_io_deq_bits_strb;
  assign io_mem_axi_0_w_bits_user = Queue_21_1_io_deq_bits_user;
  assign io_mem_axi_0_b_ready = Queue_23_1_io_enq_ready;
  assign io_mem_axi_0_ar_valid = Queue_19_1_io_deq_valid;
  assign io_mem_axi_0_ar_bits_addr = Queue_19_1_io_deq_bits_addr;
  assign io_mem_axi_0_ar_bits_len = Queue_19_1_io_deq_bits_len;
  assign io_mem_axi_0_ar_bits_size = Queue_19_1_io_deq_bits_size;
  assign io_mem_axi_0_ar_bits_burst = Queue_19_1_io_deq_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = Queue_19_1_io_deq_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = 4'h3;
  assign io_mem_axi_0_ar_bits_prot = Queue_19_1_io_deq_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = Queue_19_1_io_deq_bits_qos;
  assign io_mem_axi_0_ar_bits_region = Queue_19_1_io_deq_bits_region;
  assign io_mem_axi_0_ar_bits_id = Queue_19_1_io_deq_bits_id;
  assign io_mem_axi_0_ar_bits_user = Queue_19_1_io_deq_bits_user;
  assign io_mem_axi_0_r_ready = Queue_22_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_valid = io_mem_in_0_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block = io_mem_in_0_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id = io_mem_in_0_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat = io_mem_in_0_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type = io_mem_in_0_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type = io_mem_in_0_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union = io_mem_in_0_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data = io_mem_in_0_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_tl_grant_ready = io_mem_in_0_grant_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_aw_ready = Queue_20_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_w_ready = Queue_21_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_valid = Queue_23_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp = Queue_23_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id = Queue_23_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user = Queue_23_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_io_nasti_ar_ready = Queue_19_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_valid = Queue_22_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp = Queue_22_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data = Queue_22_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last = Queue_22_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id = Queue_22_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user = Queue_22_1_io_deq_bits_user;
  assign Queue_19_1_clk = clk;
  assign Queue_19_1_reset = reset;
  assign Queue_19_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  assign Queue_19_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  assign Queue_19_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  assign Queue_19_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  assign Queue_19_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  assign Queue_19_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  assign Queue_19_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  assign Queue_19_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  assign Queue_19_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  assign Queue_19_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  assign Queue_19_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  assign Queue_19_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  assign Queue_19_1_io_deq_ready = io_mem_axi_0_ar_ready;
  assign Queue_20_1_clk = clk;
  assign Queue_20_1_reset = reset;
  assign Queue_20_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  assign Queue_20_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  assign Queue_20_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  assign Queue_20_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  assign Queue_20_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  assign Queue_20_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  assign Queue_20_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  assign Queue_20_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  assign Queue_20_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  assign Queue_20_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  assign Queue_20_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  assign Queue_20_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  assign Queue_20_1_io_deq_ready = io_mem_axi_0_aw_ready;
  assign Queue_21_1_clk = clk;
  assign Queue_21_1_reset = reset;
  assign Queue_21_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  assign Queue_21_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  assign Queue_21_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  assign Queue_21_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  assign Queue_21_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  assign Queue_21_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  assign Queue_21_1_io_deq_ready = io_mem_axi_0_w_ready;
  assign Queue_22_1_clk = clk;
  assign Queue_22_1_reset = reset;
  assign Queue_22_1_io_enq_valid = io_mem_axi_0_r_valid;
  assign Queue_22_1_io_enq_bits_resp = io_mem_axi_0_r_bits_resp;
  assign Queue_22_1_io_enq_bits_data = io_mem_axi_0_r_bits_data;
  assign Queue_22_1_io_enq_bits_last = io_mem_axi_0_r_bits_last;
  assign Queue_22_1_io_enq_bits_id = io_mem_axi_0_r_bits_id;
  assign Queue_22_1_io_enq_bits_user = io_mem_axi_0_r_bits_user;
  assign Queue_22_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  assign Queue_23_1_clk = clk;
  assign Queue_23_1_reset = reset;
  assign Queue_23_1_io_enq_valid = io_mem_axi_0_b_valid;
  assign Queue_23_1_io_enq_bits_resp = io_mem_axi_0_b_bits_resp;
  assign Queue_23_1_io_enq_bits_id = io_mem_axi_0_b_bits_id;
  assign Queue_23_1_io_enq_bits_user = io_mem_axi_0_b_bits_user;
  assign Queue_23_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
endmodule
module Top_1(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [33:0] io_debug_req_bits_data,
  input  [1:0] io_debug_req_bits_op,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [33:0] io_debug_resp_bits_data,
  output [1:0] io_debug_resp_bits_resp
);
  wire  coreplex_clk;
  wire  coreplex_reset;
  wire  coreplex_io_mem_0_acquire_ready;
  wire  coreplex_io_mem_0_acquire_valid;
  wire [25:0] coreplex_io_mem_0_acquire_bits_addr_block;
  wire [2:0] coreplex_io_mem_0_acquire_bits_client_xact_id;
  wire [2:0] coreplex_io_mem_0_acquire_bits_addr_beat;
  wire  coreplex_io_mem_0_acquire_bits_is_builtin_type;
  wire [2:0] coreplex_io_mem_0_acquire_bits_a_type;
  wire [10:0] coreplex_io_mem_0_acquire_bits_union;
  wire [63:0] coreplex_io_mem_0_acquire_bits_data;
  wire  coreplex_io_mem_0_grant_ready;
  wire  coreplex_io_mem_0_grant_valid;
  wire [2:0] coreplex_io_mem_0_grant_bits_addr_beat;
  wire [2:0] coreplex_io_mem_0_grant_bits_client_xact_id;
  wire  coreplex_io_mem_0_grant_bits_manager_xact_id;
  wire  coreplex_io_mem_0_grant_bits_is_builtin_type;
  wire [3:0] coreplex_io_mem_0_grant_bits_g_type;
  wire [63:0] coreplex_io_mem_0_grant_bits_data;
  wire  coreplex_io_interrupts_0;
  wire  coreplex_io_interrupts_1;
  wire  coreplex_io_debug_req_ready;
  wire  coreplex_io_debug_req_valid;
  wire [4:0] coreplex_io_debug_req_bits_addr;
  wire [33:0] coreplex_io_debug_req_bits_data;
  wire [1:0] coreplex_io_debug_req_bits_op;
  wire  coreplex_io_debug_resp_ready;
  wire  coreplex_io_debug_resp_valid;
  wire [33:0] coreplex_io_debug_resp_bits_data;
  wire [1:0] coreplex_io_debug_resp_bits_resp;
  wire  coreplex_io_rtcTick;
  wire  periphery_clk;
  wire  periphery_reset;
  wire  periphery_io_mem_in_0_acquire_ready;
  wire  periphery_io_mem_in_0_acquire_valid;
  wire [25:0] periphery_io_mem_in_0_acquire_bits_addr_block;
  wire [2:0] periphery_io_mem_in_0_acquire_bits_client_xact_id;
  wire [2:0] periphery_io_mem_in_0_acquire_bits_addr_beat;
  wire  periphery_io_mem_in_0_acquire_bits_is_builtin_type;
  wire [2:0] periphery_io_mem_in_0_acquire_bits_a_type;
  wire [10:0] periphery_io_mem_in_0_acquire_bits_union;
  wire [63:0] periphery_io_mem_in_0_acquire_bits_data;
  wire  periphery_io_mem_in_0_grant_ready;
  wire  periphery_io_mem_in_0_grant_valid;
  wire [2:0] periphery_io_mem_in_0_grant_bits_addr_beat;
  wire [2:0] periphery_io_mem_in_0_grant_bits_client_xact_id;
  wire  periphery_io_mem_in_0_grant_bits_manager_xact_id;
  wire  periphery_io_mem_in_0_grant_bits_is_builtin_type;
  wire [3:0] periphery_io_mem_in_0_grant_bits_g_type;
  wire [63:0] periphery_io_mem_in_0_grant_bits_data;
  wire  periphery_io_mem_axi_0_aw_ready;
  wire  periphery_io_mem_axi_0_aw_valid;
  wire [31:0] periphery_io_mem_axi_0_aw_bits_addr;
  wire [7:0] periphery_io_mem_axi_0_aw_bits_len;
  wire [2:0] periphery_io_mem_axi_0_aw_bits_size;
  wire [1:0] periphery_io_mem_axi_0_aw_bits_burst;
  wire  periphery_io_mem_axi_0_aw_bits_lock;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_cache;
  wire [2:0] periphery_io_mem_axi_0_aw_bits_prot;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_qos;
  wire [3:0] periphery_io_mem_axi_0_aw_bits_region;
  wire [4:0] periphery_io_mem_axi_0_aw_bits_id;
  wire  periphery_io_mem_axi_0_aw_bits_user;
  wire  periphery_io_mem_axi_0_w_ready;
  wire  periphery_io_mem_axi_0_w_valid;
  wire [63:0] periphery_io_mem_axi_0_w_bits_data;
  wire  periphery_io_mem_axi_0_w_bits_last;
  wire [4:0] periphery_io_mem_axi_0_w_bits_id;
  wire [7:0] periphery_io_mem_axi_0_w_bits_strb;
  wire  periphery_io_mem_axi_0_w_bits_user;
  wire  periphery_io_mem_axi_0_b_ready;
  wire  periphery_io_mem_axi_0_b_valid;
  wire [1:0] periphery_io_mem_axi_0_b_bits_resp;
  wire [4:0] periphery_io_mem_axi_0_b_bits_id;
  wire  periphery_io_mem_axi_0_b_bits_user;
  wire  periphery_io_mem_axi_0_ar_ready;
  wire  periphery_io_mem_axi_0_ar_valid;
  wire [31:0] periphery_io_mem_axi_0_ar_bits_addr;
  wire [7:0] periphery_io_mem_axi_0_ar_bits_len;
  wire [2:0] periphery_io_mem_axi_0_ar_bits_size;
  wire [1:0] periphery_io_mem_axi_0_ar_bits_burst;
  wire  periphery_io_mem_axi_0_ar_bits_lock;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_cache;
  wire [2:0] periphery_io_mem_axi_0_ar_bits_prot;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_qos;
  wire [3:0] periphery_io_mem_axi_0_ar_bits_region;
  wire [4:0] periphery_io_mem_axi_0_ar_bits_id;
  wire  periphery_io_mem_axi_0_ar_bits_user;
  wire  periphery_io_mem_axi_0_r_ready;
  wire  periphery_io_mem_axi_0_r_valid;
  wire [1:0] periphery_io_mem_axi_0_r_bits_resp;
  wire [63:0] periphery_io_mem_axi_0_r_bits_data;
  wire  periphery_io_mem_axi_0_r_bits_last;
  wire [4:0] periphery_io_mem_axi_0_r_bits_id;
  wire  periphery_io_mem_axi_0_r_bits_user;
  reg [6:0] T_3628;
  reg [31:0] GEN_1;
  wire  T_3630;
  wire [7:0] T_3632;
  wire [6:0] T_3633;
  wire [6:0] GEN_0;
  DefaultCoreplex coreplex (
    .clk(coreplex_clk),
    .reset(coreplex_reset),
    .io_mem_0_acquire_ready(coreplex_io_mem_0_acquire_ready),
    .io_mem_0_acquire_valid(coreplex_io_mem_0_acquire_valid),
    .io_mem_0_acquire_bits_addr_block(coreplex_io_mem_0_acquire_bits_addr_block),
    .io_mem_0_acquire_bits_client_xact_id(coreplex_io_mem_0_acquire_bits_client_xact_id),
    .io_mem_0_acquire_bits_addr_beat(coreplex_io_mem_0_acquire_bits_addr_beat),
    .io_mem_0_acquire_bits_is_builtin_type(coreplex_io_mem_0_acquire_bits_is_builtin_type),
    .io_mem_0_acquire_bits_a_type(coreplex_io_mem_0_acquire_bits_a_type),
    .io_mem_0_acquire_bits_union(coreplex_io_mem_0_acquire_bits_union),
    .io_mem_0_acquire_bits_data(coreplex_io_mem_0_acquire_bits_data),
    .io_mem_0_grant_ready(coreplex_io_mem_0_grant_ready),
    .io_mem_0_grant_valid(coreplex_io_mem_0_grant_valid),
    .io_mem_0_grant_bits_addr_beat(coreplex_io_mem_0_grant_bits_addr_beat),
    .io_mem_0_grant_bits_client_xact_id(coreplex_io_mem_0_grant_bits_client_xact_id),
    .io_mem_0_grant_bits_manager_xact_id(coreplex_io_mem_0_grant_bits_manager_xact_id),
    .io_mem_0_grant_bits_is_builtin_type(coreplex_io_mem_0_grant_bits_is_builtin_type),
    .io_mem_0_grant_bits_g_type(coreplex_io_mem_0_grant_bits_g_type),
    .io_mem_0_grant_bits_data(coreplex_io_mem_0_grant_bits_data),
    .io_interrupts_0(coreplex_io_interrupts_0),
    .io_interrupts_1(coreplex_io_interrupts_1),
    .io_debug_req_ready(coreplex_io_debug_req_ready),
    .io_debug_req_valid(coreplex_io_debug_req_valid),
    .io_debug_req_bits_addr(coreplex_io_debug_req_bits_addr),
    .io_debug_req_bits_data(coreplex_io_debug_req_bits_data),
    .io_debug_req_bits_op(coreplex_io_debug_req_bits_op),
    .io_debug_resp_ready(coreplex_io_debug_resp_ready),
    .io_debug_resp_valid(coreplex_io_debug_resp_valid),
    .io_debug_resp_bits_data(coreplex_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(coreplex_io_debug_resp_bits_resp),
    .io_rtcTick(coreplex_io_rtcTick)
  );
  Periphery periphery (
    .clk(periphery_clk),
    .reset(periphery_reset),
    .io_mem_in_0_acquire_ready(periphery_io_mem_in_0_acquire_ready),
    .io_mem_in_0_acquire_valid(periphery_io_mem_in_0_acquire_valid),
    .io_mem_in_0_acquire_bits_addr_block(periphery_io_mem_in_0_acquire_bits_addr_block),
    .io_mem_in_0_acquire_bits_client_xact_id(periphery_io_mem_in_0_acquire_bits_client_xact_id),
    .io_mem_in_0_acquire_bits_addr_beat(periphery_io_mem_in_0_acquire_bits_addr_beat),
    .io_mem_in_0_acquire_bits_is_builtin_type(periphery_io_mem_in_0_acquire_bits_is_builtin_type),
    .io_mem_in_0_acquire_bits_a_type(periphery_io_mem_in_0_acquire_bits_a_type),
    .io_mem_in_0_acquire_bits_union(periphery_io_mem_in_0_acquire_bits_union),
    .io_mem_in_0_acquire_bits_data(periphery_io_mem_in_0_acquire_bits_data),
    .io_mem_in_0_grant_ready(periphery_io_mem_in_0_grant_ready),
    .io_mem_in_0_grant_valid(periphery_io_mem_in_0_grant_valid),
    .io_mem_in_0_grant_bits_addr_beat(periphery_io_mem_in_0_grant_bits_addr_beat),
    .io_mem_in_0_grant_bits_client_xact_id(periphery_io_mem_in_0_grant_bits_client_xact_id),
    .io_mem_in_0_grant_bits_manager_xact_id(periphery_io_mem_in_0_grant_bits_manager_xact_id),
    .io_mem_in_0_grant_bits_is_builtin_type(periphery_io_mem_in_0_grant_bits_is_builtin_type),
    .io_mem_in_0_grant_bits_g_type(periphery_io_mem_in_0_grant_bits_g_type),
    .io_mem_in_0_grant_bits_data(periphery_io_mem_in_0_grant_bits_data),
    .io_mem_axi_0_aw_ready(periphery_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(periphery_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(periphery_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(periphery_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(periphery_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(periphery_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(periphery_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(periphery_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(periphery_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(periphery_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(periphery_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(periphery_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(periphery_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(periphery_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(periphery_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(periphery_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(periphery_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(periphery_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(periphery_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(periphery_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(periphery_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(periphery_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(periphery_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(periphery_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(periphery_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(periphery_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(periphery_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(periphery_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(periphery_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(periphery_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(periphery_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(periphery_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(periphery_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(periphery_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(periphery_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(periphery_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(periphery_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(periphery_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(periphery_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(periphery_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(periphery_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(periphery_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(periphery_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(periphery_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(periphery_io_mem_axi_0_r_bits_user)
  );
  assign io_mem_axi_0_aw_valid = periphery_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = periphery_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = periphery_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = periphery_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = periphery_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = periphery_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = periphery_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = periphery_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = periphery_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = periphery_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = periphery_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = periphery_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = periphery_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = periphery_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = periphery_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = periphery_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = periphery_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = periphery_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = periphery_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = periphery_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = periphery_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = periphery_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = periphery_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = periphery_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = periphery_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = periphery_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = periphery_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = periphery_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = periphery_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = periphery_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = periphery_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = periphery_io_mem_axi_0_r_ready;
  assign io_debug_req_ready = coreplex_io_debug_req_ready;
  assign io_debug_resp_valid = coreplex_io_debug_resp_valid;
  assign io_debug_resp_bits_data = coreplex_io_debug_resp_bits_data;
  assign io_debug_resp_bits_resp = coreplex_io_debug_resp_bits_resp;
  assign coreplex_clk = clk;
  assign coreplex_reset = reset;
  assign coreplex_io_mem_0_acquire_ready = periphery_io_mem_in_0_acquire_ready;
  assign coreplex_io_mem_0_grant_valid = periphery_io_mem_in_0_grant_valid;
  assign coreplex_io_mem_0_grant_bits_addr_beat = periphery_io_mem_in_0_grant_bits_addr_beat;
  assign coreplex_io_mem_0_grant_bits_client_xact_id = periphery_io_mem_in_0_grant_bits_client_xact_id;
  assign coreplex_io_mem_0_grant_bits_manager_xact_id = periphery_io_mem_in_0_grant_bits_manager_xact_id;
  assign coreplex_io_mem_0_grant_bits_is_builtin_type = periphery_io_mem_in_0_grant_bits_is_builtin_type;
  assign coreplex_io_mem_0_grant_bits_g_type = periphery_io_mem_in_0_grant_bits_g_type;
  assign coreplex_io_mem_0_grant_bits_data = periphery_io_mem_in_0_grant_bits_data;
  assign coreplex_io_interrupts_0 = io_interrupts_0;
  assign coreplex_io_interrupts_1 = io_interrupts_1;
  assign coreplex_io_debug_req_valid = io_debug_req_valid;
  assign coreplex_io_debug_req_bits_addr = io_debug_req_bits_addr;
  assign coreplex_io_debug_req_bits_data = io_debug_req_bits_data;
  assign coreplex_io_debug_req_bits_op = io_debug_req_bits_op;
  assign coreplex_io_debug_resp_ready = io_debug_resp_ready;
  assign coreplex_io_rtcTick = T_3630;
  assign periphery_clk = clk;
  assign periphery_reset = reset;
  assign periphery_io_mem_in_0_acquire_valid = coreplex_io_mem_0_acquire_valid;
  assign periphery_io_mem_in_0_acquire_bits_addr_block = coreplex_io_mem_0_acquire_bits_addr_block;
  assign periphery_io_mem_in_0_acquire_bits_client_xact_id = coreplex_io_mem_0_acquire_bits_client_xact_id;
  assign periphery_io_mem_in_0_acquire_bits_addr_beat = coreplex_io_mem_0_acquire_bits_addr_beat;
  assign periphery_io_mem_in_0_acquire_bits_is_builtin_type = coreplex_io_mem_0_acquire_bits_is_builtin_type;
  assign periphery_io_mem_in_0_acquire_bits_a_type = coreplex_io_mem_0_acquire_bits_a_type;
  assign periphery_io_mem_in_0_acquire_bits_union = coreplex_io_mem_0_acquire_bits_union;
  assign periphery_io_mem_in_0_acquire_bits_data = coreplex_io_mem_0_acquire_bits_data;
  assign periphery_io_mem_in_0_grant_ready = coreplex_io_mem_0_grant_ready;
  assign periphery_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign periphery_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign periphery_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign periphery_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign periphery_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign periphery_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign periphery_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign periphery_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign periphery_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign periphery_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign periphery_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign periphery_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign periphery_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign T_3630 = T_3628 == 7'h63;
  assign T_3632 = T_3628 + 7'h1;
  assign T_3633 = T_3632[6:0];
  assign GEN_0 = T_3630 ? 7'h0 : T_3633;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_1 = {1{$random}};
  T_3628 = GEN_1[6:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_3628 <= 7'h0;
    end else begin
      if(T_3630) begin
        T_3628 <= 7'h0;
      end else begin
        T_3628 <= T_3633;
      end
    end
  end
endmodule
module Top(
  input   clk,
  input   reset,
  output  io_ps_axi_slave_aw_ready,
  input   io_ps_axi_slave_aw_valid,
  input  [31:0] io_ps_axi_slave_aw_bits_addr,
  input  [7:0] io_ps_axi_slave_aw_bits_len,
  input  [2:0] io_ps_axi_slave_aw_bits_size,
  input  [1:0] io_ps_axi_slave_aw_bits_burst,
  input   io_ps_axi_slave_aw_bits_lock,
  input  [3:0] io_ps_axi_slave_aw_bits_cache,
  input  [2:0] io_ps_axi_slave_aw_bits_prot,
  input  [3:0] io_ps_axi_slave_aw_bits_qos,
  input  [3:0] io_ps_axi_slave_aw_bits_region,
  input  [11:0] io_ps_axi_slave_aw_bits_id,
  input   io_ps_axi_slave_aw_bits_user,
  output  io_ps_axi_slave_w_ready,
  input   io_ps_axi_slave_w_valid,
  input  [31:0] io_ps_axi_slave_w_bits_data,
  input   io_ps_axi_slave_w_bits_last,
  input  [11:0] io_ps_axi_slave_w_bits_id,
  input  [3:0] io_ps_axi_slave_w_bits_strb,
  input   io_ps_axi_slave_w_bits_user,
  input   io_ps_axi_slave_b_ready,
  output  io_ps_axi_slave_b_valid,
  output [1:0] io_ps_axi_slave_b_bits_resp,
  output [11:0] io_ps_axi_slave_b_bits_id,
  output  io_ps_axi_slave_b_bits_user,
  output  io_ps_axi_slave_ar_ready,
  input   io_ps_axi_slave_ar_valid,
  input  [31:0] io_ps_axi_slave_ar_bits_addr,
  input  [7:0] io_ps_axi_slave_ar_bits_len,
  input  [2:0] io_ps_axi_slave_ar_bits_size,
  input  [1:0] io_ps_axi_slave_ar_bits_burst,
  input   io_ps_axi_slave_ar_bits_lock,
  input  [3:0] io_ps_axi_slave_ar_bits_cache,
  input  [2:0] io_ps_axi_slave_ar_bits_prot,
  input  [3:0] io_ps_axi_slave_ar_bits_qos,
  input  [3:0] io_ps_axi_slave_ar_bits_region,
  input  [11:0] io_ps_axi_slave_ar_bits_id,
  input   io_ps_axi_slave_ar_bits_user,
  input   io_ps_axi_slave_r_ready,
  output  io_ps_axi_slave_r_valid,
  output [1:0] io_ps_axi_slave_r_bits_resp,
  output [31:0] io_ps_axi_slave_r_bits_data,
  output  io_ps_axi_slave_r_bits_last,
  output [11:0] io_ps_axi_slave_r_bits_id,
  output  io_ps_axi_slave_r_bits_user,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user
);
  wire  adapter_clk;
  wire  adapter_reset;
  wire  adapter_io_nasti_aw_ready;
  wire  adapter_io_nasti_aw_valid;
  wire [31:0] adapter_io_nasti_aw_bits_addr;
  wire [7:0] adapter_io_nasti_aw_bits_len;
  wire [2:0] adapter_io_nasti_aw_bits_size;
  wire [1:0] adapter_io_nasti_aw_bits_burst;
  wire  adapter_io_nasti_aw_bits_lock;
  wire [3:0] adapter_io_nasti_aw_bits_cache;
  wire [2:0] adapter_io_nasti_aw_bits_prot;
  wire [3:0] adapter_io_nasti_aw_bits_qos;
  wire [3:0] adapter_io_nasti_aw_bits_region;
  wire [11:0] adapter_io_nasti_aw_bits_id;
  wire  adapter_io_nasti_aw_bits_user;
  wire  adapter_io_nasti_w_ready;
  wire  adapter_io_nasti_w_valid;
  wire [31:0] adapter_io_nasti_w_bits_data;
  wire  adapter_io_nasti_w_bits_last;
  wire [11:0] adapter_io_nasti_w_bits_id;
  wire [3:0] adapter_io_nasti_w_bits_strb;
  wire  adapter_io_nasti_w_bits_user;
  wire  adapter_io_nasti_b_ready;
  wire  adapter_io_nasti_b_valid;
  wire [1:0] adapter_io_nasti_b_bits_resp;
  wire [11:0] adapter_io_nasti_b_bits_id;
  wire  adapter_io_nasti_b_bits_user;
  wire  adapter_io_nasti_ar_ready;
  wire  adapter_io_nasti_ar_valid;
  wire [31:0] adapter_io_nasti_ar_bits_addr;
  wire [7:0] adapter_io_nasti_ar_bits_len;
  wire [2:0] adapter_io_nasti_ar_bits_size;
  wire [1:0] adapter_io_nasti_ar_bits_burst;
  wire  adapter_io_nasti_ar_bits_lock;
  wire [3:0] adapter_io_nasti_ar_bits_cache;
  wire [2:0] adapter_io_nasti_ar_bits_prot;
  wire [3:0] adapter_io_nasti_ar_bits_qos;
  wire [3:0] adapter_io_nasti_ar_bits_region;
  wire [11:0] adapter_io_nasti_ar_bits_id;
  wire  adapter_io_nasti_ar_bits_user;
  wire  adapter_io_nasti_r_ready;
  wire  adapter_io_nasti_r_valid;
  wire [1:0] adapter_io_nasti_r_bits_resp;
  wire [31:0] adapter_io_nasti_r_bits_data;
  wire  adapter_io_nasti_r_bits_last;
  wire [11:0] adapter_io_nasti_r_bits_id;
  wire  adapter_io_nasti_r_bits_user;
  wire  adapter_io_reset;
  wire  adapter_io_debug_req_ready;
  wire  adapter_io_debug_req_valid;
  wire [4:0] adapter_io_debug_req_bits_addr;
  wire [33:0] adapter_io_debug_req_bits_data;
  wire [1:0] adapter_io_debug_req_bits_op;
  wire  adapter_io_debug_resp_ready;
  wire  adapter_io_debug_resp_valid;
  wire [33:0] adapter_io_debug_resp_bits_data;
  wire [1:0] adapter_io_debug_resp_bits_resp;
  wire  rocket_clk;
  wire  rocket_reset;
  wire  rocket_io_mem_axi_0_aw_ready;
  wire  rocket_io_mem_axi_0_aw_valid;
  wire [31:0] rocket_io_mem_axi_0_aw_bits_addr;
  wire [7:0] rocket_io_mem_axi_0_aw_bits_len;
  wire [2:0] rocket_io_mem_axi_0_aw_bits_size;
  wire [1:0] rocket_io_mem_axi_0_aw_bits_burst;
  wire  rocket_io_mem_axi_0_aw_bits_lock;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_cache;
  wire [2:0] rocket_io_mem_axi_0_aw_bits_prot;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_qos;
  wire [3:0] rocket_io_mem_axi_0_aw_bits_region;
  wire [4:0] rocket_io_mem_axi_0_aw_bits_id;
  wire  rocket_io_mem_axi_0_aw_bits_user;
  wire  rocket_io_mem_axi_0_w_ready;
  wire  rocket_io_mem_axi_0_w_valid;
  wire [63:0] rocket_io_mem_axi_0_w_bits_data;
  wire  rocket_io_mem_axi_0_w_bits_last;
  wire [4:0] rocket_io_mem_axi_0_w_bits_id;
  wire [7:0] rocket_io_mem_axi_0_w_bits_strb;
  wire  rocket_io_mem_axi_0_w_bits_user;
  wire  rocket_io_mem_axi_0_b_ready;
  wire  rocket_io_mem_axi_0_b_valid;
  wire [1:0] rocket_io_mem_axi_0_b_bits_resp;
  wire [4:0] rocket_io_mem_axi_0_b_bits_id;
  wire  rocket_io_mem_axi_0_b_bits_user;
  wire  rocket_io_mem_axi_0_ar_ready;
  wire  rocket_io_mem_axi_0_ar_valid;
  wire [31:0] rocket_io_mem_axi_0_ar_bits_addr;
  wire [7:0] rocket_io_mem_axi_0_ar_bits_len;
  wire [2:0] rocket_io_mem_axi_0_ar_bits_size;
  wire [1:0] rocket_io_mem_axi_0_ar_bits_burst;
  wire  rocket_io_mem_axi_0_ar_bits_lock;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_cache;
  wire [2:0] rocket_io_mem_axi_0_ar_bits_prot;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_qos;
  wire [3:0] rocket_io_mem_axi_0_ar_bits_region;
  wire [4:0] rocket_io_mem_axi_0_ar_bits_id;
  wire  rocket_io_mem_axi_0_ar_bits_user;
  wire  rocket_io_mem_axi_0_r_ready;
  wire  rocket_io_mem_axi_0_r_valid;
  wire [1:0] rocket_io_mem_axi_0_r_bits_resp;
  wire [63:0] rocket_io_mem_axi_0_r_bits_data;
  wire  rocket_io_mem_axi_0_r_bits_last;
  wire [4:0] rocket_io_mem_axi_0_r_bits_id;
  wire  rocket_io_mem_axi_0_r_bits_user;
  wire  rocket_io_interrupts_0;
  wire  rocket_io_interrupts_1;
  wire  rocket_io_debug_req_ready;
  wire  rocket_io_debug_req_valid;
  wire [4:0] rocket_io_debug_req_bits_addr;
  wire [33:0] rocket_io_debug_req_bits_data;
  wire [1:0] rocket_io_debug_req_bits_op;
  wire  rocket_io_debug_resp_ready;
  wire  rocket_io_debug_resp_valid;
  wire [33:0] rocket_io_debug_resp_bits_data;
  wire [1:0] rocket_io_debug_resp_bits_resp;
  ZynqAdapter adapter (
    .clk(adapter_clk),
    .reset(adapter_reset),
    .io_nasti_aw_ready(adapter_io_nasti_aw_ready),
    .io_nasti_aw_valid(adapter_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(adapter_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(adapter_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(adapter_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(adapter_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(adapter_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(adapter_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(adapter_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(adapter_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(adapter_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(adapter_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(adapter_io_nasti_aw_bits_user),
    .io_nasti_w_ready(adapter_io_nasti_w_ready),
    .io_nasti_w_valid(adapter_io_nasti_w_valid),
    .io_nasti_w_bits_data(adapter_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(adapter_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(adapter_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(adapter_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(adapter_io_nasti_w_bits_user),
    .io_nasti_b_ready(adapter_io_nasti_b_ready),
    .io_nasti_b_valid(adapter_io_nasti_b_valid),
    .io_nasti_b_bits_resp(adapter_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(adapter_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(adapter_io_nasti_b_bits_user),
    .io_nasti_ar_ready(adapter_io_nasti_ar_ready),
    .io_nasti_ar_valid(adapter_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(adapter_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(adapter_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(adapter_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(adapter_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(adapter_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(adapter_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(adapter_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(adapter_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(adapter_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(adapter_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(adapter_io_nasti_ar_bits_user),
    .io_nasti_r_ready(adapter_io_nasti_r_ready),
    .io_nasti_r_valid(adapter_io_nasti_r_valid),
    .io_nasti_r_bits_resp(adapter_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(adapter_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(adapter_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(adapter_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(adapter_io_nasti_r_bits_user),
    .io_reset(adapter_io_reset),
    .io_debug_req_ready(adapter_io_debug_req_ready),
    .io_debug_req_valid(adapter_io_debug_req_valid),
    .io_debug_req_bits_addr(adapter_io_debug_req_bits_addr),
    .io_debug_req_bits_data(adapter_io_debug_req_bits_data),
    .io_debug_req_bits_op(adapter_io_debug_req_bits_op),
    .io_debug_resp_ready(adapter_io_debug_resp_ready),
    .io_debug_resp_valid(adapter_io_debug_resp_valid),
    .io_debug_resp_bits_data(adapter_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(adapter_io_debug_resp_bits_resp)
  );
  Top_1 rocket (
    .clk(rocket_clk),
    .reset(rocket_reset),
    .io_mem_axi_0_aw_ready(rocket_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(rocket_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(rocket_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(rocket_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(rocket_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(rocket_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(rocket_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(rocket_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(rocket_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(rocket_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(rocket_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(rocket_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(rocket_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(rocket_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(rocket_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(rocket_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(rocket_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(rocket_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(rocket_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(rocket_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(rocket_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(rocket_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(rocket_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(rocket_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(rocket_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(rocket_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(rocket_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(rocket_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(rocket_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(rocket_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(rocket_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(rocket_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(rocket_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(rocket_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(rocket_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(rocket_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(rocket_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(rocket_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(rocket_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(rocket_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(rocket_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(rocket_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(rocket_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(rocket_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(rocket_io_mem_axi_0_r_bits_user),
    .io_interrupts_0(rocket_io_interrupts_0),
    .io_interrupts_1(rocket_io_interrupts_1),
    .io_debug_req_ready(rocket_io_debug_req_ready),
    .io_debug_req_valid(rocket_io_debug_req_valid),
    .io_debug_req_bits_addr(rocket_io_debug_req_bits_addr),
    .io_debug_req_bits_data(rocket_io_debug_req_bits_data),
    .io_debug_req_bits_op(rocket_io_debug_req_bits_op),
    .io_debug_resp_ready(rocket_io_debug_resp_ready),
    .io_debug_resp_valid(rocket_io_debug_resp_valid),
    .io_debug_resp_bits_data(rocket_io_debug_resp_bits_data),
    .io_debug_resp_bits_resp(rocket_io_debug_resp_bits_resp)
  );
  assign io_ps_axi_slave_aw_ready = adapter_io_nasti_aw_ready;
  assign io_ps_axi_slave_w_ready = adapter_io_nasti_w_ready;
  assign io_ps_axi_slave_b_valid = adapter_io_nasti_b_valid;
  assign io_ps_axi_slave_b_bits_resp = adapter_io_nasti_b_bits_resp;
  assign io_ps_axi_slave_b_bits_id = adapter_io_nasti_b_bits_id;
  assign io_ps_axi_slave_b_bits_user = adapter_io_nasti_b_bits_user;
  assign io_ps_axi_slave_ar_ready = adapter_io_nasti_ar_ready;
  assign io_ps_axi_slave_r_valid = adapter_io_nasti_r_valid;
  assign io_ps_axi_slave_r_bits_resp = adapter_io_nasti_r_bits_resp;
  assign io_ps_axi_slave_r_bits_data = adapter_io_nasti_r_bits_data;
  assign io_ps_axi_slave_r_bits_last = adapter_io_nasti_r_bits_last;
  assign io_ps_axi_slave_r_bits_id = adapter_io_nasti_r_bits_id;
  assign io_ps_axi_slave_r_bits_user = adapter_io_nasti_r_bits_user;
  assign io_mem_axi_0_aw_valid = rocket_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = rocket_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = rocket_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = rocket_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = rocket_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = rocket_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = rocket_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = rocket_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = rocket_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = rocket_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = rocket_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = rocket_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = rocket_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = rocket_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = rocket_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = rocket_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = rocket_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = rocket_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = rocket_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = rocket_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = rocket_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = rocket_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = rocket_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = rocket_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = rocket_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = rocket_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = rocket_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = rocket_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = rocket_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = rocket_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = rocket_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = rocket_io_mem_axi_0_r_ready;
  assign adapter_clk = clk;
  assign adapter_reset = reset;
  assign adapter_io_nasti_aw_valid = io_ps_axi_slave_aw_valid;
  assign adapter_io_nasti_aw_bits_addr = io_ps_axi_slave_aw_bits_addr;
  assign adapter_io_nasti_aw_bits_len = io_ps_axi_slave_aw_bits_len;
  assign adapter_io_nasti_aw_bits_size = io_ps_axi_slave_aw_bits_size;
  assign adapter_io_nasti_aw_bits_burst = io_ps_axi_slave_aw_bits_burst;
  assign adapter_io_nasti_aw_bits_lock = io_ps_axi_slave_aw_bits_lock;
  assign adapter_io_nasti_aw_bits_cache = io_ps_axi_slave_aw_bits_cache;
  assign adapter_io_nasti_aw_bits_prot = io_ps_axi_slave_aw_bits_prot;
  assign adapter_io_nasti_aw_bits_qos = io_ps_axi_slave_aw_bits_qos;
  assign adapter_io_nasti_aw_bits_region = io_ps_axi_slave_aw_bits_region;
  assign adapter_io_nasti_aw_bits_id = io_ps_axi_slave_aw_bits_id;
  assign adapter_io_nasti_aw_bits_user = io_ps_axi_slave_aw_bits_user;
  assign adapter_io_nasti_w_valid = io_ps_axi_slave_w_valid;
  assign adapter_io_nasti_w_bits_data = io_ps_axi_slave_w_bits_data;
  assign adapter_io_nasti_w_bits_last = io_ps_axi_slave_w_bits_last;
  assign adapter_io_nasti_w_bits_id = io_ps_axi_slave_w_bits_id;
  assign adapter_io_nasti_w_bits_strb = io_ps_axi_slave_w_bits_strb;
  assign adapter_io_nasti_w_bits_user = io_ps_axi_slave_w_bits_user;
  assign adapter_io_nasti_b_ready = io_ps_axi_slave_b_ready;
  assign adapter_io_nasti_ar_valid = io_ps_axi_slave_ar_valid;
  assign adapter_io_nasti_ar_bits_addr = io_ps_axi_slave_ar_bits_addr;
  assign adapter_io_nasti_ar_bits_len = io_ps_axi_slave_ar_bits_len;
  assign adapter_io_nasti_ar_bits_size = io_ps_axi_slave_ar_bits_size;
  assign adapter_io_nasti_ar_bits_burst = io_ps_axi_slave_ar_bits_burst;
  assign adapter_io_nasti_ar_bits_lock = io_ps_axi_slave_ar_bits_lock;
  assign adapter_io_nasti_ar_bits_cache = io_ps_axi_slave_ar_bits_cache;
  assign adapter_io_nasti_ar_bits_prot = io_ps_axi_slave_ar_bits_prot;
  assign adapter_io_nasti_ar_bits_qos = io_ps_axi_slave_ar_bits_qos;
  assign adapter_io_nasti_ar_bits_region = io_ps_axi_slave_ar_bits_region;
  assign adapter_io_nasti_ar_bits_id = io_ps_axi_slave_ar_bits_id;
  assign adapter_io_nasti_ar_bits_user = io_ps_axi_slave_ar_bits_user;
  assign adapter_io_nasti_r_ready = io_ps_axi_slave_r_ready;
  assign adapter_io_debug_req_ready = rocket_io_debug_req_ready;
  assign adapter_io_debug_resp_valid = rocket_io_debug_resp_valid;
  assign adapter_io_debug_resp_bits_data = rocket_io_debug_resp_bits_data;
  assign adapter_io_debug_resp_bits_resp = rocket_io_debug_resp_bits_resp;
  assign rocket_clk = clk;
  assign rocket_reset = adapter_io_reset;
  assign rocket_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign rocket_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign rocket_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign rocket_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign rocket_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign rocket_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign rocket_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign rocket_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign rocket_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign rocket_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign rocket_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign rocket_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign rocket_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign rocket_io_interrupts_0 = 1'h0;
  assign rocket_io_interrupts_1 = 1'h0;
  assign rocket_io_debug_req_valid = adapter_io_debug_req_valid;
  assign rocket_io_debug_req_bits_addr = adapter_io_debug_req_bits_addr;
  assign rocket_io_debug_req_bits_data = adapter_io_debug_req_bits_data;
  assign rocket_io_debug_req_bits_op = adapter_io_debug_req_bits_op;
  assign rocket_io_debug_resp_ready = adapter_io_debug_resp_ready;
endmodule
