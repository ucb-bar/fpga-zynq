module BTB(input clk, input reset,
    input [42:0] io_req,
    output io_resp_valid,
    output io_resp_bits_taken,
    output[42:0] io_resp_bits_target,
    output[2:0] io_resp_bits_entry,
    output[3:0] io_resp_bits_bht_index,
    output[1:0] io_resp_bits_bht_value,
    input  io_update_valid,
    input  io_update_bits_prediction_valid,
    input  io_update_bits_prediction_bits_taken,
    input [42:0] io_update_bits_prediction_bits_target,
    input [2:0] io_update_bits_prediction_bits_entry,
    input [3:0] io_update_bits_prediction_bits_bht_index,
    input [1:0] io_update_bits_prediction_bits_bht_value,
    input [42:0] io_update_bits_pc,
    input [42:0] io_update_bits_target,
    input [42:0] io_update_bits_returnAddr,
    input  io_update_bits_taken,
    input  io_update_bits_isJump,
    input  io_update_bits_isCall,
    input  io_update_bits_isReturn,
    input  io_update_bits_incorrectTarget,
    input  io_invalidate
);

  reg[0:0] T0 = 1'b0;
  wire T1;
  wire T2;
  wire T3;
  reg [42:0] R4;
  wire[42:0] T5;
  wire T6;
  wire T7;
  wire updateTarget;
  reg  R8;
  wire T9;
  wire updateValid;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  reg  R16;
  wire T17;
  wire[1:0] T18;
  wire[1:0] T19;
  reg [1:0] T20 [15:0];
  wire[1:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  reg  R25;
  wire T26;
  wire T27;
  wire T28;
  reg [1:0] R29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  R37;
  wire T38;
  wire T39;
  reg [3:0] R40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  reg [3:0] R44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire[2:0] T47;
  wire[3:0] T48;
  wire[2:0] T49;
  wire[1:0] T50;
  wire T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire[3:0] T54;
  wire[3:0] T55;
  wire[7:0] hits;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[3:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[3:0] T61;
  wire[3:0] pageHit;
  reg [3:0] pageValid;
  wire[3:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] pageReplEn;
  wire[3:0] tgtPageReplEn;
  wire[3:0] tgtPageRepl;
  wire[3:0] T66;
  wire[3:0] T67;
  wire T68;
  wire[3:0] idxPageUpdateOH;
  wire[3:0] idxPageRepl;
  wire[3:0] T69;
  reg [1:0] R70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire doPageRepl;
  wire doTgtPageRepl;
  wire T75;
  wire T76;
  wire[3:0] T77;
  wire[3:0] T78;
  wire[3:0] idxPageReplEn;
  wire doIdxPageRepl;
  wire T79;
  wire T80;
  wire[3:0] updatePageHit;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[1:0] T83;
  wire T84;
  wire[29:0] T85;
  reg [42:0] R86;
  wire[42:0] T87;
  wire[29:0] T88;
  reg [29:0] pages [3:0];
  wire[29:0] T89;
  wire[29:0] T90;
  wire[29:0] T91;
  wire[29:0] T92;
  wire T93;
  wire[3:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[29:0] T99;
  wire T100;
  wire T101;
  wire T102;
  wire[29:0] T103;
  wire[29:0] T104;
  wire[29:0] T105;
  wire[29:0] T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[29:0] T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[29:0] T116;
  wire[1:0] T117;
  wire T118;
  wire[29:0] T119;
  wire T120;
  wire[29:0] T121;
  wire T122;
  wire T123;
  wire samePage;
  wire[29:0] T124;
  wire[29:0] T125;
  wire[3:0] T126;
  wire[2:0] T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[1:0] T131;
  wire T132;
  wire[29:0] T133;
  wire[29:0] T134;
  wire T135;
  wire[29:0] T136;
  wire[1:0] T137;
  wire T138;
  wire[29:0] T139;
  wire T140;
  wire[29:0] T141;
  wire[3:0] T142;
  wire[3:0] T143;
  wire[1:0] T144;
  reg [1:0] idxPages [7:0];
  wire[1:0] T145;
  wire[1:0] T146;
  wire T147;
  wire[1:0] T148;
  wire[1:0] T149;
  wire[1:0] T150;
  wire T151;
  wire[2:0] T152;
  reg [2:0] R153;
  wire[2:0] T154;
  wire[2:0] T155;
  wire[2:0] T156;
  wire T157;
  wire T158;
  wire T159;
  reg [2:0] R160;
  wire[2:0] T161;
  wire T162;
  wire[3:0] T163;
  wire[3:0] T164;
  wire[3:0] T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire[1:0] T172;
  wire T173;
  wire[3:0] T174;
  wire[3:0] T175;
  wire[3:0] T176;
  wire[1:0] T177;
  wire[3:0] T178;
  wire[1:0] T179;
  wire T180;
  wire[3:0] T181;
  wire[3:0] T182;
  wire[3:0] T183;
  wire[1:0] T184;
  wire T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[3:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[1:0] T195;
  wire T196;
  wire[3:0] T197;
  wire[3:0] T198;
  wire[3:0] T199;
  wire[1:0] T200;
  wire[7:0] T201;
  wire[7:0] T202;
  wire[7:0] T203;
  wire[3:0] T204;
  wire[1:0] T205;
  wire T206;
  wire[12:0] T207;
  wire[12:0] T208;
  reg [12:0] idxs [7:0];
  wire[12:0] T209;
  wire[12:0] T210;
  wire T211;
  wire[12:0] T212;
  wire[1:0] T213;
  wire T214;
  wire[12:0] T215;
  wire T216;
  wire[12:0] T217;
  wire[3:0] T218;
  wire[1:0] T219;
  wire T220;
  wire[12:0] T221;
  wire T222;
  wire[12:0] T223;
  wire[1:0] T224;
  wire T225;
  wire[12:0] T226;
  wire T227;
  wire[12:0] T228;
  reg [7:0] idxValid;
  wire[7:0] T229;
  wire[7:0] T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire[7:0] T234;
  wire[7:0] T235;
  wire[7:0] T236;
  wire[3:0] T237;
  wire[1:0] T238;
  wire T239;
  wire[3:0] T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[1:0] T244;
  reg [1:0] tgtPages [7:0];
  wire[1:0] T245;
  wire[1:0] T246;
  wire T247;
  wire[1:0] T248;
  wire[1:0] T249;
  wire[3:0] T250;
  wire[1:0] T251;
  wire T252;
  wire T253;
  wire[3:0] T254;
  wire[3:0] T255;
  wire[3:0] T256;
  wire[3:0] T257;
  wire[1:0] T258;
  wire[1:0] T259;
  wire T260;
  wire[3:0] T261;
  wire[3:0] T262;
  wire[3:0] T263;
  wire[3:0] T264;
  wire[1:0] T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[3:0] T270;
  wire[1:0] T271;
  wire[3:0] T272;
  wire[1:0] T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[3:0] T278;
  wire[1:0] T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[1:0] T285;
  wire[1:0] T286;
  wire T287;
  wire[3:0] T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[1:0] T292;
  wire T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[3:0] T296;
  wire[3:0] T297;
  wire[1:0] T298;
  wire[7:0] T299;
  wire[7:0] T300;
  wire[7:0] T301;
  wire[7:0] T302;
  wire[7:0] T303;
  wire[7:0] T304;
  wire T305;
  wire T306;
  wire[7:0] T307;
  wire[7:0] T308;
  wire[3:0] T309;
  wire[1:0] T310;
  wire T311;
  wire T312;
  wire[42:0] T313;
  wire[42:0] T314;
  wire[42:0] T315;
  wire[12:0] T316;
  wire[12:0] T317;
  wire[12:0] T318;
  reg [12:0] tgts [7:0];
  wire[12:0] T319;
  wire[12:0] T320;
  wire T321;
  wire[12:0] T322;
  wire[12:0] T323;
  wire[12:0] T324;
  wire T325;
  wire[12:0] T326;
  wire[12:0] T327;
  wire[12:0] T328;
  wire T329;
  wire[12:0] T330;
  wire[12:0] T331;
  wire[12:0] T332;
  wire T333;
  wire[12:0] T334;
  wire[12:0] T335;
  wire[12:0] T336;
  wire T337;
  wire[12:0] T338;
  wire[12:0] T339;
  wire[12:0] T340;
  wire T341;
  wire[12:0] T342;
  wire[12:0] T343;
  wire[12:0] T344;
  wire T345;
  wire[12:0] T346;
  wire[12:0] T347;
  wire T348;
  wire[29:0] T349;
  wire[29:0] T350;
  wire[29:0] T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire T358;
  wire[3:0] T359;
  wire[3:0] T360;
  wire T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire T364;
  wire[3:0] T365;
  wire[3:0] T366;
  wire T367;
  wire[3:0] T368;
  wire[3:0] T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire T373;
  wire[3:0] T374;
  wire T375;
  wire[29:0] T376;
  wire[29:0] T377;
  wire[29:0] T378;
  wire T379;
  wire[29:0] T380;
  wire[29:0] T381;
  wire[29:0] T382;
  wire T383;
  wire[29:0] T384;
  wire[29:0] T385;
  wire T386;
  wire[42:0] T387;
  reg [42:0] R388;
  wire[42:0] T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire T393;
  wire T394;
  reg  R395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  reg [1:0] R404;
  wire[1:0] T405;
  wire[1:0] T406;
  wire[1:0] T407;
  wire[1:0] T408;
  wire[1:0] T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  reg [42:0] R417;
  wire[42:0] T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[7:0] T424;
  reg [7:0] useRAS;
  wire[7:0] T425;
  wire[7:0] T426;
  wire[7:0] T427;
  wire[7:0] T428;
  wire[7:0] T429;
  wire[7:0] T430;
  wire[7:0] T431;
  wire T432;
  wire T433;
  reg  R434;
  wire T435;
  wire[7:0] T436;
  wire[7:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire[7:0] T445;
  reg [7:0] isJump;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T448;
  wire[7:0] T449;
  wire[7:0] T450;
  wire[7:0] T451;
  wire[7:0] T452;
  wire T453;
  wire T454;
  wire[7:0] T455;
  wire[7:0] T456;
  wire T457;
  wire T458;
  wire T459;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R4 = {2{$random}};
    R8 = {1{$random}};
    R10 = {1{$random}};
    R16 = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      T20[initvar] = {1{$random}};
    R25 = {1{$random}};
    R29 = {1{$random}};
    R37 = {1{$random}};
    R40 = {1{$random}};
    R44 = {1{$random}};
    pageValid = {1{$random}};
    R70 = {1{$random}};
    R86 = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      pages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxPages[initvar] = {1{$random}};
    R153 = {1{$random}};
    R160 = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      idxs[initvar] = {1{$random}};
    idxValid = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgtPages[initvar] = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      tgts[initvar] = {1{$random}};
    R388 = {2{$random}};
    R395 = {1{$random}};
    R404 = {1{$random}};
    R417 = {2{$random}};
    useRAS = {1{$random}};
    R434 = {1{$random}};
    isJump = {1{$random}};
  end
`endif

  assign T1 = T2 | reset;
  assign T2 = T6 | T3;
  assign T3 = io_req == R4;
  assign T5 = io_update_valid ? io_update_bits_target : R4;
  assign T6 = T7 ^ 1'h1;
  assign T7 = T12 & updateTarget;
  assign updateTarget = updateValid & R8;
  assign T9 = io_update_valid ? io_update_bits_incorrectTarget : R8;
  assign updateValid = R8 | R10;
  assign T11 = io_update_valid ? io_update_bits_prediction_valid : R10;
  assign T12 = R16 & T13;
  assign T13 = T14 ^ 1'h1;
  assign T14 = updateValid & T15;
  assign T15 = updateTarget ^ 1'h1;
  assign T17 = reset ? 1'h0 : io_update_valid;
  assign io_resp_bits_bht_value = T18;
  assign T18 = T19;
  assign T19 = T20[T42];
  assign T22 = {R25, T23};
  assign T23 = T32 | T24;
  assign T24 = T27 & R25;
  assign T26 = io_update_valid ? io_update_bits_taken : R25;
  assign T27 = T31 | T28;
  assign T28 = R29[1'h0:1'h0];
  assign T30 = io_update_valid ? io_update_bits_prediction_bits_bht_value : R29;
  assign T31 = R29[1'h1:1'h1];
  assign T32 = T34 & T33;
  assign T33 = R29[1'h0:1'h0];
  assign T34 = R29[1'h1:1'h1];
  assign T35 = T39 & T36;
  assign T36 = R37 ^ 1'h1;
  assign T38 = io_update_valid ? io_update_bits_isJump : R37;
  assign T39 = R16 & R10;
  assign T41 = io_update_valid ? io_update_bits_prediction_bits_bht_index : R40;
  assign T42 = T43;
  assign T43 = T48 ^ R44;
  assign T45 = T35 ? T46 : R44;
  assign T46 = {R25, T47};
  assign T47 = R44[2'h3:1'h1];
  assign T48 = io_req[3'h5:2'h2];
  assign io_resp_bits_bht_index = T42;
  assign io_resp_bits_entry = T49;
  assign T49 = {T312, T50};
  assign T50 = {T311, T51};
  assign T51 = T52[1'h1:1'h1];
  assign T52 = T310 | T53;
  assign T53 = T54[1'h1:1'h0];
  assign T54 = T309 | T55;
  assign T55 = hits[2'h3:1'h0];
  assign hits = T201 & T56;
  assign T56 = T57;
  assign T57 = {T178, T58};
  assign T58 = {T167, T59};
  assign T59 = {T162, T60};
  assign T60 = T61 != 4'h0;
  assign T61 = T142 & pageHit;
  assign pageHit = T129 & pageValid;
  assign T62 = reset ? 4'h0 : T63;
  assign T63 = io_invalidate ? 4'h0 : T64;
  assign T64 = T128 ? T65 : pageValid;
  assign T65 = pageValid | pageReplEn;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : 4'h0;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T66;
  assign T66 = T126 | T67;
  assign T67 = {3'h0, T68};
  assign T68 = idxPageUpdateOH[2'h3:2'h3];
  assign idxPageUpdateOH = T80 ? updatePageHit : idxPageRepl;
  assign idxPageRepl = T69;
  assign T69 = 1'h1 << R70;
  assign T71 = reset ? 2'h0 : T72;
  assign T72 = T74 ? T73 : R70;
  assign T73 = R70 + 2'h1;
  assign T74 = R16 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doTgtPageRepl = T122 & T75;
  assign T75 = T76 ^ 1'h1;
  assign T76 = T77 != 4'h0;
  assign T77 = pageHit & T78;
  assign T78 = ~ idxPageReplEn;
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : 4'h0;
  assign doIdxPageRepl = updateTarget & T79;
  assign T79 = T80 ^ 1'h1;
  assign T80 = updatePageHit != 4'h0;
  assign updatePageHit = T81 & pageValid;
  assign T81 = T82;
  assign T82 = {T117, T83};
  assign T83 = {T115, T84};
  assign T84 = T88 == T85;
  assign T85 = R86 >> 4'hd;
  assign T87 = io_update_valid ? io_update_bits_pc : R86;
  assign T88 = pages[2'h0];
  assign T90 = T93 ? T92 : T91;
  assign T91 = R86 >> 4'hd;
  assign T92 = io_req >> 4'hd;
  assign T93 = T94 != 4'h0;
  assign T94 = idxPageUpdateOH & 4'h5;
  assign T95 = T12 & T96;
  assign T96 = T98 & T97;
  assign T97 = pageReplEn[2'h3:2'h3];
  assign T98 = T93 ? doTgtPageRepl : doIdxPageRepl;
  assign T100 = T12 & T101;
  assign T101 = T98 & T102;
  assign T102 = pageReplEn[1'h1:1'h1];
  assign T104 = T93 ? T106 : T105;
  assign T105 = io_req >> 4'hd;
  assign T106 = R86 >> 4'hd;
  assign T107 = T12 & T108;
  assign T108 = T110 & T109;
  assign T109 = pageReplEn[2'h2:2'h2];
  assign T110 = T93 ? doIdxPageRepl : doTgtPageRepl;
  assign T112 = T12 & T113;
  assign T113 = T110 & T114;
  assign T114 = pageReplEn[1'h0:1'h0];
  assign T115 = T116 == T85;
  assign T116 = pages[2'h1];
  assign T117 = {T120, T118};
  assign T118 = T119 == T85;
  assign T119 = pages[2'h2];
  assign T120 = T121 == T85;
  assign T121 = pages[2'h3];
  assign T122 = updateTarget & T123;
  assign T123 = samePage ^ 1'h1;
  assign samePage = T125 == T124;
  assign T124 = io_req >> 4'hd;
  assign T125 = R86 >> 4'hd;
  assign T126 = T127 << 1'h1;
  assign T127 = idxPageUpdateOH[2'h2:1'h0];
  assign T128 = T12 & doPageRepl;
  assign T129 = T130;
  assign T130 = {T137, T131};
  assign T131 = {T135, T132};
  assign T132 = T134 == T133;
  assign T133 = io_req >> 4'hd;
  assign T134 = pages[2'h0];
  assign T135 = T136 == T133;
  assign T136 = pages[2'h1];
  assign T137 = {T140, T138};
  assign T138 = T139 == T133;
  assign T139 = pages[2'h2];
  assign T140 = T141 == T133;
  assign T141 = pages[2'h3];
  assign T142 = T143[2'h3:1'h0];
  assign T143 = 1'h1 << T144;
  assign T144 = idxPages[3'h0];
  assign T146 = {T151, T147};
  assign T147 = T148[1'h1:1'h1];
  assign T148 = T150 | T149;
  assign T149 = idxPageUpdateOH[1'h1:1'h0];
  assign T150 = idxPageUpdateOH[2'h3:2'h2];
  assign T151 = T150 != 2'h0;
  assign T152 = R10 ? R160 : R153;
  assign T154 = reset ? 3'h0 : T155;
  assign T155 = T157 ? T156 : R153;
  assign T156 = R153 + 3'h1;
  assign T157 = T12 & T158;
  assign T158 = T159 & updateValid;
  assign T159 = R10 ^ 1'h1;
  assign T161 = io_update_valid ? io_update_bits_prediction_bits_entry : R160;
  assign T162 = T163 != 4'h0;
  assign T163 = T164 & pageHit;
  assign T164 = T165[2'h3:1'h0];
  assign T165 = 1'h1 << T166;
  assign T166 = idxPages[3'h1];
  assign T167 = {T173, T168};
  assign T168 = T169 != 4'h0;
  assign T169 = T170 & pageHit;
  assign T170 = T171[2'h3:1'h0];
  assign T171 = 1'h1 << T172;
  assign T172 = idxPages[3'h2];
  assign T173 = T174 != 4'h0;
  assign T174 = T175 & pageHit;
  assign T175 = T176[2'h3:1'h0];
  assign T176 = 1'h1 << T177;
  assign T177 = idxPages[3'h3];
  assign T178 = {T190, T179};
  assign T179 = {T185, T180};
  assign T180 = T181 != 4'h0;
  assign T181 = T182 & pageHit;
  assign T182 = T183[2'h3:1'h0];
  assign T183 = 1'h1 << T184;
  assign T184 = idxPages[3'h4];
  assign T185 = T186 != 4'h0;
  assign T186 = T187 & pageHit;
  assign T187 = T188[2'h3:1'h0];
  assign T188 = 1'h1 << T189;
  assign T189 = idxPages[3'h5];
  assign T190 = {T196, T191};
  assign T191 = T192 != 4'h0;
  assign T192 = T193 & pageHit;
  assign T193 = T194[2'h3:1'h0];
  assign T194 = 1'h1 << T195;
  assign T195 = idxPages[3'h6];
  assign T196 = T197 != 4'h0;
  assign T197 = T198 & pageHit;
  assign T198 = T199[2'h3:1'h0];
  assign T199 = 1'h1 << T200;
  assign T200 = idxPages[3'h7];
  assign T201 = idxValid & T202;
  assign T202 = T203;
  assign T203 = {T218, T204};
  assign T204 = {T213, T205};
  assign T205 = {T211, T206};
  assign T206 = T208 == T207;
  assign T207 = io_req[4'hc:1'h0];
  assign T208 = idxs[3'h0];
  assign T210 = R86[4'hc:1'h0];
  assign T211 = T212 == T207;
  assign T212 = idxs[3'h1];
  assign T213 = {T216, T214};
  assign T214 = T215 == T207;
  assign T215 = idxs[3'h2];
  assign T216 = T217 == T207;
  assign T217 = idxs[3'h3];
  assign T218 = {T224, T219};
  assign T219 = {T222, T220};
  assign T220 = T221 == T207;
  assign T221 = idxs[3'h4];
  assign T222 = T223 == T207;
  assign T223 = idxs[3'h5];
  assign T224 = {T227, T225};
  assign T225 = T226 == T207;
  assign T226 = idxs[3'h6];
  assign T227 = T228 == T207;
  assign T228 = idxs[3'h7];
  assign T229 = reset ? 8'h0 : T230;
  assign T230 = io_invalidate ? 8'h0 : T231;
  assign T231 = T12 ? T299 : T232;
  assign T232 = T12 ? T233 : idxValid;
  assign T233 = idxValid & T234;
  assign T234 = ~ T235;
  assign T235 = T236;
  assign T236 = {T272, T237};
  assign T237 = {T259, T238};
  assign T238 = {T253, T239};
  assign T239 = T240 != 4'h0;
  assign T240 = pageReplEn & T241;
  assign T241 = T142 | T242;
  assign T242 = T243[2'h3:1'h0];
  assign T243 = 1'h1 << T244;
  assign T244 = tgtPages[3'h0];
  assign T246 = {T252, T247};
  assign T247 = T248[1'h1:1'h1];
  assign T248 = T251 | T249;
  assign T249 = T250[1'h1:1'h0];
  assign T250 = T76 ? pageHit : tgtPageRepl;
  assign T251 = T250[2'h3:2'h2];
  assign T252 = T251 != 2'h0;
  assign T253 = T254 != 4'h0;
  assign T254 = pageReplEn & T255;
  assign T255 = T164 | T256;
  assign T256 = T257[2'h3:1'h0];
  assign T257 = 1'h1 << T258;
  assign T258 = tgtPages[3'h1];
  assign T259 = {T266, T260};
  assign T260 = T261 != 4'h0;
  assign T261 = pageReplEn & T262;
  assign T262 = T170 | T263;
  assign T263 = T264[2'h3:1'h0];
  assign T264 = 1'h1 << T265;
  assign T265 = tgtPages[3'h2];
  assign T266 = T267 != 4'h0;
  assign T267 = pageReplEn & T268;
  assign T268 = T175 | T269;
  assign T269 = T270[2'h3:1'h0];
  assign T270 = 1'h1 << T271;
  assign T271 = tgtPages[3'h3];
  assign T272 = {T286, T273};
  assign T273 = {T280, T274};
  assign T274 = T275 != 4'h0;
  assign T275 = pageReplEn & T276;
  assign T276 = T182 | T277;
  assign T277 = T278[2'h3:1'h0];
  assign T278 = 1'h1 << T279;
  assign T279 = tgtPages[3'h4];
  assign T280 = T281 != 4'h0;
  assign T281 = pageReplEn & T282;
  assign T282 = T187 | T283;
  assign T283 = T284[2'h3:1'h0];
  assign T284 = 1'h1 << T285;
  assign T285 = tgtPages[3'h5];
  assign T286 = {T293, T287};
  assign T287 = T288 != 4'h0;
  assign T288 = pageReplEn & T289;
  assign T289 = T193 | T290;
  assign T290 = T291[2'h3:1'h0];
  assign T291 = 1'h1 << T292;
  assign T292 = tgtPages[3'h6];
  assign T293 = T294 != 4'h0;
  assign T294 = pageReplEn & T295;
  assign T295 = T198 | T296;
  assign T296 = T297[2'h3:1'h0];
  assign T297 = 1'h1 << T298;
  assign T298 = tgtPages[3'h7];
  assign T299 = T307 | T300;
  assign T300 = T304 & T301;
  assign T301 = T303 | T302;
  assign T302 = idxValid ^ idxValid;
  assign T303 = 1'h1 << T152;
  assign T304 = T305 ? 8'hff : 8'h0;
  assign T305 = T306;
  assign T306 = updateValid;
  assign T307 = T232 & T308;
  assign T308 = ~ T301;
  assign T309 = hits[3'h7:3'h4];
  assign T310 = T54[2'h3:2'h2];
  assign T311 = T310 != 2'h0;
  assign T312 = T309 != 4'h0;
  assign io_resp_bits_target = T313;
  assign T313 = T440 ? io_update_bits_returnAddr : T314;
  assign T314 = T422 ? T387 : T315;
  assign T315 = {T349, T316};
  assign T316 = T322 | T317;
  assign T317 = T321 ? T318 : 13'h0;
  assign T318 = tgts[3'h7];
  assign T320 = io_req[4'hc:1'h0];
  assign T321 = hits[3'h7:3'h7];
  assign T322 = T326 | T323;
  assign T323 = T325 ? T324 : 13'h0;
  assign T324 = tgts[3'h6];
  assign T325 = hits[3'h6:3'h6];
  assign T326 = T330 | T327;
  assign T327 = T329 ? T328 : 13'h0;
  assign T328 = tgts[3'h5];
  assign T329 = hits[3'h5:3'h5];
  assign T330 = T334 | T331;
  assign T331 = T333 ? T332 : 13'h0;
  assign T332 = tgts[3'h4];
  assign T333 = hits[3'h4:3'h4];
  assign T334 = T338 | T335;
  assign T335 = T337 ? T336 : 13'h0;
  assign T336 = tgts[3'h3];
  assign T337 = hits[2'h3:2'h3];
  assign T338 = T342 | T339;
  assign T339 = T341 ? T340 : 13'h0;
  assign T340 = tgts[3'h2];
  assign T341 = hits[2'h2:2'h2];
  assign T342 = T346 | T343;
  assign T343 = T345 ? T344 : 13'h0;
  assign T344 = tgts[3'h1];
  assign T345 = hits[1'h1:1'h1];
  assign T346 = T348 ? T347 : 13'h0;
  assign T347 = tgts[3'h0];
  assign T348 = hits[1'h0:1'h0];
  assign T349 = T376 | T350;
  assign T350 = T352 ? T351 : 30'h0;
  assign T351 = pages[2'h3];
  assign T352 = T353[2'h3:2'h3];
  assign T353 = T356 | T354;
  assign T354 = T355 ? T296 : 4'h0;
  assign T355 = hits[3'h7:3'h7];
  assign T356 = T359 | T357;
  assign T357 = T358 ? T290 : 4'h0;
  assign T358 = hits[3'h6:3'h6];
  assign T359 = T362 | T360;
  assign T360 = T361 ? T283 : 4'h0;
  assign T361 = hits[3'h5:3'h5];
  assign T362 = T365 | T363;
  assign T363 = T364 ? T277 : 4'h0;
  assign T364 = hits[3'h4:3'h4];
  assign T365 = T368 | T366;
  assign T366 = T367 ? T269 : 4'h0;
  assign T367 = hits[2'h3:2'h3];
  assign T368 = T371 | T369;
  assign T369 = T370 ? T263 : 4'h0;
  assign T370 = hits[2'h2:2'h2];
  assign T371 = T374 | T372;
  assign T372 = T373 ? T256 : 4'h0;
  assign T373 = hits[1'h1:1'h1];
  assign T374 = T375 ? T242 : 4'h0;
  assign T375 = hits[1'h0:1'h0];
  assign T376 = T380 | T377;
  assign T377 = T379 ? T378 : 30'h0;
  assign T378 = pages[2'h2];
  assign T379 = T353[2'h2:2'h2];
  assign T380 = T384 | T381;
  assign T381 = T383 ? T382 : 30'h0;
  assign T382 = pages[2'h1];
  assign T383 = T353[1'h1:1'h1];
  assign T384 = T386 ? T385 : 30'h0;
  assign T385 = pages[2'h0];
  assign T386 = T353[1'h0:1'h0];
  assign T387 = T421 ? R417 : R388;
  assign T389 = T390 ? io_update_bits_returnAddr : R388;
  assign T390 = T399 & T391;
  assign T391 = T392[1'h0:1'h0];
  assign T392 = 1'h1 << T393;
  assign T393 = T394;
  assign T394 = R395 + 1'h1;
  assign T396 = reset ? 1'h0 : T397;
  assign T397 = T401 ? T400 : T398;
  assign T398 = T399 ? T394 : R395;
  assign T399 = io_update_valid & io_update_bits_isCall;
  assign T400 = R395 - 1'h1;
  assign T401 = T413 & T402;
  assign T402 = T403 ^ 1'h1;
  assign T403 = R404 == 2'h0;
  assign T405 = reset ? 2'h0 : T406;
  assign T406 = io_invalidate ? 2'h0 : T407;
  assign T407 = T401 ? T412 : T408;
  assign T408 = T410 ? T409 : R404;
  assign T409 = R404 + 2'h1;
  assign T410 = T399 & T411;
  assign T411 = R404 < 2'h2;
  assign T412 = R404 - 2'h1;
  assign T413 = io_update_valid & T414;
  assign T414 = T416 & T415;
  assign T415 = io_update_bits_isReturn & io_update_bits_prediction_valid;
  assign T416 = io_update_bits_isCall ^ 1'h1;
  assign T418 = T419 ? io_update_bits_returnAddr : R417;
  assign T419 = T399 & T420;
  assign T420 = T392[1'h1:1'h1];
  assign T421 = R395;
  assign T422 = T438 & T423;
  assign T423 = T424 != 8'h0;
  assign T424 = hits & useRAS;
  assign T425 = T7 ? T426 : useRAS;
  assign T426 = T436 | T427;
  assign T427 = T431 & T428;
  assign T428 = T430 | T429;
  assign T429 = useRAS ^ useRAS;
  assign T430 = 1'h1 << T152;
  assign T431 = T432 ? 8'hff : 8'h0;
  assign T432 = T433;
  assign T433 = R434;
  assign T435 = io_update_valid ? io_update_bits_isReturn : R434;
  assign T436 = useRAS & T437;
  assign T437 = ~ T428;
  assign T438 = T439 ^ 1'h1;
  assign T439 = R404 == 2'h0;
  assign T440 = T399 & T423;
  assign io_resp_bits_taken = T441;
  assign T441 = T442 ? 1'h0 : io_resp_valid;
  assign T442 = T457 & T443;
  assign T443 = T444 ^ 1'h1;
  assign T444 = T445 != 8'h0;
  assign T445 = hits & isJump;
  assign T446 = T7 ? T447 : isJump;
  assign T447 = T455 | T448;
  assign T448 = T452 & T449;
  assign T449 = T451 | T450;
  assign T450 = isJump ^ isJump;
  assign T451 = 1'h1 << T152;
  assign T452 = T453 ? 8'hff : 8'h0;
  assign T453 = T454;
  assign T454 = R37;
  assign T455 = isJump & T456;
  assign T456 = ~ T449;
  assign T457 = T458 ^ 1'h1;
  assign T458 = T18[1'h0:1'h0];
  assign io_resp_valid = T459;
  assign T459 = hits != 8'h0;

  always @(posedge clk) begin
`ifndef SYNTHESIS
  if(reset) T0 <= 1'b1;
  if(!T1 && T0) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BTB request != I$ target");
    $finish;
  end
`endif
    if(io_update_valid) begin
      R4 <= io_update_bits_target;
    end
    if(io_update_valid) begin
      R8 <= io_update_bits_incorrectTarget;
    end
    if(io_update_valid) begin
      R10 <= io_update_bits_prediction_valid;
    end
    if(reset) begin
      R16 <= 1'h0;
    end else begin
      R16 <= io_update_valid;
    end
    if (T35)
      T20[R40] <= T22;
    if(io_update_valid) begin
      R25 <= io_update_bits_taken;
    end
    if(io_update_valid) begin
      R29 <= io_update_bits_prediction_bits_bht_value;
    end
    if(io_update_valid) begin
      R37 <= io_update_bits_isJump;
    end
    if(io_update_valid) begin
      R40 <= io_update_bits_prediction_bits_bht_index;
    end
    if(T35) begin
      R44 <= T46;
    end
    if(reset) begin
      pageValid <= 4'h0;
    end else if(io_invalidate) begin
      pageValid <= 4'h0;
    end else if(T128) begin
      pageValid <= T65;
    end
    if(reset) begin
      R70 <= 2'h0;
    end else if(T74) begin
      R70 <= T73;
    end
    if(io_update_valid) begin
      R86 <= io_update_bits_pc;
    end
    if (T95)
      pages[2'h3] <= T90;
    if (T100)
      pages[2'h1] <= T90;
    if (T107)
      pages[2'h2] <= T104;
    if (T112)
      pages[2'h0] <= T104;
    if (T7)
      idxPages[T152] <= T146;
    if(reset) begin
      R153 <= 3'h0;
    end else if(T157) begin
      R153 <= T156;
    end
    if(io_update_valid) begin
      R160 <= io_update_bits_prediction_bits_entry;
    end
    if (T7)
      idxs[T152] <= T210;
    if(reset) begin
      idxValid <= 8'h0;
    end else if(io_invalidate) begin
      idxValid <= 8'h0;
    end else if(T12) begin
      idxValid <= T299;
    end else if(T12) begin
      idxValid <= T233;
    end
    if (T7)
      tgtPages[T152] <= T246;
    if (T7)
      tgts[T152] <= T320;
    if(T390) begin
      R388 <= io_update_bits_returnAddr;
    end
    if(reset) begin
      R395 <= 1'h0;
    end else if(T401) begin
      R395 <= T400;
    end else if(T399) begin
      R395 <= T394;
    end
    if(reset) begin
      R404 <= 2'h0;
    end else if(io_invalidate) begin
      R404 <= 2'h0;
    end else if(T401) begin
      R404 <= T412;
    end else if(T410) begin
      R404 <= T409;
    end
    if(T419) begin
      R417 <= io_update_bits_returnAddr;
    end
    if(T7) begin
      useRAS <= T426;
    end
    if(io_update_valid) begin
      R434 <= io_update_bits_isReturn;
    end
    if(T7) begin
      isJump <= T447;
    end
  end
endmodule

module FlowThroughSerializer_0(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg  active;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire T12;
  wire[3:0] T13;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[2:0] T16;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T17;
  wire[2:0] T18;
  wire[1:0] T19;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[511:0] T22;
  wire[511:0] T23;
  reg [511:0] rbits_payload_data;
  wire[511:0] T24;
  wire[511:0] T25;
  wire[511:0] T26;
  wire[127:0] T27;
  wire[127:0] T28;
  wire[127:0] shifter_0;
  wire[127:0] T29;
  wire[127:0] shifter_1;
  wire[127:0] T30;
  wire T31;
  wire[1:0] T32;
  wire[127:0] T33;
  wire[127:0] shifter_2;
  wire[127:0] T34;
  wire[127:0] shifter_3;
  wire[127:0] T35;
  wire T36;
  wire T37;
  wire[1:0] T38;
  reg [1:0] rbits_header_dst;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  reg [1:0] rbits_header_src;
  wire[1:0] T42;
  wire[1:0] T43;
  wire T44;
  wire T45;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cnt = {1{$random}};
    active = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T12 & wrap;
  assign wrap = cnt == 2'h3;
  assign T1 = reset ? 2'h0 : T2;
  assign T2 = T0 ? 2'h0 : T3;
  assign T3 = T12 ? T11 : T4;
  assign T4 = T6 ? T5 : cnt;
  assign T5 = {1'h0, io_out_ready};
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T8 = reset ? 1'h0 : T9;
  assign T9 = T0 ? 1'h0 : T10;
  assign T10 = T6 ? 1'h1 : active;
  assign T11 = cnt + 2'h1;
  assign T12 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T13;
  assign T13 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T14 = reset ? io_in_bits_payload_g_type : T15;
  assign T15 = T6 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T17 = reset ? io_in_bits_payload_master_xact_id : T18;
  assign T18 = T6 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T19;
  assign T19 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T20 = reset ? io_in_bits_payload_client_xact_id : T21;
  assign T21 = T6 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T22;
  assign T22 = active ? T26 : T23;
  assign T23 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T24 = reset ? io_in_bits_payload_data : T25;
  assign T25 = T6 ? io_in_bits_payload_data : rbits_payload_data;
  assign T26 = {384'h0, T27};
  assign T27 = T37 ? T33 : T28;
  assign T28 = T31 ? shifter_1 : shifter_0;
  assign shifter_0 = T29;
  assign T29 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T30;
  assign T30 = rbits_payload_data[8'hff:8'h80];
  assign T31 = T32[1'h0:1'h0];
  assign T32 = cnt;
  assign T33 = T36 ? shifter_3 : shifter_2;
  assign shifter_2 = T34;
  assign T34 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T35;
  assign T35 = rbits_payload_data[9'h1ff:9'h180];
  assign T36 = T32[1'h0:1'h0];
  assign T37 = T32[1'h1:1'h1];
  assign io_out_bits_header_dst = T38;
  assign T38 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T39 = reset ? io_in_bits_header_dst : T40;
  assign T40 = T6 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T41;
  assign T41 = active ? rbits_header_src : io_in_bits_header_src;
  assign T42 = reset ? io_in_bits_header_src : T43;
  assign T43 = T6 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T44;
  assign T44 = active | io_in_valid;
  assign io_in_ready = T45;
  assign T45 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      cnt <= 2'h0;
    end else if(T0) begin
      cnt <= 2'h0;
    end else if(T12) begin
      cnt <= T11;
    end else if(T6) begin
      cnt <= T5;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T0) begin
      active <= 1'h0;
    end else if(T6) begin
      active <= 1'h1;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T6) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T6) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T6) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T6) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T6) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T6) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output io_count
);

  wire T0;
  wire[1:0] T1;
  reg  maybe_full;
  wire T2;
  wire T3;
  wire do_enq;
  wire T4;
  wire do_deq;
  wire[2:0] T5;
  wire[6:0] T6;
  reg [6:0] ram [0:0];
  wire[6:0] T7;
  wire[6:0] T8;
  wire[6:0] T9;
  wire[4:0] T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire empty;
  wire T14;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = {maybe_full, 1'h0};
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = T4 ? do_enq : maybe_full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T4 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T5;
  assign T5 = T6[2'h2:1'h0];
  assign T6 = ram[1'h0];
  assign T8 = T9;
  assign T9 = {io_enq_bits_header_src, T10};
  assign T10 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign io_deq_bits_header_dst = T11;
  assign T11 = T6[3'h4:2'h3];
  assign io_deq_bits_header_src = T12;
  assign T12 = T6[3'h6:3'h5];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign io_enq_ready = T14;
  assign T14 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T4) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T8;
  end
endmodule

module ICache(input clk, input reset,
    input  io_req_valid,
    input [12:0] io_req_bits_idx,
    input [18:0] io_req_bits_ppn,
    input  io_req_bits_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[31:0] io_resp_bits_data,
    output[127:0] io_resp_bits_datablock,
    input  io_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[2:0] FlowThroughSerializer_io_out_bits_payload_master_xact_id;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_src;
  wire T0;
  wire T1;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_g_type;
  wire FlowThroughSerializer_io_done;
  wire[2:0] ack_q_io_deq_bits_payload_master_xact_id;
  wire[1:0] ack_q_io_deq_bits_header_dst;
  wire[1:0] ack_q_io_deq_bits_header_src;
  wire ack_q_io_deq_valid;
  wire FlowThroughSerializer_io_in_ready;
  wire[3:0] T2;
  wire[2:0] T3;
  wire[5:0] T4;
  wire[2:0] T5;
  wire[511:0] T6;
  wire[1:0] T7;
  wire[25:0] T8;
  wire[25:0] T9;
  reg [31:0] s2_addr;
  wire[31:0] T10;
  wire[31:0] s1_addr;
  wire[31:0] T11;
  reg [12:0] s1_pgoff;
  wire[12:0] T12;
  wire T13;
  wire rdy;
  wire T14;
  wire T15;
  wire s2_miss;
  wire T16;
  wire s2_any_tag_hit;
  wire T17;
  wire T18;
  wire s2_disparity_0;
  wire T19;
  reg  R20;
  wire T21;
  wire T22;
  wire T23;
  wire stall;
  wire T24;
  reg  s1_valid;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  reg  R31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[5:0] T40;
  wire T41;
  reg [63:0] vb_array;
  wire[63:0] T42;
  wire[127:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[127:0] T46;
  wire[127:0] T47;
  wire[127:0] T48;
  wire[127:0] T49;
  wire[127:0] T50;
  wire[6:0] T51;
  wire[5:0] T52;
  wire[127:0] T53;
  wire T54;
  wire[127:0] T55;
  wire[127:0] T56;
  wire[127:0] T57;
  wire T58;
  wire T59;
  reg  invalidated;
  wire T60;
  wire T61;
  wire T62;
  reg [1:0] state;
  wire[1:0] T63;
  wire[1:0] T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire ack_q_io_enq_ready;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire[127:0] T76;
  wire[127:0] T77;
  wire[127:0] T78;
  wire[6:0] T79;
  wire[127:0] T80;
  wire T81;
  wire[127:0] T82;
  wire[127:0] T83;
  wire[127:0] T84;
  wire T85;
  reg  s2_valid;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire s2_tag_hit_0;
  wire T92;
  reg  R93;
  wire T94;
  wire s1_tag_match_0;
  wire T95;
  wire[19:0] T96;
  wire[19:0] T97;
  wire[19:0] T98;
  wire[19:0] T99;
  wire T100;
  wire s0_valid;
  wire T101;
  wire T102;
  wire[5:0] T103;
  wire[12:0] s0_pgoff;
  wire T104;
  wire[19:0] T105;
  wire[19:0] T106;
  wire[19:0] T107;
  wire[19:0] T108;
  reg [5:0] tag_raddr;
  wire[5:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  reg [127:0] s2_dout_0;
  wire[127:0] T116;
  wire[127:0] T117;
  wire T118;
  wire T119;
  wire FlowThroughSerializer_io_out_valid;
  wire[7:0] T120;
  wire[127:0] T122;
  wire[127:0] T123;
  wire[511:0] FlowThroughSerializer_io_out_bits_payload_data;
  wire[7:0] T124;
  wire[1:0] FlowThroughSerializer_io_cnt;
  reg [7:0] R125;
  wire[7:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire[31:0] T130;
  wire[127:0] T131;
  wire[6:0] T132;
  wire[1:0] T133;
  wire[5:0] T134;
  wire s2_hit;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_addr = {1{$random}};
    s1_pgoff = {1{$random}};
    R20 = {1{$random}};
    s1_valid = {1{$random}};
    R31 = {1{$random}};
    vb_array = {2{$random}};
    invalidated = {1{$random}};
    state = {1{$random}};
    s2_valid = {1{$random}};
    R93 = {1{$random}};
    tag_raddr = {1{$random}};
    s2_dout_0 = {4{$random}};
    R125 = {1{$random}};
  end
`endif

  assign T0 = FlowThroughSerializer_io_done & T1;
  assign T1 = FlowThroughSerializer_io_out_bits_payload_g_type != 4'h0;
  assign io_mem_finish_bits_payload_master_xact_id = ack_q_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ack_q_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ack_q_io_deq_bits_header_src;
  assign io_mem_finish_valid = ack_q_io_deq_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T2;
  assign T2 = 4'h0;
  assign io_mem_acquire_bits_payload_subword_addr = T3;
  assign T3 = 3'h0;
  assign io_mem_acquire_bits_payload_write_mask = T4;
  assign T4 = 6'h0;
  assign io_mem_acquire_bits_payload_a_type = T5;
  assign T5 = 3'h2;
  assign io_mem_acquire_bits_payload_data = T6;
  assign T6 = 512'h0;
  assign io_mem_acquire_bits_payload_client_xact_id = T7;
  assign T7 = 2'h0;
  assign io_mem_acquire_bits_payload_addr = T8;
  assign T8 = T9;
  assign T9 = s2_addr >> 3'h6;
  assign T10 = T111 ? s1_addr : s2_addr;
  assign s1_addr = T11;
  assign T11 = {io_req_bits_ppn, s1_pgoff};
  assign T12 = T13 ? io_req_bits_idx : s1_pgoff;
  assign T13 = io_req_valid & rdy;
  assign rdy = T14;
  assign T14 = T110 & T15;
  assign T15 = s2_miss ^ 1'h1;
  assign s2_miss = s2_valid & T16;
  assign T16 = s2_any_tag_hit ^ 1'h1;
  assign s2_any_tag_hit = T17;
  assign T17 = s2_tag_hit_0 & T18;
  assign T18 = s2_disparity_0 ^ 1'h1;
  assign s2_disparity_0 = T19;
  assign T19 = R31 & R20;
  assign T21 = T22 ? 1'h0 : R20;
  assign T22 = T24 & T23;
  assign T23 = stall ^ 1'h1;
  assign stall = io_resp_ready ^ 1'h1;
  assign T24 = s1_valid & rdy;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T30 | T27;
  assign T27 = T29 & T28;
  assign T28 = io_req_bits_kill ^ 1'h1;
  assign T29 = s1_valid & stall;
  assign T30 = io_req_valid & rdy;
  assign T32 = T22 ? T33 : R31;
  assign T33 = T34;
  assign T34 = T41 & T35;
  assign T35 = T36 - 1'h1;
  assign T36 = 1'h1 << T37;
  assign T37 = T38 + 7'h1;
  assign T38 = T39 - T39;
  assign T39 = {1'h0, T40};
  assign T40 = s1_pgoff[4'hb:3'h6];
  assign T41 = vb_array >> T39;
  assign T42 = T43[6'h3f:1'h0];
  assign T43 = reset ? 128'h0 : T44;
  assign T44 = T85 ? T76 : T45;
  assign T45 = io_invalidate ? 128'h0 : T46;
  assign T46 = T58 ? T48 : T47;
  assign T47 = {64'h0, vb_array};
  assign T48 = T55 | T49;
  assign T49 = T53 & T50;
  assign T50 = 1'h1 << T51;
  assign T51 = {1'h0, T52};
  assign T52 = s2_addr[4'hb:3'h6];
  assign T53 = T54 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T54 = 1'h1;
  assign T55 = T57 & T56;
  assign T56 = ~ T50;
  assign T57 = {64'h0, vb_array};
  assign T58 = FlowThroughSerializer_io_done & T59;
  assign T59 = invalidated ^ 1'h1;
  assign T60 = T62 ? 1'h0 : T61;
  assign T61 = io_invalidate ? 1'h1 : invalidated;
  assign T62 = 2'h0 == state;
  assign T63 = reset ? 2'h0 : T64;
  assign T64 = T74 ? 2'h0 : T65;
  assign T65 = T72 ? 2'h3 : T66;
  assign T66 = T69 ? 2'h2 : T67;
  assign T67 = T68 ? 2'h1 : state;
  assign T68 = T62 & s2_miss;
  assign T69 = T71 & T70;
  assign T70 = io_mem_acquire_ready & ack_q_io_enq_ready;
  assign T71 = 2'h1 == state;
  assign T72 = T73 & io_mem_grant_valid;
  assign T73 = 2'h2 == state;
  assign T74 = T75 & FlowThroughSerializer_io_done;
  assign T75 = 2'h3 == state;
  assign T76 = T82 | T77;
  assign T77 = T80 & T78;
  assign T78 = 1'h1 << T79;
  assign T79 = {1'h0, T52};
  assign T80 = T81 ? 128'hffffffffffffffffffffffffffffffff : 128'h0;
  assign T81 = 1'h0;
  assign T82 = T84 & T83;
  assign T83 = ~ T78;
  assign T84 = {64'h0, vb_array};
  assign T85 = s2_valid & s2_disparity_0;
  assign T86 = reset ? 1'h0 : T87;
  assign T87 = T89 | T88;
  assign T88 = io_resp_valid & stall;
  assign T89 = T91 & T90;
  assign T90 = io_req_bits_kill ^ 1'h1;
  assign T91 = s1_valid & rdy;
  assign s2_tag_hit_0 = T92;
  assign T92 = R31 & R93;
  assign T94 = T22 ? s1_tag_match_0 : R93;
  assign s1_tag_match_0 = T95;
  assign T95 = T97 == T96;
  assign T96 = s1_addr[5'h1f:4'hc];
  assign T97 = T98[5'h13:1'h0];
  assign T98 = T99[5'h13:1'h0];
  assign T100 = T102 & s0_valid;
  assign s0_valid = io_req_valid | T101;
  assign T101 = s1_valid & stall;
  assign T102 = FlowThroughSerializer_io_done ^ 1'h1;
  assign T103 = s0_pgoff[4'hb:3'h6];
  assign s0_pgoff = T104 ? s1_pgoff : io_req_bits_idx;
  assign T104 = s1_valid & stall;
  ICache_tag_array tag_array (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_io_done ? T52 : T103),
    .RW0E(T100 || FlowThroughSerializer_io_done),
    .RW0W(FlowThroughSerializer_io_done),
    .RW0I(T107),
    .RW0M(T106),
    .RW0O(T99)
  );
  assign T106 = 20'hfffff;
  assign T107 = T108;
  assign T108 = s2_addr[5'h1f:4'hc];
  assign T109 = T100 ? T103 : tag_raddr;
  assign T110 = state == 2'h0;
  assign T111 = T113 & T112;
  assign T112 = stall ^ 1'h1;
  assign T113 = s1_valid & rdy;
  assign io_mem_acquire_valid = T114;
  assign T114 = T115 & ack_q_io_enq_ready;
  assign T115 = state == 2'h1;
  assign io_resp_bits_datablock = s2_dout_0;
  assign T116 = T127 ? T117 : s2_dout_0;
  assign T118 = T119 & s0_valid;
  assign T119 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T120 = s0_pgoff[4'hb:3'h4];
  ICache_T121 T121 (
    .CLK(clk),
    .RW0A(FlowThroughSerializer_io_out_valid ? T124 : T120),
    .RW0E(T118 || FlowThroughSerializer_io_out_valid),
    .RW0W(FlowThroughSerializer_io_out_valid),
    .RW0I(T123),
    .RW0O(T117)
  );
  assign T123 = FlowThroughSerializer_io_out_bits_payload_data[7'h7f:1'h0];
  assign T124 = {T52, FlowThroughSerializer_io_cnt};
  assign T126 = T118 ? T120 : R125;
  assign T127 = T129 & T128;
  assign T128 = stall ^ 1'h1;
  assign T129 = s1_valid & rdy;
  assign io_resp_bits_data = T130;
  assign T130 = T131[5'h1f:1'h0];
  assign T131 = s2_dout_0 >> T132;
  assign T132 = T133 << 3'h5;
  assign T133 = T134[2'h3:2'h2];
  assign T134 = s2_addr[3'h5:1'h0];
  assign io_resp_valid = s2_hit;
  assign s2_hit = s2_valid & s2_any_tag_hit;
  FlowThroughSerializer_0 FlowThroughSerializer(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( 1'h1 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       //.io_out_bits_header_dst(  )
       .io_out_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       //.io_out_bits_payload_client_xact_id(  )
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type ),
       .io_cnt( FlowThroughSerializer_io_cnt ),
       .io_done( FlowThroughSerializer_io_done )
  );
  Queue_0 ack_q(.clk(clk), .reset(reset),
       .io_enq_ready( ack_q_io_enq_ready ),
       .io_enq_valid( T0 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( FlowThroughSerializer_io_out_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_deq_ready( io_mem_finish_ready ),
       .io_deq_valid( ack_q_io_deq_valid ),
       .io_deq_bits_header_src( ack_q_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ack_q_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ack_q_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ack_q.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(T111) begin
      s2_addr <= s1_addr;
    end
    if(T13) begin
      s1_pgoff <= io_req_bits_idx;
    end
    if(T22) begin
      R20 <= 1'h0;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T26;
    end
    if(T22) begin
      R31 <= T33;
    end
    vb_array <= T42;
    if(T62) begin
      invalidated <= 1'h0;
    end else if(io_invalidate) begin
      invalidated <= 1'h1;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T74) begin
      state <= 2'h0;
    end else if(T72) begin
      state <= 2'h3;
    end else if(T69) begin
      state <= 2'h2;
    end else if(T68) begin
      state <= 2'h1;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= T87;
    end
    if(T22) begin
      R93 <= s1_tag_match_0;
    end
    if(T100) begin
      tag_raddr <= T103;
    end
    if(T127) begin
      s2_dout_0 <= T117;
    end
    if(T118) begin
      R125 <= T120;
    end
  end
endmodule

module RocketCAM(input clk, input reset,
    input  io_clear,
    input  io_clear_hit,
    input [36:0] io_tag,
    output io_hit,
    output[3:0] io_hits,
    output[3:0] io_valid_bits,
    input  io_write,
    input [36:0] io_write_tag,
    input [1:0] io_write_addr
);

  reg [3:0] vb_array;
  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[1:0] T17;
  wire hits_0;
  wire T18;
  wire[36:0] T19;
  reg [36:0] cam_tags [3:0];
  wire[36:0] T20;
  wire T21;
  wire hits_1;
  wire T22;
  wire[36:0] T23;
  wire T24;
  wire[1:0] T25;
  wire hits_2;
  wire T26;
  wire[36:0] T27;
  wire T28;
  wire hits_3;
  wire T29;
  wire[36:0] T30;
  wire T31;
  wire T32;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    vb_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      cam_tags[initvar] = {2{$random}};
  end
`endif

  assign io_valid_bits = vb_array;
  assign T0 = reset ? 4'h0 : T1;
  assign T1 = T13 ? T11 : T2;
  assign T2 = io_clear ? 4'h0 : T3;
  assign T3 = io_write ? T4 : vb_array;
  assign T4 = T9 | T5;
  assign T5 = T7 & T6;
  assign T6 = 1'h1 << io_write_addr;
  assign T7 = T8 ? 4'hf : 4'h0;
  assign T8 = 1'h1;
  assign T9 = vb_array & T10;
  assign T10 = ~ T6;
  assign T11 = vb_array & T12;
  assign T12 = ~ io_hits;
  assign T13 = T14 & io_clear_hit;
  assign T14 = io_clear ^ 1'h1;
  assign io_hits = T15;
  assign T15 = T16;
  assign T16 = {T25, T17};
  assign T17 = {hits_1, hits_0};
  assign hits_0 = T21 & T18;
  assign T18 = T19 == io_tag;
  assign T19 = cam_tags[2'h0];
  assign T21 = vb_array[1'h0:1'h0];
  assign hits_1 = T24 & T22;
  assign T22 = T23 == io_tag;
  assign T23 = cam_tags[2'h1];
  assign T24 = vb_array[1'h1:1'h1];
  assign T25 = {hits_3, hits_2};
  assign hits_2 = T28 & T26;
  assign T26 = T27 == io_tag;
  assign T27 = cam_tags[2'h2];
  assign T28 = vb_array[2'h2:2'h2];
  assign hits_3 = T31 & T29;
  assign T29 = T30 == io_tag;
  assign T30 = cam_tags[2'h3];
  assign T31 = vb_array[2'h3:2'h3];
  assign io_hit = T32;
  assign T32 = io_hits != 4'h0;

  always @(posedge clk) begin
    if(reset) begin
      vb_array <= 4'h0;
    end else if(T13) begin
      vb_array <= T11;
    end else if(io_clear) begin
      vb_array <= 4'h0;
    end else if(io_write) begin
      vb_array <= T4;
    end
    if (io_write)
      cam_tags[io_write_addr] <= io_write_tag;
  end
endmodule

module TLB(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [6:0] io_req_bits_asid,
    input [30:0] io_req_bits_vpn,
    input  io_req_bits_passthrough,
    input  io_req_bits_instruction,
    output io_resp_miss,
    output[3:0] io_resp_hit_idx,
    output[18:0] io_resp_ppn,
    output io_resp_xcpt_ld,
    output io_resp_xcpt_st,
    output io_resp_xcpt_if,
    input  io_ptw_req_ready,
    output io_ptw_req_valid,
    output[29:0] io_ptw_req_bits,
    input  io_ptw_resp_valid,
    input  io_ptw_resp_bits_error,
    input [18:0] io_ptw_resp_bits_ppn,
    input [5:0] io_ptw_resp_bits_perm,
    input [7:0] io_ptw_status_ip,
    input [7:0] io_ptw_status_im,
    input [6:0] io_ptw_status_zero,
    input  io_ptw_status_er,
    input  io_ptw_status_vm,
    input  io_ptw_status_s64,
    input  io_ptw_status_u64,
    input  io_ptw_status_ef,
    input  io_ptw_status_pei,
    input  io_ptw_status_ei,
    input  io_ptw_status_ps,
    input  io_ptw_status_s,
    input  io_ptw_invalidate,
    input  io_ptw_sret
);

  reg [1:0] r_refill_waddr;
  wire[1:0] T0;
  wire[1:0] repl_waddr;
  wire[1:0] T1;
  wire[2:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  reg [3:0] R10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[6:0] T15;
  wire[1:0] T16;
  wire T17;
  wire[1:0] T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[3:0] tag_cam_io_hits;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire[3:0] T25;
  wire[3:0] T26;
  wire[3:0] T27;
  wire[3:0] T28;
  wire[3:0] T29;
  wire T30;
  wire tlb_hit;
  wire tag_cam_io_hit;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire[1:0] T34;
  wire T35;
  wire[3:0] T36;
  wire[3:0] tag_cam_io_valid_bits;
  wire T37;
  wire T38;
  wire has_invalid_entry;
  wire T39;
  wire T40;
  wire tlb_miss;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire[36:0] T48;
  reg [37:0] r_refill_tag;
  wire[37:0] T49;
  wire[37:0] lookup_tag;
  wire[37:0] T50;
  wire T51;
  wire T52;
  reg [1:0] state;
  wire[1:0] T53;
  wire[1:0] T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire[36:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire[29:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[3:0] T78;
  reg [3:0] ux_array;
  wire[3:0] T79;
  wire[3:0] T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire[5:0] T86;
  wire[5:0] T87;
  wire T88;
  wire T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire T92;
  wire[3:0] T93;
  reg [3:0] sx_array;
  wire[3:0] T94;
  wire[3:0] T95;
  wire[3:0] T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire T99;
  wire T100;
  wire[3:0] T101;
  wire[3:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire[3:0] T108;
  reg [3:0] uw_array;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T112;
  wire[3:0] T113;
  wire T114;
  wire T115;
  wire[3:0] T116;
  wire[3:0] T117;
  wire T118;
  wire[3:0] T119;
  reg [3:0] sw_array;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] T124;
  wire T125;
  wire T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire[3:0] T134;
  reg [3:0] ur_array;
  wire[3:0] T135;
  wire[3:0] T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire T140;
  wire T141;
  wire[3:0] T142;
  wire[3:0] T143;
  wire T144;
  wire[3:0] T145;
  reg [3:0] sr_array;
  wire[3:0] T146;
  wire[3:0] T147;
  wire[3:0] T148;
  wire[3:0] T149;
  wire[3:0] T150;
  wire T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] T154;
  wire[18:0] T155;
  wire[18:0] T156;
  wire[18:0] T157;
  wire[18:0] T158;
  wire[18:0] T159;
  reg [18:0] tag_ram [3:0];
  wire[18:0] T160;
  wire T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[18:0] T164;
  wire T165;
  wire[18:0] T166;
  wire[18:0] T167;
  wire[18:0] T168;
  wire T169;
  wire[18:0] T170;
  wire[18:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_refill_waddr = {1{$random}};
    R10 = {1{$random}};
    r_refill_tag = {2{$random}};
    state = {1{$random}};
    ux_array = {1{$random}};
    sx_array = {1{$random}};
    uw_array = {1{$random}};
    sw_array = {1{$random}};
    ur_array = {1{$random}};
    sr_array = {1{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      tag_ram[initvar] = {1{$random}};
  end
`endif

  assign T0 = T40 ? repl_waddr : r_refill_waddr;
  assign repl_waddr = has_invalid_entry ? T32 : T1;
  assign T1 = T2[1'h1:1'h0];
  assign T2 = {T8, T3};
  assign T3 = T31 & T4;
  assign T4 = T5 - 1'h1;
  assign T5 = 1'h1 << T6;
  assign T6 = T7 + 2'h1;
  assign T7 = T8 - T8;
  assign T8 = {1'h1, T9};
  assign T9 = R10[1'h1:1'h1];
  assign T11 = T30 ? T12 : R10;
  assign T12 = T25 | T13;
  assign T13 = T24 ? 4'h0 : T14;
  assign T14 = T15[2'h3:1'h0];
  assign T15 = 4'h1 << T16;
  assign T16 = {1'h1, T17};
  assign T17 = T18[1'h1:1'h1];
  assign T18 = {T23, T19};
  assign T19 = T20[1'h1:1'h1];
  assign T20 = T22 | T21;
  assign T21 = tag_cam_io_hits[1'h1:1'h0];
  assign T22 = tag_cam_io_hits[2'h3:2'h2];
  assign T23 = T22 != 2'h0;
  assign T24 = T18[1'h0:1'h0];
  assign T25 = T27 & T26;
  assign T26 = ~ T14;
  assign T27 = T29 | T28;
  assign T28 = T17 ? 4'h0 : 4'h2;
  assign T29 = R10 & 4'hd;
  assign T30 = io_req_valid & tlb_hit;
  assign tlb_hit = io_ptw_status_vm & tag_cam_io_hit;
  assign T31 = R10 >> T8;
  assign T32 = T38 ? 1'h0 : T33;
  assign T33 = T37 ? 1'h1 : T34;
  assign T34 = T35 ? 2'h2 : 2'h3;
  assign T35 = T36[2'h2:2'h2];
  assign T36 = ~ tag_cam_io_valid_bits;
  assign T37 = T36[1'h1:1'h1];
  assign T38 = T36[1'h0:1'h0];
  assign has_invalid_entry = T39 ^ 1'h1;
  assign T39 = tag_cam_io_valid_bits == 4'hf;
  assign T40 = T47 & tlb_miss;
  assign tlb_miss = T45 & T41;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T44 != T43;
  assign T43 = io_req_bits_vpn[5'h1d:5'h1d];
  assign T44 = io_req_bits_vpn[5'h1e:5'h1e];
  assign T45 = io_ptw_status_vm & T46;
  assign T46 = tag_cam_io_hit ^ 1'h1;
  assign T47 = io_req_ready & io_req_valid;
  assign T48 = r_refill_tag[6'h24:1'h0];
  assign T49 = T40 ? lookup_tag : r_refill_tag;
  assign lookup_tag = T50;
  assign T50 = {io_req_bits_asid, io_req_bits_vpn};
  assign T51 = T52 & io_ptw_resp_valid;
  assign T52 = state == 2'h2;
  assign T53 = reset ? 2'h0 : T54;
  assign T54 = io_ptw_resp_valid ? 2'h0 : T55;
  assign T55 = T64 ? 2'h3 : T56;
  assign T56 = T63 ? 2'h3 : T57;
  assign T57 = T62 ? 2'h2 : T58;
  assign T58 = T60 ? 2'h0 : T59;
  assign T59 = T40 ? 2'h1 : state;
  assign T60 = T61 & io_ptw_invalidate;
  assign T61 = state == 2'h1;
  assign T62 = T61 & io_ptw_req_ready;
  assign T63 = T62 & io_ptw_invalidate;
  assign T64 = T65 & io_ptw_invalidate;
  assign T65 = state == 2'h2;
  assign T66 = lookup_tag[6'h24:1'h0];
  assign T67 = T70 & T68;
  assign T68 = io_req_bits_instruction ? io_resp_xcpt_if : T69;
  assign T69 = io_resp_xcpt_ld & io_resp_xcpt_st;
  assign T70 = io_req_ready & io_req_valid;
  assign io_ptw_req_bits = T71;
  assign T71 = r_refill_tag[5'h1d:1'h0];
  assign io_ptw_req_valid = T72;
  assign T72 = state == 2'h1;
  assign io_resp_xcpt_if = T73;
  assign T73 = T42 | T74;
  assign T74 = tlb_hit & T75;
  assign T75 = T76 ^ 1'h1;
  assign T76 = io_ptw_status_s ? T92 : T77;
  assign T77 = T78 != 4'h0;
  assign T78 = ux_array & tag_cam_io_hits;
  assign T79 = io_ptw_resp_valid ? T80 : ux_array;
  assign T80 = T90 | T81;
  assign T81 = T83 & T82;
  assign T82 = 1'h1 << r_refill_waddr;
  assign T83 = T84 ? 4'hf : 4'h0;
  assign T84 = T85;
  assign T85 = T86[2'h2:2'h2];
  assign T86 = T87 & io_ptw_resp_bits_perm;
  assign T87 = T88 ? 6'h3f : 6'h0;
  assign T88 = T89;
  assign T89 = io_ptw_resp_bits_error ^ 1'h1;
  assign T90 = ux_array & T91;
  assign T91 = ~ T82;
  assign T92 = T93 != 4'h0;
  assign T93 = sx_array & tag_cam_io_hits;
  assign T94 = io_ptw_resp_valid ? T95 : sx_array;
  assign T95 = T101 | T96;
  assign T96 = T98 & T97;
  assign T97 = 1'h1 << r_refill_waddr;
  assign T98 = T99 ? 4'hf : 4'h0;
  assign T99 = T100;
  assign T100 = T86[3'h5:3'h5];
  assign T101 = sx_array & T102;
  assign T102 = ~ T97;
  assign io_resp_xcpt_st = T103;
  assign T103 = T42 | T104;
  assign T104 = tlb_hit & T105;
  assign T105 = T106 ^ 1'h1;
  assign T106 = io_ptw_status_s ? T118 : T107;
  assign T107 = T108 != 4'h0;
  assign T108 = uw_array & tag_cam_io_hits;
  assign T109 = io_ptw_resp_valid ? T110 : uw_array;
  assign T110 = T116 | T111;
  assign T111 = T113 & T112;
  assign T112 = 1'h1 << r_refill_waddr;
  assign T113 = T114 ? 4'hf : 4'h0;
  assign T114 = T115;
  assign T115 = T86[1'h1:1'h1];
  assign T116 = uw_array & T117;
  assign T117 = ~ T112;
  assign T118 = T119 != 4'h0;
  assign T119 = sw_array & tag_cam_io_hits;
  assign T120 = io_ptw_resp_valid ? T121 : sw_array;
  assign T121 = T127 | T122;
  assign T122 = T124 & T123;
  assign T123 = 1'h1 << r_refill_waddr;
  assign T124 = T125 ? 4'hf : 4'h0;
  assign T125 = T126;
  assign T126 = T86[3'h4:3'h4];
  assign T127 = sw_array & T128;
  assign T128 = ~ T123;
  assign io_resp_xcpt_ld = T129;
  assign T129 = T42 | T130;
  assign T130 = tlb_hit & T131;
  assign T131 = T132 ^ 1'h1;
  assign T132 = io_ptw_status_s ? T144 : T133;
  assign T133 = T134 != 4'h0;
  assign T134 = ur_array & tag_cam_io_hits;
  assign T135 = io_ptw_resp_valid ? T136 : ur_array;
  assign T136 = T142 | T137;
  assign T137 = T139 & T138;
  assign T138 = 1'h1 << r_refill_waddr;
  assign T139 = T140 ? 4'hf : 4'h0;
  assign T140 = T141;
  assign T141 = T86[1'h0:1'h0];
  assign T142 = ur_array & T143;
  assign T143 = ~ T138;
  assign T144 = T145 != 4'h0;
  assign T145 = sr_array & tag_cam_io_hits;
  assign T146 = io_ptw_resp_valid ? T147 : sr_array;
  assign T147 = T153 | T148;
  assign T148 = T150 & T149;
  assign T149 = 1'h1 << r_refill_waddr;
  assign T150 = T151 ? 4'hf : 4'h0;
  assign T151 = T152;
  assign T152 = T86[2'h3:2'h3];
  assign T153 = sr_array & T154;
  assign T154 = ~ T149;
  assign io_resp_ppn = T155;
  assign T155 = T173 ? T157 : T156;
  assign T156 = io_req_bits_vpn[5'h12:1'h0];
  assign T157 = T162 | T158;
  assign T158 = T161 ? T159 : 19'h0;
  assign T159 = tag_ram[2'h3];
  assign T161 = tag_cam_io_hits[2'h3:2'h3];
  assign T162 = T166 | T163;
  assign T163 = T165 ? T164 : 19'h0;
  assign T164 = tag_ram[2'h2];
  assign T165 = tag_cam_io_hits[2'h2:2'h2];
  assign T166 = T170 | T167;
  assign T167 = T169 ? T168 : 19'h0;
  assign T168 = tag_ram[2'h1];
  assign T169 = tag_cam_io_hits[1'h1:1'h1];
  assign T170 = T172 ? T171 : 19'h0;
  assign T171 = tag_ram[2'h0];
  assign T172 = tag_cam_io_hits[1'h0:1'h0];
  assign T173 = io_ptw_status_vm & T174;
  assign T174 = io_req_bits_passthrough ^ 1'h1;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_resp_miss = tlb_miss;
  assign io_req_ready = T175;
  assign T175 = state == 2'h0;
  RocketCAM tag_cam(.clk(clk), .reset(reset),
       .io_clear( io_ptw_invalidate ),
       .io_clear_hit( T67 ),
       .io_tag( T66 ),
       .io_hit( tag_cam_io_hit ),
       .io_hits( tag_cam_io_hits ),
       .io_valid_bits( tag_cam_io_valid_bits ),
       .io_write( T51 ),
       .io_write_tag( T48 ),
       .io_write_addr( r_refill_waddr )
  );

  always @(posedge clk) begin
    if(T40) begin
      r_refill_waddr <= repl_waddr;
    end
    if(T30) begin
      R10 <= T12;
    end
    if(T40) begin
      r_refill_tag <= lookup_tag;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(io_ptw_resp_valid) begin
      state <= 2'h0;
    end else if(T64) begin
      state <= 2'h3;
    end else if(T63) begin
      state <= 2'h3;
    end else if(T62) begin
      state <= 2'h2;
    end else if(T60) begin
      state <= 2'h0;
    end else if(T40) begin
      state <= 2'h1;
    end
    if(io_ptw_resp_valid) begin
      ux_array <= T80;
    end
    if(io_ptw_resp_valid) begin
      sx_array <= T95;
    end
    if(io_ptw_resp_valid) begin
      uw_array <= T110;
    end
    if(io_ptw_resp_valid) begin
      sw_array <= T121;
    end
    if(io_ptw_resp_valid) begin
      ur_array <= T136;
    end
    if(io_ptw_resp_valid) begin
      sr_array <= T147;
    end
    if (io_ptw_resp_valid)
      tag_ram[r_refill_waddr] <= io_ptw_resp_bits_ppn;
  end
endmodule

module Frontend(input clk, input reset,
    input  io_cpu_req_valid,
    input [43:0] io_cpu_req_bits_pc,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[43:0] io_cpu_resp_bits_pc,
    output[31:0] io_cpu_resp_bits_data,
    output io_cpu_resp_bits_xcpt_ma,
    output io_cpu_resp_bits_xcpt_if,
    output io_cpu_btb_resp_valid,
    output io_cpu_btb_resp_bits_taken,
    output[42:0] io_cpu_btb_resp_bits_target,
    output[2:0] io_cpu_btb_resp_bits_entry,
    output[3:0] io_cpu_btb_resp_bits_bht_index,
    output[1:0] io_cpu_btb_resp_bits_bht_value,
    input  io_cpu_btb_update_valid,
    input  io_cpu_btb_update_bits_prediction_valid,
    input  io_cpu_btb_update_bits_prediction_bits_taken,
    input [42:0] io_cpu_btb_update_bits_prediction_bits_target,
    input [2:0] io_cpu_btb_update_bits_prediction_bits_entry,
    input [3:0] io_cpu_btb_update_bits_prediction_bits_bht_index,
    input [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
    input [42:0] io_cpu_btb_update_bits_pc,
    input [42:0] io_cpu_btb_update_bits_target,
    input [42:0] io_cpu_btb_update_bits_returnAddr,
    input  io_cpu_btb_update_bits_taken,
    input  io_cpu_btb_update_bits_isJump,
    input  io_cpu_btb_update_bits_isCall,
    input  io_cpu_btb_update_bits_isReturn,
    input  io_cpu_btb_update_bits_incorrectTarget,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    input  io_cpu_invalidate,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    //output[1:0] io_mem_acquire_bits_header_src
    //output[1:0] io_mem_acquire_bits_header_dst
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id
);

  wire[30:0] T0;
  wire[43:0] s1_pc;
  reg [43:0] s1_pc_;
  wire[43:0] T1;
  wire[43:0] T2;
  wire[43:0] npc;
  wire[43:0] T3;
  wire[43:0] predicted_npc;
  wire[43:0] pcp4;
  wire[42:0] T4;
  wire[43:0] pcp4_0;
  wire T5;
  wire T6;
  wire T7;
  wire[43:0] btbTarget;
  wire[42:0] btb_io_resp_bits_target;
  wire T8;
  wire btb_io_resp_bits_taken;
  reg [43:0] s2_pc;
  wire[43:0] T9;
  wire[43:0] T10;
  wire T11;
  wire T12;
  wire icmiss;
  wire T13;
  wire icache_io_resp_valid;
  reg  s2_valid;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire stall;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg  s1_same_block;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire tlb_io_resp_miss;
  wire s0_same_block;
  wire T29;
  wire[43:0] T30;
  wire[43:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[18:0] tlb_io_resp_ppn;
  wire[12:0] T40;
  wire[43:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire[42:0] T46;
  wire[43:0] T47;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire icache_io_mem_finish_valid;
  wire icache_io_mem_grant_ready;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire icache_io_mem_acquire_valid;
  wire[29:0] tlb_io_ptw_req_bits;
  wire tlb_io_ptw_req_valid;
  reg [1:0] s2_btb_resp_bits_bht_value;
  wire[1:0] T48;
  wire[1:0] btb_io_resp_bits_bht_value;
  wire T49;
  wire btb_io_resp_valid;
  reg [3:0] s2_btb_resp_bits_bht_index;
  wire[3:0] T50;
  wire[3:0] btb_io_resp_bits_bht_index;
  reg [2:0] s2_btb_resp_bits_entry;
  wire[2:0] T51;
  wire[2:0] btb_io_resp_bits_entry;
  reg [42:0] s2_btb_resp_bits_target;
  wire[42:0] T52;
  reg  s2_btb_resp_bits_taken;
  wire T53;
  reg  s2_btb_resp_valid;
  wire T54;
  wire T55;
  reg  s2_xcpt_if;
  wire T56;
  wire T57;
  wire tlb_io_resp_xcpt_if;
  wire T58;
  wire[1:0] T59;
  wire[31:0] T60;
  wire[127:0] T61;
  wire[6:0] T62;
  wire[1:0] T63;
  wire[127:0] icache_io_resp_bits_datablock;
  wire[43:0] T64;
  wire T65;
  wire T66;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s1_pc_ = {2{$random}};
    s2_pc = {2{$random}};
    s2_valid = {1{$random}};
    s1_same_block = {1{$random}};
    s2_btb_resp_bits_bht_value = {1{$random}};
    s2_btb_resp_bits_bht_index = {1{$random}};
    s2_btb_resp_bits_entry = {1{$random}};
    s2_btb_resp_bits_target = {2{$random}};
    s2_btb_resp_bits_taken = {1{$random}};
    s2_btb_resp_valid = {1{$random}};
    s2_xcpt_if = {1{$random}};
  end
`endif

  assign T0 = s1_pc >> 4'hd;
  assign s1_pc = s1_pc_ & 44'hffffffffffe;
  assign T1 = io_cpu_req_valid ? io_cpu_req_bits_pc : T2;
  assign T2 = T18 ? npc : s1_pc_;
  assign npc = T3;
  assign T3 = icmiss ? s2_pc : predicted_npc;
  assign predicted_npc = btb_io_resp_bits_taken ? btbTarget : pcp4;
  assign pcp4 = {T5, T4};
  assign T4 = pcp4_0[6'h2a:1'h0];
  assign pcp4_0 = s1_pc + 44'h4;
  assign T5 = T7 & T6;
  assign T6 = pcp4_0[6'h2a:6'h2a];
  assign T7 = s1_pc[6'h2a:6'h2a];
  assign btbTarget = {T8, btb_io_resp_bits_target};
  assign T8 = btb_io_resp_bits_target[6'h2a:6'h2a];
  assign T9 = reset ? 44'h2000 : T10;
  assign T10 = T11 ? s1_pc : s2_pc;
  assign T11 = T18 & T12;
  assign T12 = icmiss ^ 1'h1;
  assign icmiss = s2_valid & T13;
  assign T13 = icache_io_resp_valid ^ 1'h1;
  assign T14 = reset ? 1'h1 : T15;
  assign T15 = io_cpu_req_valid ? 1'h0 : T16;
  assign T16 = T18 ? T17 : s2_valid;
  assign T17 = icmiss ^ 1'h1;
  assign T18 = stall ^ 1'h1;
  assign stall = io_cpu_resp_valid & T19;
  assign T19 = io_cpu_resp_ready ^ 1'h1;
  assign T20 = T22 & T21;
  assign T21 = icmiss ^ 1'h1;
  assign T22 = stall ^ 1'h1;
  assign T23 = T37 & T24;
  assign T24 = s1_same_block ^ 1'h1;
  assign T25 = io_cpu_req_valid ? 1'h0 : T26;
  assign T26 = T18 ? T27 : s1_same_block;
  assign T27 = s0_same_block & T28;
  assign T28 = tlb_io_resp_miss ^ 1'h1;
  assign s0_same_block = T32 & T29;
  assign T29 = T31 == T30;
  assign T30 = s1_pc & 44'h10;
  assign T31 = pcp4 & 44'h10;
  assign T32 = T34 & T33;
  assign T33 = btb_io_resp_bits_taken ^ 1'h1;
  assign T34 = T36 & T35;
  assign T35 = io_cpu_req_valid ^ 1'h1;
  assign T36 = icmiss ^ 1'h1;
  assign T37 = stall ^ 1'h1;
  assign T38 = T39 | icmiss;
  assign T39 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T40 = T41[4'hc:1'h0];
  assign T41 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T42 = T44 & T43;
  assign T43 = s0_same_block ^ 1'h1;
  assign T44 = stall ^ 1'h1;
  assign T45 = io_cpu_invalidate | io_cpu_ptw_invalidate;
  assign T46 = T47[6'h2a:1'h0];
  assign T47 = s1_pc & 44'hffffffffffc;
  assign io_mem_finish_bits_payload_master_xact_id = icache_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = icache_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = icache_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = icache_io_mem_finish_valid;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = icache_io_mem_acquire_bits_payload_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = icache_io_mem_acquire_bits_payload_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = icache_io_mem_acquire_bits_payload_write_mask;
  assign io_mem_acquire_bits_payload_a_type = icache_io_mem_acquire_bits_payload_a_type;
  assign io_mem_acquire_bits_payload_data = icache_io_mem_acquire_bits_payload_data;
  assign io_mem_acquire_bits_payload_client_xact_id = icache_io_mem_acquire_bits_payload_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = icache_io_mem_acquire_bits_payload_addr;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_cpu_ptw_req_bits = tlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign T48 = T49 ? btb_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T49 = T11 & btb_io_resp_valid;
  assign io_cpu_btb_resp_bits_bht_index = s2_btb_resp_bits_bht_index;
  assign T50 = T49 ? btb_io_resp_bits_bht_index : s2_btb_resp_bits_bht_index;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign T51 = T49 ? btb_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign T52 = T49 ? btb_io_resp_bits_target : s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign T53 = T49 ? btb_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign T54 = reset ? 1'h0 : T55;
  assign T55 = T11 ? btb_io_resp_valid : s2_btb_resp_valid;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign T56 = reset ? 1'h0 : T57;
  assign T57 = T11 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign io_cpu_resp_bits_xcpt_ma = T58;
  assign T58 = T59 != 2'h0;
  assign T59 = s2_pc[1'h1:1'h0];
  assign io_cpu_resp_bits_data = T60;
  assign T60 = T61[5'h1f:1'h0];
  assign T61 = icache_io_resp_bits_datablock >> T62;
  assign T62 = T63 << 3'h5;
  assign T63 = s2_pc[2'h3:2'h2];
  assign io_cpu_resp_bits_pc = T64;
  assign T64 = s2_pc & 44'hffffffffffc;
  assign io_cpu_resp_valid = T65;
  assign T65 = s2_valid & T66;
  assign T66 = s2_xcpt_if | icache_io_resp_valid;
  BTB btb(.clk(clk), .reset(reset),
       .io_req( T46 ),
       .io_resp_valid( btb_io_resp_valid ),
       .io_resp_bits_taken( btb_io_resp_bits_taken ),
       .io_resp_bits_target( btb_io_resp_bits_target ),
       .io_resp_bits_entry( btb_io_resp_bits_entry ),
       .io_resp_bits_bht_index( btb_io_resp_bits_bht_index ),
       .io_resp_bits_bht_value( btb_io_resp_bits_bht_value ),
       .io_update_valid( io_cpu_btb_update_valid ),
       .io_update_bits_prediction_valid( io_cpu_btb_update_bits_prediction_valid ),
       .io_update_bits_prediction_bits_taken( io_cpu_btb_update_bits_prediction_bits_taken ),
       .io_update_bits_prediction_bits_target( io_cpu_btb_update_bits_prediction_bits_target ),
       .io_update_bits_prediction_bits_entry( io_cpu_btb_update_bits_prediction_bits_entry ),
       .io_update_bits_prediction_bits_bht_index( io_cpu_btb_update_bits_prediction_bits_bht_index ),
       .io_update_bits_prediction_bits_bht_value( io_cpu_btb_update_bits_prediction_bits_bht_value ),
       .io_update_bits_pc( io_cpu_btb_update_bits_pc ),
       .io_update_bits_target( io_cpu_btb_update_bits_target ),
       .io_update_bits_returnAddr( io_cpu_btb_update_bits_returnAddr ),
       .io_update_bits_taken( io_cpu_btb_update_bits_taken ),
       .io_update_bits_isJump( io_cpu_btb_update_bits_isJump ),
       .io_update_bits_isCall( io_cpu_btb_update_bits_isCall ),
       .io_update_bits_isReturn( io_cpu_btb_update_bits_isReturn ),
       .io_update_bits_incorrectTarget( io_cpu_btb_update_bits_incorrectTarget ),
       .io_invalidate( T45 )
  );
  ICache icache(.clk(clk), .reset(reset),
       .io_req_valid( T42 ),
       .io_req_bits_idx( T40 ),
       .io_req_bits_ppn( tlb_io_resp_ppn ),
       .io_req_bits_kill( T38 ),
       .io_resp_ready( T23 ),
       .io_resp_valid( icache_io_resp_valid ),
       //.io_resp_bits_data(  )
       .io_resp_bits_datablock( icache_io_resp_bits_datablock ),
       .io_invalidate( io_cpu_invalidate ),
       .io_mem_acquire_ready( io_mem_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  TLB tlb(.clk(clk), .reset(reset),
       //.io_req_ready(  )
       .io_req_valid( T20 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T0 ),
       .io_req_bits_passthrough( 1'h0 ),
       .io_req_bits_instruction( 1'h1 ),
       .io_resp_miss( tlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( tlb_io_resp_ppn ),
       //.io_resp_xcpt_ld(  )
       //.io_resp_xcpt_st(  )
       .io_resp_xcpt_if( tlb_io_resp_xcpt_if ),
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( tlb_io_ptw_req_valid ),
       .io_ptw_req_bits( tlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );

  always @(posedge clk) begin
    if(io_cpu_req_valid) begin
      s1_pc_ <= io_cpu_req_bits_pc;
    end else if(T18) begin
      s1_pc_ <= npc;
    end
    if(reset) begin
      s2_pc <= 44'h2000;
    end else if(T11) begin
      s2_pc <= s1_pc;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s2_valid <= 1'h0;
    end else if(T18) begin
      s2_valid <= T17;
    end
    if(io_cpu_req_valid) begin
      s1_same_block <= 1'h0;
    end else if(T18) begin
      s1_same_block <= T27;
    end
    if(T49) begin
      s2_btb_resp_bits_bht_value <= btb_io_resp_bits_bht_value;
    end
    if(T49) begin
      s2_btb_resp_bits_bht_index <= btb_io_resp_bits_bht_index;
    end
    if(T49) begin
      s2_btb_resp_bits_entry <= btb_io_resp_bits_entry;
    end
    if(T49) begin
      s2_btb_resp_bits_target <= btb_io_resp_bits_target;
    end
    if(T49) begin
      s2_btb_resp_bits_taken <= btb_io_resp_bits_taken;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else if(T11) begin
      s2_btb_resp_valid <= btb_io_resp_valid;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else if(T11) begin
      s2_xcpt_if <= tlb_io_resp_xcpt_if;
    end
  end
endmodule

module WritebackUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [19:0] io_req_bits_tag,
    input [5:0] io_req_bits_idx,
    input  io_req_bits_way_en,
    input [1:0] io_req_bits_client_xact_id,
    input [2:0] io_req_bits_master_xact_id,
    input [2:0] io_req_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_data_req_ready,
    output io_data_req_valid,
    output io_data_req_bits_way_en,
    output[11:0] io_data_req_bits_addr,
    input [127:0] io_data_resp,
    input  io_release_ready,
    output io_release_valid,
    output[25:0] io_release_bits_addr,
    output[1:0] io_release_bits_client_xact_id,
    output[2:0] io_release_bits_master_xact_id,
    output[511:0] io_release_bits_data,
    output[2:0] io_release_bits_r_type
);

  reg [2:0] req_r_type;
  wire[2:0] T0;
  wire T1;
  reg [511:0] R2;
  wire[511:0] T3;
  wire[511:0] T4;
  wire[383:0] T5;
  wire T6;
  reg  r2_data_req_fired;
  wire T7;
  wire T8;
  reg  r1_data_req_fired;
  wire T9;
  wire T10;
  wire T11;
  reg  active;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  reg [2:0] cnt;
  wire[2:0] T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire[2:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  reg [2:0] req_master_xact_id;
  wire[2:0] T30;
  reg [1:0] req_client_xact_id;
  wire[1:0] T31;
  wire[25:0] T32;
  wire[25:0] T33;
  reg [5:0] req_idx;
  wire[5:0] T34;
  reg [19:0] req_tag;
  wire[19:0] T35;
  wire[11:0] T36;
  wire[7:0] T37;
  wire[1:0] T38;
  reg  req_way_en;
  wire T39;
  wire fire;
  wire T40;
  wire T41;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_r_type = {1{$random}};
    R2 = {16{$random}};
    r2_data_req_fired = {1{$random}};
    r1_data_req_fired = {1{$random}};
    active = {1{$random}};
    cnt = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_idx = {1{$random}};
    req_tag = {1{$random}};
    req_way_en = {1{$random}};
  end
`endif

  assign io_release_bits_r_type = req_r_type;
  assign T0 = T1 ? io_req_bits_r_type : req_r_type;
  assign T1 = io_req_ready & io_req_valid;
  assign io_release_bits_data = R2;
  assign T3 = T6 ? T4 : R2;
  assign T4 = {io_data_resp, T5};
  assign T5 = R2[9'h1ff:8'h80];
  assign T6 = active & r2_data_req_fired;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = active ? r1_data_req_fired : r2_data_req_fired;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = T23 ? 1'h1 : T11;
  assign T11 = active ? 1'h0 : r1_data_req_fired;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T1 ? 1'h1 : T14;
  assign T14 = T16 ? T15 : active;
  assign T15 = io_release_ready ^ 1'h1;
  assign T16 = active & T17;
  assign T17 = T27 & T18;
  assign T18 = cnt == 3'h4;
  assign T19 = reset ? 3'h0 : T20;
  assign T20 = T1 ? 3'h0 : T21;
  assign T21 = T23 ? T22 : cnt;
  assign T22 = cnt + 3'h1;
  assign T23 = active & T24;
  assign T24 = T26 & T25;
  assign T25 = io_meta_read_ready & io_meta_read_valid;
  assign T26 = io_data_req_ready & io_data_req_valid;
  assign T27 = T29 & T28;
  assign T28 = r2_data_req_fired ^ 1'h1;
  assign T29 = r1_data_req_fired ^ 1'h1;
  assign io_release_bits_master_xact_id = req_master_xact_id;
  assign T30 = T1 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign T31 = T1 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_release_bits_addr = T32;
  assign T32 = T33;
  assign T33 = {req_tag, req_idx};
  assign T34 = T1 ? io_req_bits_idx : req_idx;
  assign T35 = T1 ? io_req_bits_tag : req_tag;
  assign io_release_valid = T16;
  assign io_data_req_bits_addr = T36;
  assign T36 = T37 << 3'h4;
  assign T37 = {req_idx, T38};
  assign T38 = cnt[1'h1:1'h0];
  assign io_data_req_bits_way_en = req_way_en;
  assign T39 = T1 ? io_req_bits_way_en : req_way_en;
  assign io_data_req_valid = fire;
  assign fire = active & T40;
  assign T40 = cnt < 3'h4;
  assign io_meta_read_bits_tag = req_tag;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_valid = fire;
  assign io_req_ready = T41;
  assign T41 = active ^ 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      req_r_type <= io_req_bits_r_type;
    end
    if(T6) begin
      R2 <= T4;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else if(active) begin
      r2_data_req_fired <= r1_data_req_fired;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else if(T23) begin
      r1_data_req_fired <= 1'h1;
    end else if(active) begin
      r1_data_req_fired <= 1'h0;
    end
    if(reset) begin
      active <= 1'h0;
    end else if(T1) begin
      active <= 1'h1;
    end else if(T16) begin
      active <= T15;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else if(T1) begin
      cnt <= 3'h0;
    end else if(T23) begin
      cnt <= T22;
    end
    if(T1) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T1) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T1) begin
      req_idx <= io_req_bits_idx;
    end
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      req_way_en <= io_req_bits_way_en;
    end
  end
endmodule

module ProbeUnit(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [25:0] io_req_bits_addr,
    input [2:0] io_req_bits_master_xact_id,
    input [1:0] io_req_bits_p_type,
    input [1:0] io_req_bits_client_xact_id,
    input  io_rep_ready,
    output io_rep_valid,
    output[25:0] io_rep_bits_addr,
    output[1:0] io_rep_bits_client_xact_id,
    output[2:0] io_rep_bits_master_xact_id,
    output[511:0] io_rep_bits_data,
    output[2:0] io_rep_bits_r_type,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    input  io_way_en,
    input  io_mshr_rdy,
    input [1:0] io_line_state_state
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire T4;
  reg [1:0] req_p_type;
  wire[1:0] T5;
  wire T6;
  wire T7;
  reg [3:0] state;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire[3:0] T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire[3:0] T28;
  wire T29;
  reg [1:0] line_state_state;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  reg  way_en;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire[2:0] T43;
  wire[2:0] T44;
  wire[2:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire[1:0] T51;
  reg [2:0] req_master_xact_id;
  wire[2:0] T52;
  reg [1:0] req_client_xact_id;
  wire[1:0] T53;
  wire[5:0] T54;
  reg [25:0] req_addr;
  wire[25:0] T55;
  wire[19:0] T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[19:0] T65;
  wire[5:0] T66;
  wire T67;
  wire[19:0] T68;
  wire[5:0] T69;
  wire T70;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire[2:0] T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[511:0] T88;
  wire[2:0] T89;
  wire[1:0] T90;
  wire[25:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_p_type = {1{$random}};
    state = {1{$random}};
    line_state_state = {1{$random}};
    way_en = {1{$random}};
    req_master_xact_id = {1{$random}};
    req_client_xact_id = {1{$random}};
    req_addr = {1{$random}};
  end
`endif

  assign io_wb_req_bits_r_type = T0;
  assign T0 = T49 ? T43 : T1;
  assign T1 = T42 ? 3'h4 : T2;
  assign T2 = T41 ? 3'h5 : T3;
  assign T3 = T4 ? 3'h6 : 3'h4;
  assign T4 = req_p_type == 2'h2;
  assign T5 = T6 ? io_req_bits_p_type : req_p_type;
  assign T6 = T7 & io_req_valid;
  assign T7 = state == 4'h1;
  assign T8 = reset ? 4'h1 : T9;
  assign T9 = T40 ? 4'h1 : T10;
  assign T10 = T6 ? 4'h2 : T11;
  assign T11 = T38 ? 4'h3 : T12;
  assign T12 = T37 ? 4'h4 : T13;
  assign T13 = T35 ? 4'h2 : T14;
  assign T14 = T31 ? 4'h5 : T15;
  assign T15 = T32 ? T28 : T16;
  assign T16 = T26 ? 4'h1 : T17;
  assign T17 = T24 ? 4'h7 : T18;
  assign T18 = T22 ? 4'h8 : T19;
  assign T19 = T20 ? 4'h1 : state;
  assign T20 = T21 & io_meta_write_ready;
  assign T21 = state == 4'h8;
  assign T22 = T23 & io_wb_req_ready;
  assign T23 = state == 4'h7;
  assign T24 = T25 & io_wb_req_ready;
  assign T25 = state == 4'h6;
  assign T26 = T27 & io_rep_ready;
  assign T27 = state == 4'h5;
  assign T28 = T29 ? 4'h6 : 4'h8;
  assign T29 = line_state_state == 2'h3;
  assign T30 = T31 ? io_line_state_state : line_state_state;
  assign T31 = state == 4'h4;
  assign T32 = T26 & T33;
  assign T33 = way_en != 1'h0;
  assign T34 = T31 ? io_way_en : way_en;
  assign T35 = T31 & T36;
  assign T36 = io_mshr_rdy ^ 1'h1;
  assign T37 = state == 4'h3;
  assign T38 = T39 & io_meta_read_ready;
  assign T39 = state == 4'h2;
  assign T40 = state == 4'h0;
  assign T41 = req_p_type == 2'h1;
  assign T42 = req_p_type == 2'h0;
  assign T43 = T48 ? 3'h1 : T44;
  assign T44 = T47 ? 3'h2 : T45;
  assign T45 = T46 ? 3'h3 : 3'h1;
  assign T46 = req_p_type == 2'h2;
  assign T47 = req_p_type == 2'h1;
  assign T48 = req_p_type == 2'h0;
  assign T49 = T50 == 2'h3;
  assign T50 = T33 ? line_state_state : T51;
  assign T51 = 2'h0;
  assign io_wb_req_bits_master_xact_id = req_master_xact_id;
  assign T52 = T6 ? io_req_bits_master_xact_id : req_master_xact_id;
  assign io_wb_req_bits_client_xact_id = req_client_xact_id;
  assign T53 = T6 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign io_wb_req_bits_way_en = way_en;
  assign io_wb_req_bits_idx = T54;
  assign T54 = req_addr[3'h5:1'h0];
  assign T55 = T6 ? io_req_bits_addr : req_addr;
  assign io_wb_req_bits_tag = T56;
  assign T56 = req_addr >> 3'h6;
  assign io_wb_req_valid = T57;
  assign T57 = state == 4'h6;
  assign io_meta_write_bits_data_coh_state = T58;
  assign T58 = T59;
  assign T59 = T64 ? 2'h0 : T60;
  assign T60 = T63 ? 2'h1 : T61;
  assign T61 = T62 ? line_state_state : line_state_state;
  assign T62 = req_p_type == 2'h2;
  assign T63 = req_p_type == 2'h1;
  assign T64 = req_p_type == 2'h0;
  assign io_meta_write_bits_data_tag = T65;
  assign T65 = req_addr >> 3'h6;
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_idx = T66;
  assign T66 = req_addr[3'h5:1'h0];
  assign io_meta_write_valid = T67;
  assign T67 = state == 4'h8;
  assign io_meta_read_bits_tag = T68;
  assign T68 = req_addr >> 3'h6;
  assign io_meta_read_bits_idx = T69;
  assign T69 = req_addr[3'h5:1'h0];
  assign io_meta_read_valid = T70;
  assign T70 = state == 4'h2;
  assign io_rep_bits_r_type = T71;
  assign T71 = T72;
  assign T72 = T85 ? T79 : T73;
  assign T73 = T78 ? 3'h4 : T74;
  assign T74 = T77 ? 3'h5 : T75;
  assign T75 = T76 ? 3'h6 : 3'h4;
  assign T76 = req_p_type == 2'h2;
  assign T77 = req_p_type == 2'h1;
  assign T78 = req_p_type == 2'h0;
  assign T79 = T84 ? 3'h1 : T80;
  assign T80 = T83 ? 3'h2 : T81;
  assign T81 = T82 ? 3'h3 : 3'h1;
  assign T82 = req_p_type == 2'h2;
  assign T83 = req_p_type == 2'h1;
  assign T84 = req_p_type == 2'h0;
  assign T85 = T86 == 2'h3;
  assign T86 = T33 ? line_state_state : T87;
  assign T87 = 2'h0;
  assign io_rep_bits_data = T88;
  assign T88 = 512'h0;
  assign io_rep_bits_master_xact_id = T89;
  assign T89 = req_master_xact_id;
  assign io_rep_bits_client_xact_id = T90;
  assign T90 = req_client_xact_id;
  assign io_rep_bits_addr = T91;
  assign T91 = req_addr;
  assign io_rep_valid = T92;
  assign T92 = T96 & T93;
  assign T93 = T94 ^ 1'h1;
  assign T94 = T33 & T95;
  assign T95 = line_state_state == 2'h3;
  assign T96 = state == 4'h5;
  assign io_req_ready = T97;
  assign T97 = state == 4'h1;

  always @(posedge clk) begin
    if(T6) begin
      req_p_type <= io_req_bits_p_type;
    end
    if(reset) begin
      state <= 4'h1;
    end else if(T40) begin
      state <= 4'h1;
    end else if(T6) begin
      state <= 4'h2;
    end else if(T38) begin
      state <= 4'h3;
    end else if(T37) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h2;
    end else if(T31) begin
      state <= 4'h5;
    end else if(T32) begin
      state <= T28;
    end else if(T26) begin
      state <= 4'h1;
    end else if(T24) begin
      state <= 4'h7;
    end else if(T22) begin
      state <= 4'h8;
    end else if(T20) begin
      state <= 4'h1;
    end
    if(T31) begin
      line_state_state <= io_line_state_state;
    end
    if(T31) begin
      way_en <= io_way_en;
    end
    if(T6) begin
      req_master_xact_id <= io_req_bits_master_xact_id;
    end
    if(T6) begin
      req_client_xact_id <= io_req_bits_client_xact_id;
    end
    if(T6) begin
      req_addr <= io_req_bits_addr;
    end
  end
endmodule

module Arbiter_0(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input [19:0] io_in_1_bits_tag,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input [19:0] io_in_0_bits_tag,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[19:0] io_out_bits_tag,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[19:0] T2;
  wire T3;
  wire[5:0] T4;
  wire T5;
  wire T6;
  wire T7;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_tag = T2;
  assign T2 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign T3 = T0;
  assign io_out_bits_idx = T4;
  assign T4 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T5;
  assign T5 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T6;
  assign T6 = T7 & io_out_ready;
  assign T7 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_1(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [19:0] io_in_1_bits_data_tag,
    input [1:0] io_in_1_bits_data_coh_state,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [19:0] io_in_0_bits_data_tag,
    input [1:0] io_in_0_bits_data_coh_state,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[19:0] io_out_bits_data_tag,
    output[1:0] io_out_bits_data_coh_state,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[1:0] T2;
  wire T3;
  wire[19:0] T4;
  wire T5;
  wire[5:0] T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data_coh_state = T2;
  assign T2 = T3 ? io_in_1_bits_data_coh_state : io_in_0_bits_data_coh_state;
  assign T3 = T0;
  assign io_out_bits_data_tag = T4;
  assign T4 = T3 ? io_in_1_bits_data_tag : io_in_0_bits_data_tag;
  assign io_out_bits_way_en = T5;
  assign T5 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T6;
  assign T6 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_2(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_a_type,
    input [5:0] io_in_1_bits_write_mask,
    input [2:0] io_in_1_bits_subword_addr,
    input [3:0] io_in_1_bits_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_a_type,
    input [5:0] io_in_0_bits_write_mask,
    input [2:0] io_in_0_bits_subword_addr,
    input [3:0] io_in_0_bits_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_a_type,
    output[5:0] io_out_bits_write_mask,
    output[2:0] io_out_bits_subword_addr,
    output[3:0] io_out_bits_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[3:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[2:0] T6;
  wire[511:0] T7;
  wire[1:0] T8;
  wire[25:0] T9;
  wire T10;
  wire T11;
  wire T12;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_atomic_opcode = T2;
  assign T2 = T3 ? io_in_1_bits_atomic_opcode : io_in_0_bits_atomic_opcode;
  assign T3 = T0;
  assign io_out_bits_subword_addr = T4;
  assign T4 = T3 ? io_in_1_bits_subword_addr : io_in_0_bits_subword_addr;
  assign io_out_bits_write_mask = T5;
  assign T5 = T3 ? io_in_1_bits_write_mask : io_in_0_bits_write_mask;
  assign io_out_bits_a_type = T6;
  assign T6 = T3 ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign io_out_bits_data = T7;
  assign T7 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_client_xact_id = T8;
  assign T8 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T9;
  assign T9 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T10;
  assign T10 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T11;
  assign T11 = T12 & io_out_ready;
  assign T12 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_3(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire T6;
  wire T7;
  wire T8;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_payload_master_xact_id = T2;
  assign T2 = T3 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T3 = T0;
  assign io_out_bits_header_dst = T4;
  assign T4 = T3 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T5;
  assign T5 = T3 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T6;
  assign T6 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T7;
  assign T7 = T8 & io_out_ready;
  assign T8 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_4(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [19:0] io_in_1_bits_tag,
    input [5:0] io_in_1_bits_idx,
    input  io_in_1_bits_way_en,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [19:0] io_in_0_bits_tag,
    input [5:0] io_in_0_bits_idx,
    input  io_in_0_bits_way_en,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[19:0] io_out_bits_tag,
    output[5:0] io_out_bits_idx,
    output io_out_bits_way_en,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[2:0] T4;
  wire[1:0] T5;
  wire T6;
  wire[5:0] T7;
  wire[19:0] T8;
  wire T9;
  wire T10;
  wire T11;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_master_xact_id = T4;
  assign T4 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_bits_idx = T7;
  assign T7 = T3 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign io_out_bits_tag = T8;
  assign T8 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_valid = T9;
  assign T9 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T10;
  assign T10 = T11 & io_out_ready;
  assign T11 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_5(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_kill,
    input [2:0] io_in_1_bits_typ,
    input  io_in_1_bits_phys,
    input [43:0] io_in_1_bits_addr,
    input [63:0] io_in_1_bits_data,
    input [7:0] io_in_1_bits_tag,
    input [4:0] io_in_1_bits_cmd,
    input [4:0] io_in_1_bits_sdq_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_kill,
    input [2:0] io_in_0_bits_typ,
    input  io_in_0_bits_phys,
    input [43:0] io_in_0_bits_addr,
    input [63:0] io_in_0_bits_data,
    input [7:0] io_in_0_bits_tag,
    input [4:0] io_in_0_bits_cmd,
    input [4:0] io_in_0_bits_sdq_id,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_kill,
    output[2:0] io_out_bits_typ,
    output io_out_bits_phys,
    output[43:0] io_out_bits_addr,
    output[63:0] io_out_bits_data,
    output[7:0] io_out_bits_tag,
    output[4:0] io_out_bits_cmd,
    output[4:0] io_out_bits_sdq_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[4:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[7:0] T5;
  wire[63:0] T6;
  wire[43:0] T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_sdq_id = T2;
  assign T2 = T3 ? io_in_1_bits_sdq_id : io_in_0_bits_sdq_id;
  assign T3 = T0;
  assign io_out_bits_cmd = T4;
  assign T4 = T3 ? io_in_1_bits_cmd : io_in_0_bits_cmd;
  assign io_out_bits_tag = T5;
  assign T5 = T3 ? io_in_1_bits_tag : io_in_0_bits_tag;
  assign io_out_bits_data = T6;
  assign T6 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_phys = T8;
  assign T8 = T3 ? io_in_1_bits_phys : io_in_0_bits_phys;
  assign io_out_bits_typ = T9;
  assign T9 = T3 ? io_in_1_bits_typ : io_in_0_bits_typ;
  assign io_out_bits_kill = T10;
  assign T10 = T3 ? io_in_1_bits_kill : io_in_0_bits_kill;
  assign io_out_valid = T11;
  assign T11 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = io_in_0_valid ^ 1'h1;
endmodule

module Arbiter_6(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits = T2;
  assign T2 = T3 ? io_in_1_bits : io_in_0_bits;
  assign T3 = T0;
  assign io_out_valid = T4;
  assign T4 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T5;
  assign T5 = T6 & io_out_ready;
  assign T6 = io_in_0_valid ^ 1'h1;
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_kill,
    input [2:0] io_enq_bits_typ,
    input  io_enq_bits_phys,
    input [43:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input [7:0] io_enq_bits_tag,
    input [4:0] io_enq_bits_cmd,
    input [4:0] io_enq_bits_sdq_id,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_kill,
    output[2:0] io_deq_bits_typ,
    output io_deq_bits_phys,
    output[43:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data,
    output[7:0] io_deq_bits_tag,
    output[4:0] io_deq_bits_cmd,
    output[4:0] io_deq_bits_sdq_id,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire do_deq;
  reg [3:0] R5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire do_enq;
  wire T9;
  wire ptr_match;
  reg  maybe_full;
  wire T10;
  wire T11;
  wire T12;
  wire[4:0] T13;
  wire[130:0] T14;
  reg [130:0] ram [15:0];
  wire[130:0] T15;
  wire[130:0] T16;
  wire[130:0] T17;
  wire[81:0] T18;
  wire[9:0] T19;
  wire[71:0] T20;
  wire[48:0] T21;
  wire[44:0] T22;
  wire[3:0] T23;
  wire[4:0] T24;
  wire[7:0] T25;
  wire[63:0] T26;
  wire[43:0] T27;
  wire T28;
  wire[2:0] T29;
  wire T30;
  wire T31;
  wire empty;
  wire T32;
  wire T33;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {5{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T9, ptr_diff};
  assign ptr_diff = R5 - R1;
  assign T2 = reset ? 4'h0 : T3;
  assign T3 = do_deq ? T4 : R1;
  assign T4 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 4'h0 : T7;
  assign T7 = do_enq ? T8 : R5;
  assign T8 = R5 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T9 = maybe_full & ptr_match;
  assign ptr_match = R5 == R1;
  assign T10 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign io_deq_bits_sdq_id = T13;
  assign T13 = T14[3'h4:1'h0];
  assign T14 = ram[R1];
  assign T16 = T17;
  assign T17 = {T21, T18};
  assign T18 = {T20, T19};
  assign T19 = {io_enq_bits_cmd, io_enq_bits_sdq_id};
  assign T20 = {io_enq_bits_data, io_enq_bits_tag};
  assign T21 = {T23, T22};
  assign T22 = {io_enq_bits_phys, io_enq_bits_addr};
  assign T23 = {io_enq_bits_kill, io_enq_bits_typ};
  assign io_deq_bits_cmd = T24;
  assign T24 = T14[4'h9:3'h5];
  assign io_deq_bits_tag = T25;
  assign T25 = T14[5'h11:4'ha];
  assign io_deq_bits_data = T26;
  assign T26 = T14[7'h51:5'h12];
  assign io_deq_bits_addr = T27;
  assign T27 = T14[7'h7d:7'h52];
  assign io_deq_bits_phys = T28;
  assign T28 = T14[7'h7e:7'h7e];
  assign io_deq_bits_typ = T29;
  assign T29 = T14[8'h81:7'h7f];
  assign io_deq_bits_kill = T30;
  assign T30 = T14[8'h82:8'h82];
  assign io_deq_valid = T31;
  assign T31 = empty ^ 1'h1;
  assign empty = ptr_match & T32;
  assign T32 = maybe_full ^ 1'h1;
  assign io_enq_ready = T33;
  assign T33 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T4;
    end
    if(reset) begin
      R5 <= 4'h0;
    end else if(do_enq) begin
      R5 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R5] <= T16;
  end
endmodule

module MSHR_0(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire rpq_io_deq_valid;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  reg [1:0] refill_count;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire reply;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire idx_match;
  wire[5:0] T125;
  wire[5:0] T126;
  reg [43:0] req_addr;
  wire[43:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg [1:0] meta_hazard;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg  req_way_en;
  wire T144;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T145;
  wire T146;
  wire ackq_io_enq_ready;
  wire T147;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire T148;
  wire ackq_io_deq_valid;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire[4:0] T149;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[63:0] rpq_io_deq_bits_data;
  wire[43:0] T150;
  wire[31:0] T151;
  wire[31:0] T152;
  wire[11:0] T153;
  wire[5:0] T154;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire T155;
  wire T156;
  wire[1:0] T157;
  reg [1:0] line_state_state;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T161;
  wire[1:0] T162;
  wire[1:0] T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] meta_on_flush_state;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[127:0] T182;
  reg [63:0] req_data;
  wire[63:0] T183;
  wire[11:0] T184;
  wire[7:0] T185;
  reg [2:0] acquire_type;
  wire[2:0] T186;
  wire[2:0] T187;
  wire[2:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire[2:0] T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[25:0] T213;
  wire[25:0] T214;
  wire T215;
  wire T216;
  wire[19:0] T217;
  wire[31:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire rpq_io_enq_ready;
  wire T222;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T63 | T1;
  assign T1 = state == 4'h5;
  assign T2 = reset ? 4'h0 : T3;
  assign T3 = T61 ? T59 : T4;
  assign T4 = T57 ? 4'h4 : T5;
  assign T5 = T35 ? 4'h6 : T6;
  assign T6 = T34 ? 4'h2 : T7;
  assign T7 = T32 ? 4'h3 : T8;
  assign T8 = T30 ? 4'h4 : T9;
  assign T9 = T29 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T27 & refill_done;
  assign refill_done = reply & T21;
  assign T21 = refill_count == 2'h3;
  assign T22 = T28 ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_count;
  assign T24 = refill_count + 2'h1;
  assign T25 = T27 & reply;
  assign reply = io_mem_grant_valid & T26;
  assign T26 = io_mem_grant_bits_payload_client_xact_id == 2'h0;
  assign T27 = state == 4'h5;
  assign T28 = io_req_pri_val & io_req_pri_rdy;
  assign T29 = io_mem_req_ready & io_mem_req_valid;
  assign T30 = T31 & io_meta_write_ready;
  assign T31 = state == 4'h3;
  assign T32 = T33 & reply;
  assign T33 = state == 4'h2;
  assign T34 = io_wb_req_ready & io_wb_req_valid;
  assign T35 = T56 & T36;
  assign T36 = T45 ? T42 : T37;
  assign T37 = T39 | T38;
  assign T38 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T39 = T41 | T40;
  assign T40 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T42 = T44 | T43;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T44 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T45 = T47 | T46;
  assign T46 = io_req_bits_cmd == 5'h6;
  assign T47 = T49 | T48;
  assign T48 = io_req_bits_cmd == 5'h3;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h4;
  assign T52 = io_req_bits_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h7;
  assign T55 = io_req_bits_cmd == 5'h1;
  assign T56 = T28 & io_req_bits_tag_match;
  assign T57 = T56 & T58;
  assign T58 = T36 ^ 1'h1;
  assign T59 = T60 ? 4'h1 : 4'h3;
  assign T60 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T61 = T28 & T62;
  assign T62 = io_req_bits_tag_match ^ 1'h1;
  assign T63 = T65 | T64;
  assign T64 = state == 4'h4;
  assign T65 = state == 4'h0;
  assign T66 = T68 & T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T128 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T120 | T84;
  assign T84 = T117 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 3'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T110 & T101;
  assign T101 = T103 | T102;
  assign T102 = 3'h6 == io_mem_req_bits_a_type;
  assign T103 = T105 | T104;
  assign T104 = 3'h5 == io_mem_req_bits_a_type;
  assign T105 = T107 | T106;
  assign T106 = 3'h4 == io_mem_req_bits_a_type;
  assign T107 = T109 | T108;
  assign T108 = 3'h3 == io_mem_req_bits_a_type;
  assign T109 = 3'h2 == io_mem_req_bits_a_type;
  assign T110 = T114 | T111;
  assign T111 = T113 | T112;
  assign T112 = io_req_bits_cmd == 5'h4;
  assign T113 = io_req_bits_cmd[2'h3:2'h3];
  assign T114 = T116 | T115;
  assign T115 = io_req_bits_cmd == 5'h6;
  assign T116 = io_req_bits_cmd == 5'h0;
  assign T117 = T119 | T118;
  assign T118 = state == 4'h5;
  assign T119 = state == 4'h4;
  assign T120 = T122 | T121;
  assign T121 = state == 4'h3;
  assign T122 = T124 | T123;
  assign T123 = state == 4'h2;
  assign T124 = state == 4'h1;
  assign idx_match = T126 == T125;
  assign T125 = io_req_bits_addr[4'hb:3'h6];
  assign T126 = req_addr[4'hb:3'h6];
  assign T127 = T28 ? io_req_bits_addr : req_addr;
  assign T128 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T129;
  assign T129 = T143 | T130;
  assign T130 = T138 & T131;
  assign T131 = meta_hazard == 2'h0;
  assign T132 = reset ? 2'h0 : T133;
  assign T133 = T137 ? 2'h1 : T134;
  assign T134 = T136 ? T135 : meta_hazard;
  assign T135 = meta_hazard + 2'h1;
  assign T136 = meta_hazard != 2'h0;
  assign T137 = io_meta_write_ready & io_meta_write_valid;
  assign T138 = T140 & T139;
  assign T139 = state != 4'h3;
  assign T140 = T142 & T141;
  assign T141 = state != 4'h2;
  assign T142 = state != 4'h1;
  assign T143 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h0;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T144 = T28 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = T126;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T145 = T28 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T146;
  assign T146 = T147 & ackq_io_enq_ready;
  assign T147 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T148;
  assign T148 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T149;
  assign T149 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T150;
  assign T150 = {12'h0, T151};
  assign T151 = T152;
  assign T152 = {io_tag, T153};
  assign T153 = {T126, T154};
  assign T154 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T155;
  assign T155 = T156 & rpq_io_deq_valid;
  assign T156 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T157;
  assign T157 = T177 ? meta_on_flush_state : line_state_state;
  assign T158 = T35 ? meta_on_hit_state : T159;
  assign T159 = T28 ? meta_on_flush_state : T160;
  assign T160 = T25 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T161;
  assign T161 = T168 ? 2'h1 : T162;
  assign T162 = T167 ? T165 : T163;
  assign T163 = T164 ? 2'h3 : 2'h0;
  assign T164 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T165 = T166 ? 2'h3 : 2'h2;
  assign T166 = io_mem_req_bits_a_type == 3'h1;
  assign T167 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T168 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_flush_state = 2'h0;
  assign meta_on_hit_state = T169;
  assign T169 = T170 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T170 = T174 | T171;
  assign T171 = T173 | T172;
  assign T172 = io_req_bits_cmd == 5'h4;
  assign T173 = io_req_bits_cmd[2'h3:2'h3];
  assign T174 = T176 | T175;
  assign T175 = io_req_bits_cmd == 5'h7;
  assign T176 = io_req_bits_cmd == 5'h1;
  assign T177 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = T126;
  assign io_meta_write_valid = T178;
  assign T178 = T180 | T179;
  assign T179 = state == 4'h3;
  assign T180 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = T126;
  assign io_meta_read_valid = T181;
  assign T181 = state == 4'h8;
  assign io_mem_resp_data = T182;
  assign T182 = {64'h0, req_data};
  assign T183 = T28 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T184;
  assign T184 = T185 << 3'h4;
  assign T185 = {T126, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T186 = T28 ? T201 : T187;
  assign T187 = T200 ? T188 : acquire_type;
  assign T188 = T189 ? 3'h1 : io_mem_req_bits_a_type;
  assign T189 = T191 | T190;
  assign T190 = io_req_bits_cmd == 5'h6;
  assign T191 = T193 | T192;
  assign T192 = io_req_bits_cmd == 5'h3;
  assign T193 = T197 | T194;
  assign T194 = T196 | T195;
  assign T195 = io_req_bits_cmd == 5'h4;
  assign T196 = io_req_bits_cmd[2'h3:2'h3];
  assign T197 = T199 | T198;
  assign T198 = io_req_bits_cmd == 5'h7;
  assign T199 = io_req_bits_cmd == 5'h1;
  assign T200 = io_req_sec_val & io_req_sec_rdy;
  assign T201 = T202 ? 3'h1 : 3'h0;
  assign T202 = T204 | T203;
  assign T203 = io_req_bits_cmd == 5'h6;
  assign T204 = T206 | T205;
  assign T205 = io_req_bits_cmd == 5'h3;
  assign T206 = T210 | T207;
  assign T207 = T209 | T208;
  assign T208 = io_req_bits_cmd == 5'h4;
  assign T209 = io_req_bits_cmd[2'h3:2'h3];
  assign T210 = T212 | T211;
  assign T211 = io_req_bits_cmd == 5'h7;
  assign T212 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h0;
  assign io_mem_req_bits_addr = T213;
  assign T213 = T214;
  assign T214 = {io_tag, T126};
  assign io_mem_req_valid = T215;
  assign T215 = T216 & ackq_io_enq_ready;
  assign T216 = state == 4'h4;
  assign io_tag = T217;
  assign T217 = T218[5'h13:1'h0];
  assign T218 = req_addr >> 4'hc;
  assign io_idx_match = T219;
  assign T219 = T220 & idx_match;
  assign T220 = state != 4'h0;
  assign io_req_sec_rdy = T221;
  assign T221 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T222;
  assign T222 = state == 4'h0;
  Queue_1 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_0 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T66 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T61) begin
      state <= T59;
    end else if(T57) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h6;
    end else if(T34) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h3;
    end else if(T30) begin
      state <= 4'h4;
    end else if(T29) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(T28) begin
      refill_count <= 2'h0;
    end else if(T25) begin
      refill_count <= T24;
    end
    if(T28) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T137) begin
      meta_hazard <= 2'h1;
    end else if(T136) begin
      meta_hazard <= T135;
    end
    if(T28) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T28) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T35) begin
      line_state_state <= meta_on_hit_state;
    end else if(T28) begin
      line_state_state <= meta_on_flush_state;
    end else if(T25) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T28) begin
      req_data <= io_req_bits_data;
    end
    if(T28) begin
      acquire_type <= T201;
    end else if(T200) begin
      acquire_type <= T188;
    end
  end
endmodule

module MSHR_1(input clk, input reset,
    input  io_req_pri_val,
    output io_req_pri_rdy,
    input  io_req_sec_val,
    output io_req_sec_rdy,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    input [4:0] io_req_sdq_id,
    output io_idx_match,
    output[19:0] io_tag,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    //output[511:0] io_mem_req_bits_data
    output[2:0] io_mem_req_bits_a_type,
    //output[5:0] io_mem_req_bits_write_mask
    //output[2:0] io_mem_req_bits_subword_addr
    //output[3:0] io_mem_req_bits_atomic_opcode
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy
);

  wire T0;
  wire can_finish;
  wire T1;
  reg [3:0] state;
  wire[3:0] T2;
  wire[3:0] T3;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[3:0] T6;
  wire[3:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire rpq_io_deq_valid;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire refill_done;
  wire T21;
  reg [1:0] refill_count;
  wire[1:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire reply;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire[3:0] T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire wb_done;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire sec_rdy;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire idx_match;
  wire[5:0] T125;
  wire[5:0] T126;
  reg [43:0] req_addr;
  wire[43:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg [1:0] meta_hazard;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg  req_way_en;
  wire T144;
  reg [19:0] req_old_meta_tag;
  wire[19:0] T145;
  wire T146;
  wire ackq_io_enq_ready;
  wire T147;
  wire[2:0] ackq_io_deq_bits_payload_master_xact_id;
  wire[1:0] ackq_io_deq_bits_header_dst;
  wire[1:0] ackq_io_deq_bits_header_src;
  wire T148;
  wire ackq_io_deq_valid;
  wire[4:0] rpq_io_deq_bits_sdq_id;
  wire[4:0] T149;
  wire[4:0] rpq_io_deq_bits_cmd;
  wire[7:0] rpq_io_deq_bits_tag;
  wire[63:0] rpq_io_deq_bits_data;
  wire[43:0] T150;
  wire[31:0] T151;
  wire[31:0] T152;
  wire[11:0] T153;
  wire[5:0] T154;
  wire[43:0] rpq_io_deq_bits_addr;
  wire[2:0] rpq_io_deq_bits_typ;
  wire rpq_io_deq_bits_kill;
  wire T155;
  wire T156;
  wire[1:0] T157;
  reg [1:0] line_state_state;
  wire[1:0] T158;
  wire[1:0] T159;
  wire[1:0] T160;
  wire[1:0] meta_on_grant_state;
  wire[1:0] T161;
  wire[1:0] T162;
  wire[1:0] T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[1:0] meta_on_flush_state;
  wire[1:0] meta_on_hit_state;
  wire[1:0] T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire[127:0] T182;
  reg [63:0] req_data;
  wire[63:0] T183;
  wire[11:0] T184;
  wire[7:0] T185;
  reg [2:0] acquire_type;
  wire[2:0] T186;
  wire[2:0] T187;
  wire[2:0] T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire[2:0] T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire[25:0] T213;
  wire[25:0] T214;
  wire T215;
  wire T216;
  wire[19:0] T217;
  wire[31:0] T218;
  wire T219;
  wire T220;
  wire T221;
  wire rpq_io_enq_ready;
  wire T222;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    refill_count = {1{$random}};
    req_addr = {2{$random}};
    meta_hazard = {1{$random}};
    req_way_en = {1{$random}};
    req_old_meta_tag = {1{$random}};
    line_state_state = {1{$random}};
    req_data = {2{$random}};
    acquire_type = {1{$random}};
  end
`endif

  assign T0 = io_mem_finish_ready & can_finish;
  assign can_finish = T63 | T1;
  assign T1 = state == 4'h5;
  assign T2 = reset ? 4'h0 : T3;
  assign T3 = T61 ? T59 : T4;
  assign T4 = T57 ? 4'h4 : T5;
  assign T5 = T35 ? 4'h6 : T6;
  assign T6 = T34 ? 4'h2 : T7;
  assign T7 = T32 ? 4'h3 : T8;
  assign T8 = T30 ? 4'h4 : T9;
  assign T9 = T29 ? 4'h5 : T10;
  assign T10 = T20 ? 4'h6 : T11;
  assign T11 = T18 ? 4'h7 : T12;
  assign T12 = T17 ? 4'h8 : T13;
  assign T13 = T14 ? 4'h0 : state;
  assign T14 = T16 & T15;
  assign T15 = rpq_io_deq_valid ^ 1'h1;
  assign T16 = state == 4'h8;
  assign T17 = state == 4'h7;
  assign T18 = T19 & io_meta_write_ready;
  assign T19 = state == 4'h6;
  assign T20 = T27 & refill_done;
  assign refill_done = reply & T21;
  assign T21 = refill_count == 2'h3;
  assign T22 = T28 ? 2'h0 : T23;
  assign T23 = T25 ? T24 : refill_count;
  assign T24 = refill_count + 2'h1;
  assign T25 = T27 & reply;
  assign reply = io_mem_grant_valid & T26;
  assign T26 = io_mem_grant_bits_payload_client_xact_id == 2'h1;
  assign T27 = state == 4'h5;
  assign T28 = io_req_pri_val & io_req_pri_rdy;
  assign T29 = io_mem_req_ready & io_mem_req_valid;
  assign T30 = T31 & io_meta_write_ready;
  assign T31 = state == 4'h3;
  assign T32 = T33 & reply;
  assign T33 = state == 4'h2;
  assign T34 = io_wb_req_ready & io_wb_req_valid;
  assign T35 = T56 & T36;
  assign T36 = T45 ? T42 : T37;
  assign T37 = T39 | T38;
  assign T38 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T39 = T41 | T40;
  assign T40 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T41 = io_req_bits_old_meta_coh_state == 2'h1;
  assign T42 = T44 | T43;
  assign T43 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T44 = io_req_bits_old_meta_coh_state == 2'h2;
  assign T45 = T47 | T46;
  assign T46 = io_req_bits_cmd == 5'h6;
  assign T47 = T49 | T48;
  assign T48 = io_req_bits_cmd == 5'h3;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = io_req_bits_cmd == 5'h4;
  assign T52 = io_req_bits_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = io_req_bits_cmd == 5'h7;
  assign T55 = io_req_bits_cmd == 5'h1;
  assign T56 = T28 & io_req_bits_tag_match;
  assign T57 = T56 & T58;
  assign T58 = T36 ^ 1'h1;
  assign T59 = T60 ? 4'h1 : 4'h3;
  assign T60 = io_req_bits_old_meta_coh_state == 2'h3;
  assign T61 = T28 & T62;
  assign T62 = io_req_bits_tag_match ^ 1'h1;
  assign T63 = T65 | T64;
  assign T64 = state == 4'h4;
  assign T65 = state == 4'h0;
  assign T66 = T68 & T67;
  assign T67 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T68 = wb_done | refill_done;
  assign wb_done = reply & T69;
  assign T69 = state == 4'h2;
  assign T70 = T75 ? 1'h0 : T71;
  assign T71 = T73 | T72;
  assign T72 = state == 4'h0;
  assign T73 = io_replay_ready & T74;
  assign T74 = state == 4'h8;
  assign T75 = io_meta_read_ready ^ 1'h1;
  assign T76 = T81 & T77;
  assign T77 = T78 ^ 1'h1;
  assign T78 = T80 | T79;
  assign T79 = io_req_bits_cmd == 5'h3;
  assign T80 = io_req_bits_cmd == 5'h2;
  assign T81 = T128 | T82;
  assign T82 = io_req_sec_val & sec_rdy;
  assign sec_rdy = idx_match & T83;
  assign T83 = T120 | T84;
  assign T84 = T117 & T85;
  assign T85 = T86 ^ 1'h1;
  assign T86 = T100 | T87;
  assign T87 = T89 & T88;
  assign T88 = io_mem_req_bits_a_type != 3'h1;
  assign T89 = T91 | T90;
  assign T90 = io_req_bits_cmd == 5'h6;
  assign T91 = T93 | T92;
  assign T92 = io_req_bits_cmd == 5'h3;
  assign T93 = T97 | T94;
  assign T94 = T96 | T95;
  assign T95 = io_req_bits_cmd == 5'h4;
  assign T96 = io_req_bits_cmd[2'h3:2'h3];
  assign T97 = T99 | T98;
  assign T98 = io_req_bits_cmd == 5'h7;
  assign T99 = io_req_bits_cmd == 5'h1;
  assign T100 = T110 & T101;
  assign T101 = T103 | T102;
  assign T102 = 3'h6 == io_mem_req_bits_a_type;
  assign T103 = T105 | T104;
  assign T104 = 3'h5 == io_mem_req_bits_a_type;
  assign T105 = T107 | T106;
  assign T106 = 3'h4 == io_mem_req_bits_a_type;
  assign T107 = T109 | T108;
  assign T108 = 3'h3 == io_mem_req_bits_a_type;
  assign T109 = 3'h2 == io_mem_req_bits_a_type;
  assign T110 = T114 | T111;
  assign T111 = T113 | T112;
  assign T112 = io_req_bits_cmd == 5'h4;
  assign T113 = io_req_bits_cmd[2'h3:2'h3];
  assign T114 = T116 | T115;
  assign T115 = io_req_bits_cmd == 5'h6;
  assign T116 = io_req_bits_cmd == 5'h0;
  assign T117 = T119 | T118;
  assign T118 = state == 4'h5;
  assign T119 = state == 4'h4;
  assign T120 = T122 | T121;
  assign T121 = state == 4'h3;
  assign T122 = T124 | T123;
  assign T123 = state == 4'h2;
  assign T124 = state == 4'h1;
  assign idx_match = T126 == T125;
  assign T125 = io_req_bits_addr[4'hb:3'h6];
  assign T126 = req_addr[4'hb:3'h6];
  assign T127 = T28 ? io_req_bits_addr : req_addr;
  assign T128 = io_req_pri_val & io_req_pri_rdy;
  assign io_probe_rdy = T129;
  assign T129 = T143 | T130;
  assign T130 = T138 & T131;
  assign T131 = meta_hazard == 2'h0;
  assign T132 = reset ? 2'h0 : T133;
  assign T133 = T137 ? 2'h1 : T134;
  assign T134 = T136 ? T135 : meta_hazard;
  assign T135 = meta_hazard + 2'h1;
  assign T136 = meta_hazard != 2'h0;
  assign T137 = io_meta_write_ready & io_meta_write_valid;
  assign T138 = T140 & T139;
  assign T139 = state != 4'h3;
  assign T140 = T142 & T141;
  assign T141 = state != 4'h2;
  assign T142 = state != 4'h1;
  assign T143 = idx_match ^ 1'h1;
  assign io_wb_req_bits_r_type = 3'h0;
  assign io_wb_req_bits_master_xact_id = 3'h0;
  assign io_wb_req_bits_client_xact_id = 2'h1;
  assign io_wb_req_bits_way_en = req_way_en;
  assign T144 = T28 ? io_req_bits_way_en : req_way_en;
  assign io_wb_req_bits_idx = T126;
  assign io_wb_req_bits_tag = req_old_meta_tag;
  assign T145 = T28 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign io_wb_req_valid = T146;
  assign T146 = T147 & ackq_io_enq_ready;
  assign T147 = state == 4'h1;
  assign io_mem_finish_bits_payload_master_xact_id = ackq_io_deq_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = ackq_io_deq_bits_header_dst;
  assign io_mem_finish_bits_header_src = ackq_io_deq_bits_header_src;
  assign io_mem_finish_valid = T148;
  assign T148 = ackq_io_deq_valid & can_finish;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_replay_bits_cmd = T149;
  assign T149 = T75 ? 5'h5 : rpq_io_deq_bits_cmd;
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_data = rpq_io_deq_bits_data;
  assign io_replay_bits_addr = T150;
  assign T150 = {12'h0, T151};
  assign T151 = T152;
  assign T152 = {io_tag, T153};
  assign T153 = {T126, T154};
  assign T154 = rpq_io_deq_bits_addr[3'h5:1'h0];
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_kill = rpq_io_deq_bits_kill;
  assign io_replay_valid = T155;
  assign T155 = T156 & rpq_io_deq_valid;
  assign T156 = state == 4'h8;
  assign io_meta_write_bits_data_coh_state = T157;
  assign T157 = T177 ? meta_on_flush_state : line_state_state;
  assign T158 = T35 ? meta_on_hit_state : T159;
  assign T159 = T28 ? meta_on_flush_state : T160;
  assign T160 = T25 ? meta_on_grant_state : line_state_state;
  assign meta_on_grant_state = T161;
  assign T161 = T168 ? 2'h1 : T162;
  assign T162 = T167 ? T165 : T163;
  assign T163 = T164 ? 2'h3 : 2'h0;
  assign T164 = io_mem_grant_bits_payload_g_type == 4'h5;
  assign T165 = T166 ? 2'h3 : 2'h2;
  assign T166 = io_mem_req_bits_a_type == 3'h1;
  assign T167 = io_mem_grant_bits_payload_g_type == 4'h2;
  assign T168 = io_mem_grant_bits_payload_g_type == 4'h1;
  assign meta_on_flush_state = 2'h0;
  assign meta_on_hit_state = T169;
  assign T169 = T170 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign T170 = T174 | T171;
  assign T171 = T173 | T172;
  assign T172 = io_req_bits_cmd == 5'h4;
  assign T173 = io_req_bits_cmd[2'h3:2'h3];
  assign T174 = T176 | T175;
  assign T175 = io_req_bits_cmd == 5'h7;
  assign T176 = io_req_bits_cmd == 5'h1;
  assign T177 = state == 4'h3;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_idx = T126;
  assign io_meta_write_valid = T178;
  assign T178 = T180 | T179;
  assign T179 = state == 4'h3;
  assign T180 = state == 4'h6;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_read_bits_idx = T126;
  assign io_meta_read_valid = T181;
  assign T181 = state == 4'h8;
  assign io_mem_resp_data = T182;
  assign T182 = {64'h0, req_data};
  assign T183 = T28 ? io_req_bits_data : req_data;
  assign io_mem_resp_addr = T184;
  assign T184 = T185 << 3'h4;
  assign T185 = {T126, refill_count};
  assign io_mem_resp_way_en = req_way_en;
  assign io_mem_req_bits_a_type = acquire_type;
  assign T186 = T28 ? T201 : T187;
  assign T187 = T200 ? T188 : acquire_type;
  assign T188 = T189 ? 3'h1 : io_mem_req_bits_a_type;
  assign T189 = T191 | T190;
  assign T190 = io_req_bits_cmd == 5'h6;
  assign T191 = T193 | T192;
  assign T192 = io_req_bits_cmd == 5'h3;
  assign T193 = T197 | T194;
  assign T194 = T196 | T195;
  assign T195 = io_req_bits_cmd == 5'h4;
  assign T196 = io_req_bits_cmd[2'h3:2'h3];
  assign T197 = T199 | T198;
  assign T198 = io_req_bits_cmd == 5'h7;
  assign T199 = io_req_bits_cmd == 5'h1;
  assign T200 = io_req_sec_val & io_req_sec_rdy;
  assign T201 = T202 ? 3'h1 : 3'h0;
  assign T202 = T204 | T203;
  assign T203 = io_req_bits_cmd == 5'h6;
  assign T204 = T206 | T205;
  assign T205 = io_req_bits_cmd == 5'h3;
  assign T206 = T210 | T207;
  assign T207 = T209 | T208;
  assign T208 = io_req_bits_cmd == 5'h4;
  assign T209 = io_req_bits_cmd[2'h3:2'h3];
  assign T210 = T212 | T211;
  assign T211 = io_req_bits_cmd == 5'h7;
  assign T212 = io_req_bits_cmd == 5'h1;
  assign io_mem_req_bits_client_xact_id = 2'h1;
  assign io_mem_req_bits_addr = T213;
  assign T213 = T214;
  assign T214 = {io_tag, T126};
  assign io_mem_req_valid = T215;
  assign T215 = T216 & ackq_io_enq_ready;
  assign T216 = state == 4'h4;
  assign io_tag = T217;
  assign T217 = T218[5'h13:1'h0];
  assign T218 = req_addr >> 4'hc;
  assign io_idx_match = T219;
  assign T219 = T220 & idx_match;
  assign T220 = state != 4'h0;
  assign io_req_sec_rdy = T221;
  assign T221 = sec_rdy & rpq_io_enq_ready;
  assign io_req_pri_rdy = T222;
  assign T222 = state == 4'h0;
  Queue_1 rpq(.clk(clk), .reset(reset),
       .io_enq_ready( rpq_io_enq_ready ),
       .io_enq_valid( T76 ),
       .io_enq_bits_kill( io_req_bits_kill ),
       .io_enq_bits_typ( io_req_bits_typ ),
       .io_enq_bits_phys( io_req_bits_phys ),
       .io_enq_bits_addr( io_req_bits_addr ),
       .io_enq_bits_data( io_req_bits_data ),
       .io_enq_bits_tag( io_req_bits_tag ),
       .io_enq_bits_cmd( io_req_bits_cmd ),
       .io_enq_bits_sdq_id( io_req_sdq_id ),
       .io_deq_ready( T70 ),
       .io_deq_valid( rpq_io_deq_valid ),
       .io_deq_bits_kill( rpq_io_deq_bits_kill ),
       .io_deq_bits_typ( rpq_io_deq_bits_typ ),
       //.io_deq_bits_phys(  )
       .io_deq_bits_addr( rpq_io_deq_bits_addr ),
       .io_deq_bits_data( rpq_io_deq_bits_data ),
       .io_deq_bits_tag( rpq_io_deq_bits_tag ),
       .io_deq_bits_cmd( rpq_io_deq_bits_cmd ),
       .io_deq_bits_sdq_id( rpq_io_deq_bits_sdq_id )
       //.io_count(  )
  );
  Queue_0 ackq(.clk(clk), .reset(reset),
       .io_enq_ready( ackq_io_enq_ready ),
       .io_enq_valid( T66 ),
       //.io_enq_bits_header_src(  )
       .io_enq_bits_header_dst( io_mem_grant_bits_header_src ),
       .io_enq_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_deq_ready( T0 ),
       .io_deq_valid( ackq_io_deq_valid ),
       .io_deq_bits_header_src( ackq_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( ackq_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( ackq_io_deq_bits_payload_master_xact_id )
       //.io_count(  )
  );
  `ifndef SYNTHESIS
    assign ackq.io_enq_bits_header_src = {1{$random}};
  `endif

  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else if(T61) begin
      state <= T59;
    end else if(T57) begin
      state <= 4'h4;
    end else if(T35) begin
      state <= 4'h6;
    end else if(T34) begin
      state <= 4'h2;
    end else if(T32) begin
      state <= 4'h3;
    end else if(T30) begin
      state <= 4'h4;
    end else if(T29) begin
      state <= 4'h5;
    end else if(T20) begin
      state <= 4'h6;
    end else if(T18) begin
      state <= 4'h7;
    end else if(T17) begin
      state <= 4'h8;
    end else if(T14) begin
      state <= 4'h0;
    end
    if(T28) begin
      refill_count <= 2'h0;
    end else if(T25) begin
      refill_count <= T24;
    end
    if(T28) begin
      req_addr <= io_req_bits_addr;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else if(T137) begin
      meta_hazard <= 2'h1;
    end else if(T136) begin
      meta_hazard <= T135;
    end
    if(T28) begin
      req_way_en <= io_req_bits_way_en;
    end
    if(T28) begin
      req_old_meta_tag <= io_req_bits_old_meta_tag;
    end
    if(T35) begin
      line_state_state <= meta_on_hit_state;
    end else if(T28) begin
      line_state_state <= meta_on_flush_state;
    end else if(T25) begin
      line_state_state <= meta_on_grant_state;
    end
    if(T28) begin
      req_data <= io_req_bits_data;
    end
    if(T28) begin
      acquire_type <= T201;
    end else if(T200) begin
      acquire_type <= T188;
    end
  end
endmodule

module MSHRFile(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input  io_req_bits_kill,
    input [2:0] io_req_bits_typ,
    input  io_req_bits_phys,
    input [43:0] io_req_bits_addr,
    input [63:0] io_req_bits_data,
    input [7:0] io_req_bits_tag,
    input [4:0] io_req_bits_cmd,
    input  io_req_bits_tag_match,
    input [19:0] io_req_bits_old_meta_tag,
    input [1:0] io_req_bits_old_meta_coh_state,
    input  io_req_bits_way_en,
    output io_secondary_miss,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output[25:0] io_mem_req_bits_addr,
    output[1:0] io_mem_req_bits_client_xact_id,
    output[511:0] io_mem_req_bits_data,
    output[2:0] io_mem_req_bits_a_type,
    output[5:0] io_mem_req_bits_write_mask,
    output[2:0] io_mem_req_bits_subword_addr,
    output[3:0] io_mem_req_bits_atomic_opcode,
    output io_mem_resp_way_en,
    output[11:0] io_mem_resp_addr,
    output[1:0] io_mem_resp_wmask,
    output[127:0] io_mem_resp_data,
    input  io_meta_read_ready,
    output io_meta_read_valid,
    output[5:0] io_meta_read_bits_idx,
    output[19:0] io_meta_read_bits_tag,
    input  io_meta_write_ready,
    output io_meta_write_valid,
    output[5:0] io_meta_write_bits_idx,
    output io_meta_write_bits_way_en,
    output[19:0] io_meta_write_bits_data_tag,
    output[1:0] io_meta_write_bits_data_coh_state,
    input  io_replay_ready,
    output io_replay_valid,
    output io_replay_bits_kill,
    output[2:0] io_replay_bits_typ,
    output io_replay_bits_phys,
    output[43:0] io_replay_bits_addr,
    output[63:0] io_replay_bits_data,
    output[7:0] io_replay_bits_tag,
    output[4:0] io_replay_bits_cmd,
    output[4:0] io_replay_bits_sdq_id,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    input  io_wb_req_ready,
    output io_wb_req_valid,
    output[19:0] io_wb_req_bits_tag,
    output[5:0] io_wb_req_bits_idx,
    output io_wb_req_bits_way_en,
    output[1:0] io_wb_req_bits_client_xact_id,
    output[2:0] io_wb_req_bits_master_xact_id,
    output[2:0] io_wb_req_bits_r_type,
    output io_probe_rdy,
    output io_fence_rdy
);

  wire wb_req_arb_io_in_1_ready;
  wire mem_finish_arb_io_in_1_ready;
  wire replay_arb_io_in_1_ready;
  wire meta_write_arb_io_in_1_ready;
  wire meta_read_arb_io_in_1_ready;
  wire mem_req_arb_io_in_1_ready;
  wire[4:0] T0;
  wire[4:0] T1;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[4:0] T7;
  wire[4:0] T8;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[4:0] T11;
  wire[4:0] T12;
  wire[4:0] T13;
  wire[4:0] T14;
  wire[4:0] T15;
  wire T16;
  wire[16:0] T17;
  wire[16:0] T18;
  reg [16:0] sdq_val;
  wire[16:0] T19;
  wire[31:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[31:0] T23;
  wire[31:0] T24;
  wire[16:0] T25;
  wire[16:0] T26;
  wire[16:0] T27;
  wire sdq_enq;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire[16:0] T36;
  wire[16:0] T37;
  wire[16:0] T38;
  wire[16:0] T39;
  wire[16:0] T40;
  wire[16:0] T41;
  wire[16:0] T42;
  wire[16:0] T43;
  wire[16:0] T44;
  wire[16:0] T45;
  wire[16:0] T46;
  wire[16:0] T47;
  wire[16:0] T48;
  wire[16:0] T49;
  wire[16:0] T50;
  wire[16:0] T51;
  wire[16:0] T52;
  wire T53;
  wire[16:0] T54;
  wire[16:0] T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire[31:0] T72;
  wire[31:0] T73;
  wire[31:0] T74;
  wire[31:0] T75;
  wire[16:0] T76;
  wire[16:0] T77;
  wire free_sdq;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire[31:0] T86;
  wire[31:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire tag_match;
  wire[31:0] T105;
  wire[31:0] T106;
  wire[19:0] T107;
  wire[19:0] T108;
  wire[19:0] tagList_1;
  wire[19:0] MSHR_1_io_tag;
  wire idxMatch_1;
  wire MSHR_1_io_idx_match;
  wire[19:0] T109;
  wire[19:0] tagList_0;
  wire[19:0] MSHR_0_io_tag;
  wire idxMatch_0;
  wire MSHR_0_io_idx_match;
  wire T110;
  wire sdq_rdy;
  wire T111;
  wire alloc_arb_io_in_1_ready;
  wire wb_req_arb_io_in_0_ready;
  wire mem_finish_arb_io_in_0_ready;
  wire replay_arb_io_in_0_ready;
  wire meta_write_arb_io_in_0_ready;
  wire meta_read_arb_io_in_0_ready;
  wire mem_req_arb_io_in_0_ready;
  wire T112;
  wire T113;
  wire alloc_arb_io_in_0_ready;
  wire T114;
  wire T115;
  wire idx_match;
  wire T116;
  wire MSHR_0_io_req_pri_rdy;
  wire MSHR_1_io_req_pri_rdy;
  wire[4:0] MSHR_0_io_replay_bits_sdq_id;
  wire[4:0] MSHR_0_io_replay_bits_cmd;
  wire[7:0] MSHR_0_io_replay_bits_tag;
  wire[63:0] MSHR_0_io_replay_bits_data;
  wire[43:0] MSHR_0_io_replay_bits_addr;
  wire MSHR_0_io_replay_bits_phys;
  wire[2:0] MSHR_0_io_replay_bits_typ;
  wire MSHR_0_io_replay_bits_kill;
  wire MSHR_0_io_replay_valid;
  wire[4:0] MSHR_1_io_replay_bits_sdq_id;
  wire[4:0] MSHR_1_io_replay_bits_cmd;
  wire[7:0] MSHR_1_io_replay_bits_tag;
  wire[63:0] MSHR_1_io_replay_bits_data;
  wire[43:0] MSHR_1_io_replay_bits_addr;
  wire MSHR_1_io_replay_bits_phys;
  wire[2:0] MSHR_1_io_replay_bits_typ;
  wire MSHR_1_io_replay_bits_kill;
  wire MSHR_1_io_replay_valid;
  wire[2:0] MSHR_0_io_wb_req_bits_r_type;
  wire[2:0] MSHR_0_io_wb_req_bits_master_xact_id;
  wire[1:0] MSHR_0_io_wb_req_bits_client_xact_id;
  wire MSHR_0_io_wb_req_bits_way_en;
  wire[5:0] MSHR_0_io_wb_req_bits_idx;
  wire[19:0] MSHR_0_io_wb_req_bits_tag;
  wire MSHR_0_io_wb_req_valid;
  wire[2:0] MSHR_1_io_wb_req_bits_r_type;
  wire[2:0] MSHR_1_io_wb_req_bits_master_xact_id;
  wire[1:0] MSHR_1_io_wb_req_bits_client_xact_id;
  wire MSHR_1_io_wb_req_bits_way_en;
  wire[5:0] MSHR_1_io_wb_req_bits_idx;
  wire[19:0] MSHR_1_io_wb_req_bits_tag;
  wire MSHR_1_io_wb_req_valid;
  wire[2:0] MSHR_0_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_dst;
  wire[1:0] MSHR_0_io_mem_finish_bits_header_src;
  wire MSHR_0_io_mem_finish_valid;
  wire[2:0] MSHR_1_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_dst;
  wire[1:0] MSHR_1_io_mem_finish_bits_header_src;
  wire MSHR_1_io_mem_finish_valid;
  wire[2:0] MSHR_0_io_mem_req_bits_a_type;
  wire[1:0] MSHR_0_io_mem_req_bits_client_xact_id;
  wire[25:0] MSHR_0_io_mem_req_bits_addr;
  wire MSHR_0_io_mem_req_valid;
  wire[2:0] MSHR_1_io_mem_req_bits_a_type;
  wire[1:0] MSHR_1_io_mem_req_bits_client_xact_id;
  wire[25:0] MSHR_1_io_mem_req_bits_addr;
  wire MSHR_1_io_mem_req_valid;
  wire[1:0] MSHR_0_io_meta_write_bits_data_coh_state;
  wire[19:0] MSHR_0_io_meta_write_bits_data_tag;
  wire MSHR_0_io_meta_write_bits_way_en;
  wire[5:0] MSHR_0_io_meta_write_bits_idx;
  wire MSHR_0_io_meta_write_valid;
  wire[1:0] MSHR_1_io_meta_write_bits_data_coh_state;
  wire[19:0] MSHR_1_io_meta_write_bits_data_tag;
  wire MSHR_1_io_meta_write_bits_way_en;
  wire[5:0] MSHR_1_io_meta_write_bits_idx;
  wire MSHR_1_io_meta_write_valid;
  wire[19:0] MSHR_0_io_meta_read_bits_tag;
  wire[5:0] MSHR_0_io_meta_read_bits_idx;
  wire MSHR_0_io_meta_read_valid;
  wire[19:0] MSHR_1_io_meta_read_bits_tag;
  wire[5:0] MSHR_1_io_meta_read_bits_idx;
  wire MSHR_1_io_meta_read_valid;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire MSHR_0_io_probe_rdy;
  wire T124;
  wire MSHR_1_io_probe_rdy;
  wire[2:0] wb_req_arb_io_out_bits_r_type;
  wire[2:0] wb_req_arb_io_out_bits_master_xact_id;
  wire[1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire wb_req_arb_io_out_bits_way_en;
  wire[5:0] wb_req_arb_io_out_bits_idx;
  wire[19:0] wb_req_arb_io_out_bits_tag;
  wire wb_req_arb_io_out_valid;
  wire[2:0] mem_finish_arb_io_out_bits_payload_master_xact_id;
  wire[1:0] mem_finish_arb_io_out_bits_header_dst;
  wire[1:0] mem_finish_arb_io_out_bits_header_src;
  wire mem_finish_arb_io_out_valid;
  wire[4:0] replay_arb_io_out_bits_sdq_id;
  wire[4:0] replay_arb_io_out_bits_cmd;
  wire[7:0] replay_arb_io_out_bits_tag;
  wire[63:0] T125;
  reg [63:0] sdq [16:0];
  wire[63:0] T126;
  wire T127;
  wire T128;
  wire[4:0] T129;
  reg [4:0] R130;
  wire[4:0] T131;
  wire[43:0] replay_arb_io_out_bits_addr;
  wire replay_arb_io_out_bits_phys;
  wire[2:0] replay_arb_io_out_bits_typ;
  wire replay_arb_io_out_bits_kill;
  wire replay_arb_io_out_valid;
  wire[1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire[19:0] meta_write_arb_io_out_bits_data_tag;
  wire meta_write_arb_io_out_bits_way_en;
  wire[5:0] meta_write_arb_io_out_bits_idx;
  wire meta_write_arb_io_out_valid;
  wire[19:0] meta_read_arb_io_out_bits_tag;
  wire[5:0] meta_read_arb_io_out_bits_idx;
  wire meta_read_arb_io_out_valid;
  wire[127:0] T132;
  wire[127:0] memRespMux_0_data;
  wire[127:0] MSHR_0_io_mem_resp_data;
  wire[127:0] memRespMux_1_data;
  wire[127:0] MSHR_1_io_mem_resp_data;
  wire T133;
  wire T134;
  wire[1:0] T135;
  wire[1:0] memRespMux_0_wmask;
  wire[1:0] MSHR_0_io_mem_resp_wmask;
  wire[1:0] memRespMux_1_wmask;
  wire[1:0] MSHR_1_io_mem_resp_wmask;
  wire[11:0] T136;
  wire[11:0] memRespMux_0_addr;
  wire[11:0] MSHR_0_io_mem_resp_addr;
  wire[11:0] memRespMux_1_addr;
  wire[11:0] MSHR_1_io_mem_resp_addr;
  wire T137;
  wire memRespMux_0_way_en;
  wire MSHR_0_io_mem_resp_way_en;
  wire memRespMux_1_way_en;
  wire MSHR_1_io_mem_resp_way_en;
  wire[3:0] mem_req_arb_io_out_bits_atomic_opcode;
  wire[2:0] mem_req_arb_io_out_bits_subword_addr;
  wire[5:0] mem_req_arb_io_out_bits_write_mask;
  wire[2:0] mem_req_arb_io_out_bits_a_type;
  wire[511:0] mem_req_arb_io_out_bits_data;
  wire[1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire[25:0] mem_req_arb_io_out_bits_addr;
  wire mem_req_arb_io_out_valid;
  wire T138;
  wire T139;
  wire pri_rdy;
  wire T140;
  wire sec_rdy;
  wire MSHR_1_io_req_sec_rdy;
  wire MSHR_0_io_req_sec_rdy;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    sdq_val = {1{$random}};
    for (initvar = 0; initvar < 17; initvar = initvar+1)
      sdq[initvar] = {2{$random}};
    R130 = {1{$random}};
  end
`endif

  assign T0 = T103 ? 1'h0 : T1;
  assign T1 = T102 ? 1'h1 : T2;
  assign T2 = T101 ? 2'h2 : T3;
  assign T3 = T100 ? 2'h3 : T4;
  assign T4 = T99 ? 3'h4 : T5;
  assign T5 = T98 ? 3'h5 : T6;
  assign T6 = T97 ? 3'h6 : T7;
  assign T7 = T96 ? 3'h7 : T8;
  assign T8 = T95 ? 4'h8 : T9;
  assign T9 = T94 ? 4'h9 : T10;
  assign T10 = T93 ? 4'ha : T11;
  assign T11 = T92 ? 4'hb : T12;
  assign T12 = T91 ? 4'hc : T13;
  assign T13 = T90 ? 4'hd : T14;
  assign T14 = T89 ? 4'he : T15;
  assign T15 = T16 ? 4'hf : 5'h10;
  assign T16 = T17[4'hf:4'hf];
  assign T17 = ~ T18;
  assign T18 = sdq_val[5'h10:1'h0];
  assign T19 = T20[5'h10:1'h0];
  assign T20 = reset ? 32'h0 : T21;
  assign T21 = T88 ? T23 : T22;
  assign T22 = {15'h0, sdq_val};
  assign T23 = T72 | T24;
  assign T24 = {15'h0, T25};
  assign T25 = T36 & T26;
  assign T26 = 17'h0 - T27;
  assign T27 = {16'h0, sdq_enq};
  assign sdq_enq = T35 & T28;
  assign T28 = T32 | T29;
  assign T29 = T31 | T30;
  assign T30 = io_req_bits_cmd == 5'h4;
  assign T31 = io_req_bits_cmd[2'h3:2'h3];
  assign T32 = T34 | T33;
  assign T33 = io_req_bits_cmd == 5'h7;
  assign T34 = io_req_bits_cmd == 5'h1;
  assign T35 = io_req_valid & io_req_ready;
  assign T36 = T71 ? 17'h1 : T37;
  assign T37 = T70 ? 17'h2 : T38;
  assign T38 = T69 ? 17'h4 : T39;
  assign T39 = T68 ? 17'h8 : T40;
  assign T40 = T67 ? 17'h10 : T41;
  assign T41 = T66 ? 17'h20 : T42;
  assign T42 = T65 ? 17'h40 : T43;
  assign T43 = T64 ? 17'h80 : T44;
  assign T44 = T63 ? 17'h100 : T45;
  assign T45 = T62 ? 17'h200 : T46;
  assign T46 = T61 ? 17'h400 : T47;
  assign T47 = T60 ? 17'h800 : T48;
  assign T48 = T59 ? 17'h1000 : T49;
  assign T49 = T58 ? 17'h2000 : T50;
  assign T50 = T57 ? 17'h4000 : T51;
  assign T51 = T56 ? 17'h8000 : T52;
  assign T52 = T53 ? 17'h10000 : 17'h0;
  assign T53 = T54[5'h10:5'h10];
  assign T54 = ~ T55;
  assign T55 = sdq_val[5'h10:1'h0];
  assign T56 = T54[4'hf:4'hf];
  assign T57 = T54[4'he:4'he];
  assign T58 = T54[4'hd:4'hd];
  assign T59 = T54[4'hc:4'hc];
  assign T60 = T54[4'hb:4'hb];
  assign T61 = T54[4'ha:4'ha];
  assign T62 = T54[4'h9:4'h9];
  assign T63 = T54[4'h8:4'h8];
  assign T64 = T54[3'h7:3'h7];
  assign T65 = T54[3'h6:3'h6];
  assign T66 = T54[3'h5:3'h5];
  assign T67 = T54[3'h4:3'h4];
  assign T68 = T54[2'h3:2'h3];
  assign T69 = T54[2'h2:2'h2];
  assign T70 = T54[1'h1:1'h1];
  assign T71 = T54[1'h0:1'h0];
  assign T72 = T87 & T73;
  assign T73 = ~ T74;
  assign T74 = T86 & T75;
  assign T75 = {15'h0, T76};
  assign T76 = 17'h0 - T77;
  assign T77 = {16'h0, free_sdq};
  assign free_sdq = T85 & T78;
  assign T78 = T82 | T79;
  assign T79 = T81 | T80;
  assign T80 = io_replay_bits_cmd == 5'h4;
  assign T81 = io_replay_bits_cmd[2'h3:2'h3];
  assign T82 = T84 | T83;
  assign T83 = io_replay_bits_cmd == 5'h7;
  assign T84 = io_replay_bits_cmd == 5'h1;
  assign T85 = io_replay_ready & io_replay_valid;
  assign T86 = 1'h1 << io_replay_bits_sdq_id;
  assign T87 = {15'h0, sdq_val};
  assign T88 = io_replay_valid | sdq_enq;
  assign T89 = T17[4'he:4'he];
  assign T90 = T17[4'hd:4'hd];
  assign T91 = T17[4'hc:4'hc];
  assign T92 = T17[4'hb:4'hb];
  assign T93 = T17[4'ha:4'ha];
  assign T94 = T17[4'h9:4'h9];
  assign T95 = T17[4'h8:4'h8];
  assign T96 = T17[3'h7:3'h7];
  assign T97 = T17[3'h6:3'h6];
  assign T98 = T17[3'h5:3'h5];
  assign T99 = T17[3'h4:3'h4];
  assign T100 = T17[2'h3:2'h3];
  assign T101 = T17[2'h2:2'h2];
  assign T102 = T17[1'h1:1'h1];
  assign T103 = T17[1'h0:1'h0];
  assign T104 = T110 & tag_match;
  assign tag_match = T106 == T105;
  assign T105 = io_req_bits_addr >> 4'hc;
  assign T106 = {12'h0, T107};
  assign T107 = T109 | T108;
  assign T108 = idxMatch_1 ? tagList_1 : 20'h0;
  assign tagList_1 = MSHR_1_io_tag;
  assign idxMatch_1 = MSHR_1_io_idx_match;
  assign T109 = idxMatch_0 ? tagList_0 : 20'h0;
  assign tagList_0 = MSHR_0_io_tag;
  assign idxMatch_0 = MSHR_0_io_idx_match;
  assign T110 = io_req_valid & sdq_rdy;
  assign sdq_rdy = T111 ^ 1'h1;
  assign T111 = sdq_val == 17'h1ffff;
  assign T112 = T113 & tag_match;
  assign T113 = io_req_valid & sdq_rdy;
  assign T114 = T116 & T115;
  assign T115 = idx_match ^ 1'h1;
  assign idx_match = MSHR_0_io_idx_match | MSHR_1_io_idx_match;
  assign T116 = io_req_valid & sdq_rdy;
  assign io_fence_rdy = T117;
  assign T117 = T120 ? 1'h0 : T118;
  assign T118 = T119 == 1'h0;
  assign T119 = MSHR_0_io_req_pri_rdy ^ 1'h1;
  assign T120 = MSHR_1_io_req_pri_rdy ^ 1'h1;
  assign io_probe_rdy = T121;
  assign T121 = T124 ? 1'h0 : T122;
  assign T122 = T123 == 1'h0;
  assign T123 = MSHR_0_io_probe_rdy ^ 1'h1;
  assign T124 = MSHR_1_io_probe_rdy ^ 1'h1;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_master_xact_id = wb_req_arb_io_out_bits_master_xact_id;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_wb_req_bits_idx = wb_req_arb_io_out_bits_idx;
  assign io_wb_req_bits_tag = wb_req_arb_io_out_bits_tag;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_mem_finish_bits_payload_master_xact_id = mem_finish_arb_io_out_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mem_finish_arb_io_out_bits_header_dst;
  assign io_mem_finish_bits_header_src = mem_finish_arb_io_out_bits_header_src;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_replay_bits_sdq_id = replay_arb_io_out_bits_sdq_id;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_data = T125;
  assign T125 = sdq[R130];
  assign T127 = sdq_enq & T128;
  assign T128 = T129 < 5'h11;
  assign T129 = T0[3'h4:1'h0];
  assign T131 = free_sdq ? replay_arb_io_out_bits_sdq_id : R130;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_kill = replay_arb_io_out_bits_kill;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_mem_resp_data = T132;
  assign T132 = T133 ? memRespMux_1_data : memRespMux_0_data;
  assign memRespMux_0_data = MSHR_0_io_mem_resp_data;
  assign memRespMux_1_data = MSHR_1_io_mem_resp_data;
  assign T133 = T134;
  assign T134 = io_mem_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_mem_resp_wmask = T135;
  assign T135 = T133 ? memRespMux_1_wmask : memRespMux_0_wmask;
  assign memRespMux_0_wmask = MSHR_0_io_mem_resp_wmask;
  assign memRespMux_1_wmask = MSHR_1_io_mem_resp_wmask;
  assign io_mem_resp_addr = T136;
  assign T136 = T133 ? memRespMux_1_addr : memRespMux_0_addr;
  assign memRespMux_0_addr = MSHR_0_io_mem_resp_addr;
  assign memRespMux_1_addr = MSHR_1_io_mem_resp_addr;
  assign io_mem_resp_way_en = T137;
  assign T137 = T133 ? memRespMux_1_way_en : memRespMux_0_way_en;
  assign memRespMux_0_way_en = MSHR_0_io_mem_resp_way_en;
  assign memRespMux_1_way_en = MSHR_1_io_mem_resp_way_en;
  assign io_mem_req_bits_atomic_opcode = mem_req_arb_io_out_bits_atomic_opcode;
  assign io_mem_req_bits_subword_addr = mem_req_arb_io_out_bits_subword_addr;
  assign io_mem_req_bits_write_mask = mem_req_arb_io_out_bits_write_mask;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr = mem_req_arb_io_out_bits_addr;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_secondary_miss = idx_match;
  assign io_req_ready = T138;
  assign T138 = T139 & sdq_rdy;
  assign T139 = idx_match ? T140 : pri_rdy;
  assign pri_rdy = MSHR_0_io_req_pri_rdy | MSHR_1_io_req_pri_rdy;
  assign T140 = tag_match & sec_rdy;
  assign sec_rdy = MSHR_0_io_req_sec_rdy | MSHR_1_io_req_sec_rdy;
  Arbiter_0 meta_read_arb(
       .io_in_1_ready( meta_read_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_read_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_in_1_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_in_0_ready( meta_read_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_read_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_in_0_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_out_ready( io_meta_read_ready ),
       .io_out_valid( meta_read_arb_io_out_valid ),
       .io_out_bits_idx( meta_read_arb_io_out_bits_idx ),
       .io_out_bits_tag( meta_read_arb_io_out_bits_tag )
       //.io_chosen(  )
  );
  Arbiter_1 meta_write_arb(
       .io_in_1_ready( meta_write_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_meta_write_valid ),
       .io_in_1_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( meta_write_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_meta_write_valid ),
       .io_in_0_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_out_ready( io_meta_write_ready ),
       .io_out_valid( meta_write_arb_io_out_valid ),
       .io_out_bits_idx( meta_write_arb_io_out_bits_idx ),
       .io_out_bits_way_en( meta_write_arb_io_out_bits_way_en ),
       .io_out_bits_data_tag( meta_write_arb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( meta_write_arb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  Arbiter_2 mem_req_arb(
       .io_in_1_ready( mem_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_req_valid ),
       .io_in_1_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_in_1_bits_data(  )
       .io_in_1_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_in_1_bits_write_mask(  )
       //.io_in_1_bits_subword_addr(  )
       //.io_in_1_bits_atomic_opcode(  )
       .io_in_0_ready( mem_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_req_valid ),
       .io_in_0_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_in_0_bits_data(  )
       .io_in_0_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_in_0_bits_write_mask(  )
       //.io_in_0_bits_subword_addr(  )
       //.io_in_0_bits_atomic_opcode(  )
       .io_out_ready( io_mem_req_ready ),
       .io_out_valid( mem_req_arb_io_out_valid ),
       .io_out_bits_addr( mem_req_arb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( mem_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_data( mem_req_arb_io_out_bits_data ),
       .io_out_bits_a_type( mem_req_arb_io_out_bits_a_type ),
       .io_out_bits_write_mask( mem_req_arb_io_out_bits_write_mask ),
       .io_out_bits_subword_addr( mem_req_arb_io_out_bits_subword_addr ),
       .io_out_bits_atomic_opcode( mem_req_arb_io_out_bits_atomic_opcode )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign mem_req_arb.io_in_1_bits_data = {16{$random}};
    assign mem_req_arb.io_in_1_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_1_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_1_bits_atomic_opcode = {1{$random}};
    assign mem_req_arb.io_in_0_bits_data = {16{$random}};
    assign mem_req_arb.io_in_0_bits_write_mask = {1{$random}};
    assign mem_req_arb.io_in_0_bits_subword_addr = {1{$random}};
    assign mem_req_arb.io_in_0_bits_atomic_opcode = {1{$random}};
  `endif
  Arbiter_3 mem_finish_arb(
       .io_in_1_ready( mem_finish_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_mem_finish_valid ),
       .io_in_1_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_in_1_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( mem_finish_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_mem_finish_valid ),
       .io_in_0_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_in_0_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_mem_finish_ready ),
       .io_out_valid( mem_finish_arb_io_out_valid ),
       .io_out_bits_header_src( mem_finish_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( mem_finish_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( mem_finish_arb_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  Arbiter_4 wb_req_arb(
       .io_in_1_ready( wb_req_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_wb_req_valid ),
       .io_in_1_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_in_0_ready( wb_req_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_wb_req_valid ),
       .io_in_0_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_out_ready( io_wb_req_ready ),
       .io_out_valid( wb_req_arb_io_out_valid ),
       .io_out_bits_tag( wb_req_arb_io_out_bits_tag ),
       .io_out_bits_idx( wb_req_arb_io_out_bits_idx ),
       .io_out_bits_way_en( wb_req_arb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wb_req_arb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wb_req_arb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wb_req_arb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  Arbiter_5 replay_arb(
       .io_in_1_ready( replay_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_replay_valid ),
       .io_in_1_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_in_1_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_in_1_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_in_1_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_in_1_bits_data( MSHR_1_io_replay_bits_data ),
       .io_in_1_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_in_1_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_in_1_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_in_0_ready( replay_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_replay_valid ),
       .io_in_0_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_in_0_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_in_0_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_in_0_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_in_0_bits_data( MSHR_0_io_replay_bits_data ),
       .io_in_0_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_in_0_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_in_0_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_out_ready( io_replay_ready ),
       .io_out_valid( replay_arb_io_out_valid ),
       .io_out_bits_kill( replay_arb_io_out_bits_kill ),
       .io_out_bits_typ( replay_arb_io_out_bits_typ ),
       .io_out_bits_phys( replay_arb_io_out_bits_phys ),
       .io_out_bits_addr( replay_arb_io_out_bits_addr ),
       //.io_out_bits_data(  )
       .io_out_bits_tag( replay_arb_io_out_bits_tag ),
       .io_out_bits_cmd( replay_arb_io_out_bits_cmd ),
       .io_out_bits_sdq_id( replay_arb_io_out_bits_sdq_id )
       //.io_chosen(  )
  );
  Arbiter_6 alloc_arb(
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( MSHR_1_io_req_pri_rdy ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( MSHR_0_io_req_pri_rdy ),
       //.io_in_0_bits(  )
       .io_out_ready( T114 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  MSHR_0 MSHR_0(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_0_ready ),
       .io_req_pri_rdy( MSHR_0_io_req_pri_rdy ),
       .io_req_sec_val( T112 ),
       .io_req_sec_rdy( MSHR_0_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T0 ),
       .io_idx_match( MSHR_0_io_idx_match ),
       .io_tag( MSHR_0_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_0_ready ),
       .io_mem_req_valid( MSHR_0_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_0_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_0_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_0_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_0_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_0_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_0_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_0_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_0_ready ),
       .io_meta_read_valid( MSHR_0_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_0_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_0_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_0_ready ),
       .io_meta_write_valid( MSHR_0_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_0_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_0_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_0_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_0_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_0_ready ),
       .io_replay_valid( MSHR_0_io_replay_valid ),
       .io_replay_bits_kill( MSHR_0_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_0_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_0_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_0_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_0_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_0_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_0_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_0_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_0_ready ),
       .io_mem_finish_valid( MSHR_0_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_0_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_0_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_0_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_0_ready ),
       .io_wb_req_valid( MSHR_0_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_0_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_0_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_0_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_0_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_0_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_0_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_0_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_0.io_mem_resp_wmask = {1{$random}};
  `endif
  MSHR_1 MSHR_1(.clk(clk), .reset(reset),
       .io_req_pri_val( alloc_arb_io_in_1_ready ),
       .io_req_pri_rdy( MSHR_1_io_req_pri_rdy ),
       .io_req_sec_val( T104 ),
       .io_req_sec_rdy( MSHR_1_io_req_sec_rdy ),
       .io_req_bits_kill( io_req_bits_kill ),
       .io_req_bits_typ( io_req_bits_typ ),
       .io_req_bits_phys( io_req_bits_phys ),
       .io_req_bits_addr( io_req_bits_addr ),
       .io_req_bits_data( io_req_bits_data ),
       .io_req_bits_tag( io_req_bits_tag ),
       .io_req_bits_cmd( io_req_bits_cmd ),
       .io_req_bits_tag_match( io_req_bits_tag_match ),
       .io_req_bits_old_meta_tag( io_req_bits_old_meta_tag ),
       .io_req_bits_old_meta_coh_state( io_req_bits_old_meta_coh_state ),
       .io_req_bits_way_en( io_req_bits_way_en ),
       .io_req_sdq_id( T0 ),
       .io_idx_match( MSHR_1_io_idx_match ),
       .io_tag( MSHR_1_io_tag ),
       .io_mem_req_ready( mem_req_arb_io_in_1_ready ),
       .io_mem_req_valid( MSHR_1_io_mem_req_valid ),
       .io_mem_req_bits_addr( MSHR_1_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( MSHR_1_io_mem_req_bits_client_xact_id ),
       //.io_mem_req_bits_data(  )
       .io_mem_req_bits_a_type( MSHR_1_io_mem_req_bits_a_type ),
       //.io_mem_req_bits_write_mask(  )
       //.io_mem_req_bits_subword_addr(  )
       //.io_mem_req_bits_atomic_opcode(  )
       .io_mem_resp_way_en( MSHR_1_io_mem_resp_way_en ),
       .io_mem_resp_addr( MSHR_1_io_mem_resp_addr ),
       .io_mem_resp_wmask( MSHR_1_io_mem_resp_wmask ),
       .io_mem_resp_data( MSHR_1_io_mem_resp_data ),
       .io_meta_read_ready( meta_read_arb_io_in_1_ready ),
       .io_meta_read_valid( MSHR_1_io_meta_read_valid ),
       .io_meta_read_bits_idx( MSHR_1_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( MSHR_1_io_meta_read_bits_tag ),
       .io_meta_write_ready( meta_write_arb_io_in_1_ready ),
       .io_meta_write_valid( MSHR_1_io_meta_write_valid ),
       .io_meta_write_bits_idx( MSHR_1_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( MSHR_1_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( MSHR_1_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( MSHR_1_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( replay_arb_io_in_1_ready ),
       .io_replay_valid( MSHR_1_io_replay_valid ),
       .io_replay_bits_kill( MSHR_1_io_replay_bits_kill ),
       .io_replay_bits_typ( MSHR_1_io_replay_bits_typ ),
       .io_replay_bits_phys( MSHR_1_io_replay_bits_phys ),
       .io_replay_bits_addr( MSHR_1_io_replay_bits_addr ),
       .io_replay_bits_data( MSHR_1_io_replay_bits_data ),
       .io_replay_bits_tag( MSHR_1_io_replay_bits_tag ),
       .io_replay_bits_cmd( MSHR_1_io_replay_bits_cmd ),
       .io_replay_bits_sdq_id( MSHR_1_io_replay_bits_sdq_id ),
       .io_mem_grant_valid( io_mem_grant_valid ),
       .io_mem_grant_bits_header_src( io_mem_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_mem_finish_ready( mem_finish_arb_io_in_1_ready ),
       .io_mem_finish_valid( MSHR_1_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( MSHR_1_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( MSHR_1_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( MSHR_1_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wb_req_arb_io_in_1_ready ),
       .io_wb_req_valid( MSHR_1_io_wb_req_valid ),
       .io_wb_req_bits_tag( MSHR_1_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( MSHR_1_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( MSHR_1_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( MSHR_1_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( MSHR_1_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( MSHR_1_io_wb_req_bits_r_type ),
       .io_probe_rdy( MSHR_1_io_probe_rdy )
  );
  `ifndef SYNTHESIS
    assign MSHR_1.io_mem_resp_wmask = {1{$random}};
  `endif

  always @(posedge clk) begin
    sdq_val <= T19;
    if (T127)
      sdq[T0] <= io_req_bits_data;
    if(free_sdq) begin
      R130 <= replay_arb_io_out_bits_sdq_id;
    end
  end
endmodule

module MetadataArray(input clk, input reset,
    output io_read_ready,
    input  io_read_valid,
    input [5:0] io_read_bits_idx,
    output io_write_ready,
    input  io_write_valid,
    input [5:0] io_write_bits_idx,
    input  io_write_bits_way_en,
    input [19:0] io_write_bits_data_tag,
    input [1:0] io_write_bits_data_coh_state,
    output[19:0] io_resp_0_tag,
    output[1:0] io_resp_0_coh_state
);

  wire[1:0] T0;
  wire[21:0] T1;
  wire[21:0] T2;
  wire[21:0] T3;
  wire[21:0] T4;
  wire[21:0] T5;
  wire[21:0] T6;
  wire T7;
  wire wmask;
  wire T8;
  reg [6:0] rst_cnt;
  wire[6:0] T9;
  wire[6:0] T10;
  wire[6:0] T11;
  wire[21:0] wdata;
  wire[21:0] T12;
  wire[1:0] T13;
  wire[1:0] rstVal_coh_state;
  wire[1:0] T14;
  wire[19:0] T15;
  wire[19:0] rstVal_tag;
  wire T16;
  wire[5:0] T17;
  wire[6:0] waddr;
  wire[6:0] T18;
  reg [5:0] R19;
  wire[5:0] T20;
  wire[19:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    rst_cnt = {1{$random}};
    R19 = {1{$random}};
  end
`endif

  assign io_resp_0_coh_state = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = T2[5'h15:1'h0];
  MetadataArray_tag_arr tag_arr (
    .CLK(clk),
    .W0A(T17),
    .W0E(T16),
    .W0I(wdata),
    .W0M(T4),
    .R1A(io_read_bits_idx),
    .R1E(io_read_valid),
    .R1O(T2)
  );
  assign T4 = T5;
  assign T5 = 22'h0 - T6;
  assign T6 = {21'h0, T7};
  assign T7 = wmask;
  assign wmask = T8 ? 1'h1 : io_write_bits_way_en;
  assign T8 = rst_cnt < 7'h40;
  assign T9 = reset ? 7'h0 : T10;
  assign T10 = T8 ? T11 : rst_cnt;
  assign T11 = rst_cnt + 7'h1;
  assign wdata = T12;
  assign T12 = {T15, T13};
  assign T13 = T8 ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign rstVal_coh_state = T14;
  assign T14 = 2'h0;
  assign T15 = T8 ? rstVal_tag : io_write_bits_data_tag;
  assign rstVal_tag = 20'h0;
  assign T16 = T8 | io_write_valid;
  assign T17 = waddr[3'h5:1'h0];
  assign waddr = T8 ? rst_cnt : T18;
  assign T18 = {1'h0, io_write_bits_idx};
  assign T20 = io_read_valid ? io_read_bits_idx : R19;
  assign io_resp_0_tag = T21;
  assign T21 = T1[5'h15:2'h2];
  assign io_write_ready = T22;
  assign T22 = T8 ^ 1'h1;
  assign io_read_ready = T23;
  assign T23 = T25 & T24;
  assign T24 = io_write_valid ^ 1'h1;
  assign T25 = T8 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else if(T8) begin
      rst_cnt <= T11;
    end
    if(io_read_valid) begin
      R19 <= io_read_bits_idx;
    end
  end
endmodule

module Arbiter_7(
    output io_in_4_ready,
    input  io_in_4_valid,
    input [5:0] io_in_4_bits_idx,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [5:0] io_in_3_bits_idx,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [5:0] io_in_2_bits_idx,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [5:0] io_in_1_bits_idx,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [5:0] io_in_0_bits_idx,
    input  io_out_ready,
    output io_out_valid,
    output[5:0] io_out_bits_idx,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[5:0] T5;
  wire[5:0] T6;
  wire[5:0] T7;
  wire T8;
  wire[2:0] T9;
  wire[5:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : 3'h4;
  assign io_out_bits_idx = T5;
  assign T5 = T13 ? io_in_4_bits_idx : T6;
  assign T6 = T12 ? T10 : T7;
  assign T7 = T8 ? io_in_1_bits_idx : io_in_0_bits_idx;
  assign T8 = T9[1'h0:1'h0];
  assign T9 = T0;
  assign T10 = T11 ? io_in_3_bits_idx : io_in_2_bits_idx;
  assign T11 = T9[1'h0:1'h0];
  assign T12 = T9[1'h1:1'h1];
  assign T13 = T9[2'h2:2'h2];
  assign io_out_valid = T14;
  assign T14 = T21 ? io_in_4_valid : T15;
  assign T15 = T20 ? T18 : T16;
  assign T16 = T17 ? io_in_1_valid : io_in_0_valid;
  assign T17 = T9[1'h0:1'h0];
  assign T18 = T19 ? io_in_3_valid : io_in_2_valid;
  assign T19 = T9[1'h0:1'h0];
  assign T20 = T9[1'h1:1'h1];
  assign T21 = T9[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T22;
  assign T22 = T23 & io_out_ready;
  assign T23 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T24;
  assign T24 = T25 & io_out_ready;
  assign T25 = T26 ^ 1'h1;
  assign T26 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T27;
  assign T27 = T28 & io_out_ready;
  assign T28 = T29 ^ 1'h1;
  assign T29 = T30 | io_in_2_valid;
  assign T30 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T31;
  assign T31 = T32 & io_out_ready;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T34 | io_in_3_valid;
  assign T34 = T35 | io_in_2_valid;
  assign T35 = io_in_0_valid | io_in_1_valid;
endmodule

module DataArray(input clk,
    output io_read_ready,
    input  io_read_valid,
    input  io_read_bits_way_en,
    input [11:0] io_read_bits_addr,
    output io_write_ready,
    input  io_write_valid,
    input  io_write_bits_way_en,
    input [11:0] io_write_bits_addr,
    input [1:0] io_write_bits_wmask,
    input [127:0] io_write_bits_data,
    output[127:0] io_resp_0
);

  wire[127:0] T0;
  wire T1;
  wire[7:0] raddr;
  wire[127:0] T3;
  wire[127:0] T4;
  wire[127:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire T11;
  wire T12;
  wire[7:0] waddr;
  reg [7:0] R13;
  wire[7:0] T14;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R13 = {1{$random}};
  end
`endif

  assign io_resp_0 = T0;
  assign T1 = io_read_bits_way_en & io_read_valid;
  assign raddr = io_read_bits_addr >> 3'h4;
  DataArray_T2 T2 (
    .CLK(clk),
    .W0A(waddr),
    .W0E(T12),
    .W0I(io_write_bits_data),
    .W0M(T4),
    .R1A(raddr),
    .R1E(T1),
    .R1O(T0)
  );
  assign T4 = T5;
  assign T5 = {T9, T6};
  assign T6 = 64'h0 - T7;
  assign T7 = {63'h0, T8};
  assign T8 = io_write_bits_wmask[1'h0:1'h0];
  assign T9 = 64'h0 - T10;
  assign T10 = {63'h0, T11};
  assign T11 = io_write_bits_wmask[1'h1:1'h1];
  assign T12 = io_write_bits_way_en & io_write_valid;
  assign waddr = io_write_bits_addr >> 3'h4;
  assign T14 = T1 ? raddr : R13;
  assign io_write_ready = 1'h1;
  assign io_read_ready = 1'h1;

  always @(posedge clk) begin
    if(T1) begin
      R13 <= raddr;
    end
  end
endmodule

module Arbiter_8(
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits_way_en,
    input [11:0] io_in_3_bits_addr,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits_way_en,
    input [11:0] io_in_2_bits_addr,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[11:0] T4;
  wire[11:0] T5;
  wire T6;
  wire[1:0] T7;
  wire[11:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 2'h0 : T2;
  assign T2 = io_in_1_valid ? 2'h1 : T3;
  assign T3 = io_in_2_valid ? 2'h2 : 2'h3;
  assign io_out_bits_addr = T4;
  assign T4 = T10 ? T8 : T5;
  assign T5 = T6 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = T0;
  assign T8 = T9 ? io_in_3_bits_addr : io_in_2_bits_addr;
  assign T9 = T7[1'h0:1'h0];
  assign T10 = T7[1'h1:1'h1];
  assign io_out_bits_way_en = T11;
  assign T11 = T16 ? T14 : T12;
  assign T12 = T13 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign T13 = T7[1'h0:1'h0];
  assign T14 = T15 ? io_in_3_bits_way_en : io_in_2_bits_way_en;
  assign T15 = T7[1'h0:1'h0];
  assign T16 = T7[1'h1:1'h1];
  assign io_out_valid = T17;
  assign T17 = T22 ? T20 : T18;
  assign T18 = T19 ? io_in_1_valid : io_in_0_valid;
  assign T19 = T7[1'h0:1'h0];
  assign T20 = T21 ? io_in_3_valid : io_in_2_valid;
  assign T21 = T7[1'h0:1'h0];
  assign T22 = T7[1'h1:1'h1];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T25;
  assign T25 = T26 & io_out_ready;
  assign T26 = T27 ^ 1'h1;
  assign T27 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T30 ^ 1'h1;
  assign T30 = T31 | io_in_2_valid;
  assign T31 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_9(
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits_way_en,
    input [11:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_wmask,
    input [127:0] io_in_1_bits_data,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits_way_en,
    input [11:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_wmask,
    input [127:0] io_in_0_bits_data,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits_way_en,
    output[11:0] io_out_bits_addr,
    output[1:0] io_out_bits_wmask,
    output[127:0] io_out_bits_data,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[127:0] T2;
  wire T3;
  wire[1:0] T4;
  wire[11:0] T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_data = T2;
  assign T2 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign T3 = T0;
  assign io_out_bits_wmask = T4;
  assign T4 = T3 ? io_in_1_bits_wmask : io_in_0_bits_wmask;
  assign io_out_bits_addr = T5;
  assign T5 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_bits_way_en = T6;
  assign T6 = T3 ? io_in_1_bits_way_en : io_in_0_bits_way_en;
  assign io_out_valid = T7;
  assign T7 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T8;
  assign T8 = T9 & io_out_ready;
  assign T9 = io_in_0_valid ^ 1'h1;
endmodule

module AMOALU(
    input [5:0] io_addr,
    input [3:0] io_cmd,
    input [2:0] io_typ,
    input [63:0] io_lhs,
    input [63:0] io_rhs,
    output[63:0] io_out
);

  wire[63:0] T0;
  wire[87:0] T1;
  wire[87:0] T2;
  wire[87:0] T3;
  wire[87:0] T4;
  wire[87:0] wmask;
  wire[87:0] T5;
  wire[47:0] T6;
  wire[23:0] T7;
  wire[15:0] T8;
  wire[7:0] T9;
  wire[7:0] T10;
  wire T11;
  wire[10:0] T12;
  wire[10:0] T13;
  wire[10:0] T14;
  wire[10:0] T15;
  wire[2:0] T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire[10:0] T21;
  wire[8:0] T22;
  wire[2:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire[10:0] T28;
  wire[7:0] T29;
  wire[2:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire T39;
  wire[23:0] T40;
  wire[15:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire T50;
  wire[39:0] T51;
  wire[23:0] T52;
  wire[15:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire T62;
  wire[15:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire T69;
  wire[87:0] T70;
  wire[87:0] T71;
  wire[63:0] out;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] rhs;
  wire[63:0] T78;
  wire[31:0] T79;
  wire[63:0] T80;
  wire[31:0] T81;
  wire[15:0] T82;
  wire[63:0] T83;
  wire[31:0] T84;
  wire[15:0] T85;
  wire[7:0] T86;
  wire T87;
  wire max;
  wire T88;
  wire[4:0] T89;
  wire T90;
  wire[4:0] T91;
  wire min;
  wire T92;
  wire[4:0] T93;
  wire T94;
  wire[4:0] T95;
  wire less;
  wire T96;
  wire cmp_rhs;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire word;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire cmp_lhs;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire sgned;
  wire T113;
  wire[4:0] T114;
  wire T115;
  wire[4:0] T116;
  wire lt;
  wire T117;
  wire T118;
  wire T119;
  wire[31:0] T120;
  wire[31:0] T121;
  wire eq_hi;
  wire[31:0] T122;
  wire[31:0] T123;
  wire T124;
  wire[31:0] T125;
  wire[31:0] T126;
  wire T127;
  wire T128;
  wire T129;
  wire[63:0] T130;
  wire T131;
  wire[4:0] T132;
  wire[63:0] T133;
  wire T134;
  wire[4:0] T135;
  wire[63:0] T136;
  wire T137;
  wire[4:0] T138;
  wire[63:0] adder_out;
  wire[63:0] T139;
  wire[63:0] mask;
  wire[63:0] T140;
  wire[31:0] T141;
  wire T142;
  wire[63:0] T143;
  wire[63:0] T144;
  wire T145;
  wire[4:0] T146;


  assign io_out = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = T70 | T2;
  assign T2 = T4 & T3;
  assign T3 = {24'h0, io_lhs};
  assign T4 = ~ wmask;
  assign wmask = T5;
  assign T5 = {T51, T6};
  assign T6 = {T40, T7};
  assign T7 = {T37, T8};
  assign T8 = {T34, T9};
  assign T9 = 8'h0 - T10;
  assign T10 = {7'h0, T11};
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T31 ? T28 : T13;
  assign T13 = T25 ? T21 : T14;
  assign T14 = T18 ? T15 : 11'hff;
  assign T15 = 4'hf << T16;
  assign T16 = {T17, 2'h0};
  assign T17 = io_addr[2'h2:2'h2];
  assign T18 = T20 | T19;
  assign T19 = io_typ == 3'h6;
  assign T20 = io_typ == 3'h2;
  assign T21 = {2'h0, T22};
  assign T22 = 2'h3 << T23;
  assign T23 = {T24, 1'h0};
  assign T24 = io_addr[2'h2:1'h1];
  assign T25 = T27 | T26;
  assign T26 = io_typ == 3'h5;
  assign T27 = io_typ == 3'h1;
  assign T28 = {3'h0, T29};
  assign T29 = 1'h1 << T30;
  assign T30 = io_addr[2'h2:1'h0];
  assign T31 = T33 | T32;
  assign T32 = io_typ == 3'h4;
  assign T33 = io_typ == 3'h0;
  assign T34 = 8'h0 - T35;
  assign T35 = {7'h0, T36};
  assign T36 = T12[1'h1:1'h1];
  assign T37 = 8'h0 - T38;
  assign T38 = {7'h0, T39};
  assign T39 = T12[2'h2:2'h2];
  assign T40 = {T48, T41};
  assign T41 = {T45, T42};
  assign T42 = 8'h0 - T43;
  assign T43 = {7'h0, T44};
  assign T44 = T12[2'h3:2'h3];
  assign T45 = 8'h0 - T46;
  assign T46 = {7'h0, T47};
  assign T47 = T12[3'h4:3'h4];
  assign T48 = 8'h0 - T49;
  assign T49 = {7'h0, T50};
  assign T50 = T12[3'h5:3'h5];
  assign T51 = {T63, T52};
  assign T52 = {T60, T53};
  assign T53 = {T57, T54};
  assign T54 = 8'h0 - T55;
  assign T55 = {7'h0, T56};
  assign T56 = T12[3'h6:3'h6];
  assign T57 = 8'h0 - T58;
  assign T58 = {7'h0, T59};
  assign T59 = T12[3'h7:3'h7];
  assign T60 = 8'h0 - T61;
  assign T61 = {7'h0, T62};
  assign T62 = T12[4'h8:4'h8];
  assign T63 = {T67, T64};
  assign T64 = 8'h0 - T65;
  assign T65 = {7'h0, T66};
  assign T66 = T12[4'h9:4'h9];
  assign T67 = 8'h0 - T68;
  assign T68 = {7'h0, T69};
  assign T69 = T12[4'ha:4'ha];
  assign T70 = wmask & T71;
  assign T71 = {24'h0, out};
  assign out = T145 ? adder_out : T72;
  assign T72 = T137 ? T136 : T73;
  assign T73 = T134 ? T133 : T74;
  assign T74 = T131 ? T130 : T75;
  assign T75 = T87 ? io_lhs : T76;
  assign T76 = T31 ? T83 : T77;
  assign T77 = T25 ? T80 : rhs;
  assign rhs = T18 ? T78 : io_rhs;
  assign T78 = {T79, T79};
  assign T79 = io_rhs[5'h1f:1'h0];
  assign T80 = {T81, T81};
  assign T81 = {T82, T82};
  assign T82 = io_rhs[4'hf:1'h0];
  assign T83 = {T84, T84};
  assign T84 = {T85, T85};
  assign T85 = {T86, T86};
  assign T86 = io_rhs[3'h7:1'h0];
  assign T87 = less ? min : max;
  assign max = T90 | T88;
  assign T88 = T89 == 5'hf;
  assign T89 = {1'h0, io_cmd};
  assign T90 = T91 == 5'hd;
  assign T91 = {1'h0, io_cmd};
  assign min = T94 | T92;
  assign T92 = T93 == 5'he;
  assign T93 = {1'h0, io_cmd};
  assign T94 = T95 == 5'hc;
  assign T95 = {1'h0, io_cmd};
  assign less = T129 ? lt : T96;
  assign T96 = sgned ? cmp_lhs : cmp_rhs;
  assign cmp_rhs = T99 ? T98 : T97;
  assign T97 = rhs[6'h3f:6'h3f];
  assign T98 = rhs[5'h1f:5'h1f];
  assign T99 = word & T100;
  assign T100 = T101 ^ 1'h1;
  assign T101 = io_addr[2'h2:2'h2];
  assign word = T103 | T102;
  assign T102 = io_typ == 3'h4;
  assign T103 = T105 | T104;
  assign T104 = io_typ == 3'h0;
  assign T105 = T107 | T106;
  assign T106 = io_typ == 3'h6;
  assign T107 = io_typ == 3'h2;
  assign cmp_lhs = T110 ? T109 : T108;
  assign T108 = io_lhs[6'h3f:6'h3f];
  assign T109 = io_lhs[5'h1f:5'h1f];
  assign T110 = word & T111;
  assign T111 = T112 ^ 1'h1;
  assign T112 = io_addr[2'h2:2'h2];
  assign sgned = T115 | T113;
  assign T113 = T114 == 5'hd;
  assign T114 = {1'h0, io_cmd};
  assign T115 = T116 == 5'hc;
  assign T116 = {1'h0, io_cmd};
  assign lt = word ? T127 : T117;
  assign T117 = T124 | T118;
  assign T118 = eq_hi & T119;
  assign T119 = T121 < T120;
  assign T120 = rhs[5'h1f:1'h0];
  assign T121 = io_lhs[5'h1f:1'h0];
  assign eq_hi = T123 == T122;
  assign T122 = rhs[6'h3f:6'h20];
  assign T123 = io_lhs[6'h3f:6'h20];
  assign T124 = T126 < T125;
  assign T125 = rhs[6'h3f:6'h20];
  assign T126 = io_lhs[6'h3f:6'h20];
  assign T127 = T128 ? T124 : T119;
  assign T128 = io_addr[2'h2:2'h2];
  assign T129 = cmp_lhs == cmp_rhs;
  assign T130 = io_lhs ^ rhs;
  assign T131 = T132 == 5'h9;
  assign T132 = {1'h0, io_cmd};
  assign T133 = io_lhs | rhs;
  assign T134 = T135 == 5'ha;
  assign T135 = {1'h0, io_cmd};
  assign T136 = io_lhs & rhs;
  assign T137 = T138 == 5'hb;
  assign T138 = {1'h0, io_cmd};
  assign adder_out = T143 + T139;
  assign T139 = rhs & mask;
  assign mask = 64'hffffffffffffffff ^ T140;
  assign T140 = {32'h0, T141};
  assign T141 = T142 << 5'h1f;
  assign T142 = io_addr[2'h2:2'h2];
  assign T143 = T144;
  assign T144 = io_lhs & mask;
  assign T145 = T146 == 5'h8;
  assign T146 = {1'h0, io_cmd};
endmodule

module Arbiter_10(
    output io_in_1_ready,
    input  io_in_1_valid,
    input [25:0] io_in_1_bits_addr,
    input [1:0] io_in_1_bits_client_xact_id,
    input [2:0] io_in_1_bits_master_xact_id,
    input [511:0] io_in_1_bits_data,
    input [2:0] io_in_1_bits_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [25:0] io_in_0_bits_addr,
    input [1:0] io_in_0_bits_client_xact_id,
    input [2:0] io_in_0_bits_master_xact_id,
    input [511:0] io_in_0_bits_data,
    input [2:0] io_in_0_bits_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[25:0] io_out_bits_addr,
    output[1:0] io_out_bits_client_xact_id,
    output[2:0] io_out_bits_master_xact_id,
    output[511:0] io_out_bits_data,
    output[2:0] io_out_bits_r_type,
    output io_chosen
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire T3;
  wire[511:0] T4;
  wire[2:0] T5;
  wire[1:0] T6;
  wire[25:0] T7;
  wire T8;
  wire T9;
  wire T10;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid == 1'h0;
  assign io_out_bits_r_type = T2;
  assign T2 = T3 ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign T3 = T0;
  assign io_out_bits_data = T4;
  assign T4 = T3 ? io_in_1_bits_data : io_in_0_bits_data;
  assign io_out_bits_master_xact_id = T5;
  assign T5 = T3 ? io_in_1_bits_master_xact_id : io_in_0_bits_master_xact_id;
  assign io_out_bits_client_xact_id = T6;
  assign T6 = T3 ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign io_out_bits_addr = T7;
  assign T7 = T3 ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign io_out_valid = T8;
  assign T8 = T3 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T9;
  assign T9 = T10 & io_out_ready;
  assign T10 = io_in_0_valid ^ 1'h1;
endmodule

module FlowThroughSerializer_1(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [1:0] io_in_bits_header_src,
    input [1:0] io_in_bits_header_dst,
    input [511:0] io_in_bits_payload_data,
    input [1:0] io_in_bits_payload_client_xact_id,
    input [2:0] io_in_bits_payload_master_xact_id,
    input [3:0] io_in_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_cnt,
    output io_done
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  reg  active;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire wrap;
  reg [1:0] cnt;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire[3:0] T23;
  reg [3:0] rbits_payload_g_type;
  wire[3:0] T24;
  wire[3:0] T25;
  wire[2:0] T26;
  reg [2:0] rbits_payload_master_xact_id;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[1:0] T29;
  reg [1:0] rbits_payload_client_xact_id;
  wire[1:0] T30;
  wire[1:0] T31;
  wire[511:0] T32;
  wire[511:0] T33;
  reg [511:0] rbits_payload_data;
  wire[511:0] T34;
  wire[511:0] T35;
  wire[511:0] T36;
  wire[127:0] T37;
  wire[127:0] T38;
  wire[127:0] shifter_0;
  wire[127:0] T39;
  wire[127:0] shifter_1;
  wire[127:0] T40;
  wire T41;
  wire[1:0] T42;
  wire[127:0] T43;
  wire[127:0] shifter_2;
  wire[127:0] T44;
  wire[127:0] shifter_3;
  wire[127:0] T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  reg [1:0] rbits_header_dst;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  reg [1:0] rbits_header_src;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire T55;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    active = {1{$random}};
    cnt = {1{$random}};
    rbits_payload_g_type = {1{$random}};
    rbits_payload_master_xact_id = {1{$random}};
    rbits_payload_client_xact_id = {1{$random}};
    rbits_payload_data = {16{$random}};
    rbits_header_dst = {1{$random}};
    rbits_header_src = {1{$random}};
  end
`endif

  assign io_done = T0;
  assign T0 = T15 ? 1'h1 : T1;
  assign T1 = T6 ? T2 : 1'h0;
  assign T2 = T3 ^ 1'h1;
  assign T3 = T5 | T4;
  assign T4 = io_in_bits_payload_g_type == 4'h2;
  assign T5 = io_in_bits_payload_g_type == 4'h1;
  assign T6 = T7 & io_in_valid;
  assign T7 = active ^ 1'h1;
  assign T8 = reset ? 1'h0 : T9;
  assign T9 = T15 ? 1'h0 : T10;
  assign T10 = T11 ? 1'h1 : active;
  assign T11 = T6 & T12;
  assign T12 = T14 | T13;
  assign T13 = io_in_bits_payload_g_type == 4'h2;
  assign T14 = io_in_bits_payload_g_type == 4'h1;
  assign T15 = T22 & wrap;
  assign wrap = cnt == 2'h3;
  assign T16 = reset ? 2'h0 : T17;
  assign T17 = T15 ? 2'h0 : T18;
  assign T18 = T22 ? T21 : T19;
  assign T19 = T11 ? T20 : cnt;
  assign T20 = {1'h0, io_out_ready};
  assign T21 = cnt + 2'h1;
  assign T22 = active & io_out_ready;
  assign io_cnt = cnt;
  assign io_out_bits_payload_g_type = T23;
  assign T23 = active ? rbits_payload_g_type : io_in_bits_payload_g_type;
  assign T24 = reset ? io_in_bits_payload_g_type : T25;
  assign T25 = T11 ? io_in_bits_payload_g_type : rbits_payload_g_type;
  assign io_out_bits_payload_master_xact_id = T26;
  assign T26 = active ? rbits_payload_master_xact_id : io_in_bits_payload_master_xact_id;
  assign T27 = reset ? io_in_bits_payload_master_xact_id : T28;
  assign T28 = T11 ? io_in_bits_payload_master_xact_id : rbits_payload_master_xact_id;
  assign io_out_bits_payload_client_xact_id = T29;
  assign T29 = active ? rbits_payload_client_xact_id : io_in_bits_payload_client_xact_id;
  assign T30 = reset ? io_in_bits_payload_client_xact_id : T31;
  assign T31 = T11 ? io_in_bits_payload_client_xact_id : rbits_payload_client_xact_id;
  assign io_out_bits_payload_data = T32;
  assign T32 = active ? T36 : T33;
  assign T33 = active ? rbits_payload_data : io_in_bits_payload_data;
  assign T34 = reset ? io_in_bits_payload_data : T35;
  assign T35 = T11 ? io_in_bits_payload_data : rbits_payload_data;
  assign T36 = {384'h0, T37};
  assign T37 = T47 ? T43 : T38;
  assign T38 = T41 ? shifter_1 : shifter_0;
  assign shifter_0 = T39;
  assign T39 = rbits_payload_data[7'h7f:1'h0];
  assign shifter_1 = T40;
  assign T40 = rbits_payload_data[8'hff:8'h80];
  assign T41 = T42[1'h0:1'h0];
  assign T42 = cnt;
  assign T43 = T46 ? shifter_3 : shifter_2;
  assign shifter_2 = T44;
  assign T44 = rbits_payload_data[9'h17f:9'h100];
  assign shifter_3 = T45;
  assign T45 = rbits_payload_data[9'h1ff:9'h180];
  assign T46 = T42[1'h0:1'h0];
  assign T47 = T42[1'h1:1'h1];
  assign io_out_bits_header_dst = T48;
  assign T48 = active ? rbits_header_dst : io_in_bits_header_dst;
  assign T49 = reset ? io_in_bits_header_dst : T50;
  assign T50 = T11 ? io_in_bits_header_dst : rbits_header_dst;
  assign io_out_bits_header_src = T51;
  assign T51 = active ? rbits_header_src : io_in_bits_header_src;
  assign T52 = reset ? io_in_bits_header_src : T53;
  assign T53 = T11 ? io_in_bits_header_src : rbits_header_src;
  assign io_out_valid = T54;
  assign T54 = active | io_in_valid;
  assign io_in_ready = T55;
  assign T55 = active ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else if(T15) begin
      active <= 1'h0;
    end else if(T11) begin
      active <= 1'h1;
    end
    if(reset) begin
      cnt <= 2'h0;
    end else if(T15) begin
      cnt <= 2'h0;
    end else if(T22) begin
      cnt <= T21;
    end else if(T11) begin
      cnt <= T20;
    end
    if(reset) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end else if(T11) begin
      rbits_payload_g_type <= io_in_bits_payload_g_type;
    end
    if(reset) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end else if(T11) begin
      rbits_payload_master_xact_id <= io_in_bits_payload_master_xact_id;
    end
    if(reset) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end else if(T11) begin
      rbits_payload_client_xact_id <= io_in_bits_payload_client_xact_id;
    end
    if(reset) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end else if(T11) begin
      rbits_payload_data <= io_in_bits_payload_data;
    end
    if(reset) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end else if(T11) begin
      rbits_header_dst <= io_in_bits_header_dst;
    end
    if(reset) begin
      rbits_header_src <= io_in_bits_header_src;
    end else if(T11) begin
      rbits_header_src <= io_in_bits_header_src;
    end
  end
endmodule

module HellaCache(input clk, input reset,
    output io_cpu_req_ready,
    input  io_cpu_req_valid,
    input  io_cpu_req_bits_kill,
    input [2:0] io_cpu_req_bits_typ,
    input  io_cpu_req_bits_phys,
    input [43:0] io_cpu_req_bits_addr,
    input [63:0] io_cpu_req_bits_data,
    input [7:0] io_cpu_req_bits_tag,
    input [4:0] io_cpu_req_bits_cmd,
    output io_cpu_resp_valid,
    output io_cpu_resp_bits_nack,
    output io_cpu_resp_bits_replay,
    output[2:0] io_cpu_resp_bits_typ,
    output io_cpu_resp_bits_has_data,
    output[63:0] io_cpu_resp_bits_data,
    output[63:0] io_cpu_resp_bits_data_subword,
    output[7:0] io_cpu_resp_bits_tag,
    output[3:0] io_cpu_resp_bits_cmd,
    output[43:0] io_cpu_resp_bits_addr,
    output[63:0] io_cpu_resp_bits_store_data,
    output io_cpu_replay_next_valid,
    output[7:0] io_cpu_replay_next_bits,
    output io_cpu_xcpt_ma_ld,
    output io_cpu_xcpt_ma_st,
    output io_cpu_xcpt_pf_ld,
    output io_cpu_xcpt_pf_st,
    input  io_cpu_ptw_req_ready,
    output io_cpu_ptw_req_valid,
    output[29:0] io_cpu_ptw_req_bits,
    input  io_cpu_ptw_resp_valid,
    input  io_cpu_ptw_resp_bits_error,
    input [18:0] io_cpu_ptw_resp_bits_ppn,
    input [5:0] io_cpu_ptw_resp_bits_perm,
    input [7:0] io_cpu_ptw_status_ip,
    input [7:0] io_cpu_ptw_status_im,
    input [6:0] io_cpu_ptw_status_zero,
    input  io_cpu_ptw_status_er,
    input  io_cpu_ptw_status_vm,
    input  io_cpu_ptw_status_s64,
    input  io_cpu_ptw_status_u64,
    input  io_cpu_ptw_status_ef,
    input  io_cpu_ptw_status_pei,
    input  io_cpu_ptw_status_ei,
    input  io_cpu_ptw_status_ps,
    input  io_cpu_ptw_status_s,
    input  io_cpu_ptw_invalidate,
    input  io_cpu_ptw_sret,
    output io_cpu_ordered,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    output[1:0] io_mem_finish_bits_header_src,
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    output[1:0] io_mem_release_bits_header_src,
    output[1:0] io_mem_release_bits_header_dst,
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type
);

  wire wb_io_req_ready;
  wire[2:0] prober_io_wb_req_bits_r_type;
  wire[2:0] prober_io_wb_req_bits_master_xact_id;
  wire[1:0] prober_io_wb_req_bits_client_xact_id;
  wire prober_io_wb_req_bits_way_en;
  wire[5:0] prober_io_wb_req_bits_idx;
  wire[19:0] prober_io_wb_req_bits_tag;
  wire prober_io_wb_req_valid;
  wire[2:0] mshrs_io_wb_req_bits_r_type;
  wire[2:0] mshrs_io_wb_req_bits_master_xact_id;
  wire[1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire mshrs_io_wb_req_bits_way_en;
  wire[5:0] mshrs_io_wb_req_bits_idx;
  wire[19:0] mshrs_io_wb_req_bits_tag;
  wire mshrs_io_wb_req_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire[3:0] FlowThroughSerializer_io_out_bits_payload_g_type;
  wire T4;
  wire writeArb_io_in_1_ready;
  wire T5;
  wire[2:0] wb_io_release_bits_r_type;
  wire[511:0] wb_io_release_bits_data;
  wire[2:0] wb_io_release_bits_master_xact_id;
  wire[1:0] wb_io_release_bits_client_xact_id;
  wire[25:0] wb_io_release_bits_addr;
  wire wb_io_release_valid;
  wire[2:0] prober_io_rep_bits_r_type;
  wire[511:0] prober_io_rep_bits_data;
  wire[2:0] prober_io_rep_bits_master_xact_id;
  wire[1:0] prober_io_rep_bits_client_xact_id;
  wire[25:0] prober_io_rep_bits_addr;
  wire prober_io_rep_valid;
  reg [63:0] s2_req_data;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] mshrs_io_replay_bits_data;
  reg  s1_replay;
  wire T9;
  wire T10;
  wire readArb_io_in_1_ready;
  wire mshrs_io_replay_valid;
  wire T11;
  wire s1_write;
  wire T12;
  wire T13;
  reg [4:0] s1_req_cmd;
  wire[4:0] T14;
  wire[4:0] T15;
  wire[4:0] T16;
  wire[4:0] mshrs_io_replay_bits_cmd;
  reg [4:0] s2_req_cmd;
  wire[4:0] T17;
  reg  s1_clk_en;
  wire metaReadArb_io_out_valid;
  wire s2_recycle;
  wire T18;
  reg  s2_recycle_next;
  wire T19;
  wire T20;
  wire T21;
  wire s2_recycle_ecc;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  reg [43:0] s2_req_addr;
  wire[43:0] T28;
  wire[43:0] T29;
  wire[31:0] s1_addr;
  wire[12:0] T30;
  reg [43:0] s1_req_addr;
  wire[43:0] T31;
  wire[43:0] T32;
  wire[43:0] T33;
  wire[43:0] T34;
  wire[43:0] T35;
  wire[43:0] T36;
  wire[31:0] T37;
  wire[25:0] T38;
  wire[5:0] wb_io_meta_read_bits_idx;
  wire[19:0] wb_io_meta_read_bits_tag;
  wire wb_io_meta_read_valid;
  wire[43:0] T39;
  wire[31:0] T40;
  wire[25:0] T41;
  wire[5:0] prober_io_meta_read_bits_idx;
  wire[19:0] prober_io_meta_read_bits_tag;
  wire prober_io_meta_read_valid;
  wire[43:0] mshrs_io_replay_bits_addr;
  wire[18:0] dtlb_io_resp_ppn;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire s2_hit;
  wire T45;
  wire[1:0] T46;
  wire[1:0] T47;
  reg [1:0] s2_hit_state_state;
  wire[1:0] T48;
  wire[1:0] meta_io_resp_0_coh_state;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  reg  s2_tag_match_way;
  wire T78;
  wire s1_tag_match_way;
  wire T79;
  wire T80;
  wire T81;
  wire s1_tag_eq_way;
  wire T82;
  wire[19:0] T83;
  wire[19:0] meta_io_resp_0_tag;
  wire T84;
  wire s2_replay;
  wire T85;
  reg  R86;
  wire T87;
  reg  s2_valid;
  wire T88;
  wire s1_valid_masked;
  wire T89;
  reg  s1_valid;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  reg [63:0] s1_req_data;
  wire[63:0] T98;
  wire[63:0] T99;
  wire[63:0] T100;
  wire T101;
  reg  s1_recycled;
  wire T102;
  wire[63:0] T103;
  wire[127:0] s2_data_word;
  wire[127:0] s2_data_word_prebypass;
  wire[6:0] T104;
  wire[127:0] s2_data_uncorrected;
  wire[127:0] T105;
  wire[63:0] T106;
  wire[127:0] s2_data_muxed;
  wire[127:0] T107;
  wire[127:0] T108;
  reg [63:0] R109;
  wire[63:0] T110;
  wire[127:0] T111;
  wire[127:0] T112;
  wire[127:0] T113;
  wire[127:0] data_io_resp_0;
  wire T114;
  wire T115;
  reg [63:0] R116;
  wire[63:0] T117;
  wire[63:0] T118;
  wire[63:0] T119;
  wire[127:0] T120;
  reg [63:0] s2_store_bypass_data;
  wire[63:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  reg [63:0] s4_req_data;
  wire[63:0] T124;
  reg [63:0] s3_req_data;
  wire[63:0] T125;
  wire[127:0] T126;
  wire[127:0] T127;
  wire[63:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[127:0] T139;
  wire[127:0] T140;
  wire[63:0] amoalu_io_out;
  wire[127:0] s2_data_corrected;
  wire[127:0] T141;
  wire T142;
  reg  s3_valid;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire s2_sc_fail;
  wire T154;
  wire s2_lrsc_addr_match;
  wire T155;
  wire[37:0] T156;
  reg [37:0] lrsc_addr;
  wire[37:0] T157;
  wire[37:0] T158;
  wire T159;
  wire s2_lr;
  wire T160;
  wire T161;
  wire s2_valid_masked;
  wire T162;
  wire T163;
  wire s2_nack;
  wire s2_nack_miss;
  wire T164;
  wire mshrs_io_req_ready;
  wire T165;
  wire T166;
  wire s2_nack_victim;
  wire mshrs_io_secondary_miss;
  reg  s2_nack_hit;
  wire T167;
  wire s1_nack;
  wire T168;
  wire T169;
  wire prober_io_req_ready;
  wire T170;
  wire[5:0] prober_io_meta_write_bits_idx;
  wire[5:0] T171;
  wire T172;
  wire dtlb_io_resp_miss;
  wire T173;
  wire T174;
  reg [4:0] lrsc_count;
  wire[4:0] T175;
  wire[4:0] T176;
  wire[4:0] T177;
  wire[4:0] T178;
  wire[4:0] T179;
  wire[4:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire s2_sc;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  reg [4:0] s3_req_cmd;
  wire[4:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire[40:0] T197;
  reg [43:0] s3_req_addr;
  wire[43:0] T198;
  wire[40:0] T199;
  wire[28:0] T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire[40:0] T211;
  wire[40:0] T212;
  wire[28:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  reg [4:0] s4_req_cmd;
  wire[4:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire[40:0] T230;
  reg [43:0] s4_req_addr;
  wire[43:0] T231;
  wire[40:0] T232;
  wire[28:0] T233;
  reg  s4_valid;
  wire T234;
  wire T235;
  reg  s2_store_bypass;
  wire T236;
  wire T237;
  reg [2:0] s2_req_typ;
  wire[2:0] T238;
  reg [2:0] s1_req_typ;
  wire[2:0] T239;
  wire[2:0] T240;
  wire[2:0] T241;
  wire[2:0] mshrs_io_replay_bits_typ;
  wire[3:0] T242;
  wire[5:0] T243;
  wire data_io_write_ready;
  wire[127:0] T244;
  wire[1:0] T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  reg  s3_way;
  wire T249;
  wire[127:0] T250;
  wire[511:0] FlowThroughSerializer_io_out_bits_payload_data;
  wire[11:0] mshrs_io_mem_resp_addr;
  wire mshrs_io_mem_resp_way_en;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire FlowThroughSerializer_io_out_valid;
  wire T255;
  wire T256;
  wire[11:0] T257;
  wire[11:0] T258;
  wire[11:0] wb_io_data_req_bits_addr;
  wire wb_io_data_req_bits_way_en;
  wire wb_io_data_req_valid;
  wire[11:0] T259;
  wire[127:0] T260;
  wire[127:0] T261;
  wire[63:0] T262;
  wire[127:0] writeArb_io_out_bits_data;
  wire[63:0] T263;
  wire[1:0] writeArb_io_out_bits_wmask;
  wire[11:0] writeArb_io_out_bits_addr;
  wire writeArb_io_out_bits_way_en;
  wire writeArb_io_out_valid;
  wire[11:0] readArb_io_out_bits_addr;
  wire readArb_io_out_bits_way_en;
  wire readArb_io_out_valid;
  wire meta_io_write_ready;
  wire[1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire[19:0] mshrs_io_meta_write_bits_data_tag;
  wire mshrs_io_meta_write_bits_way_en;
  wire[5:0] mshrs_io_meta_write_bits_idx;
  wire mshrs_io_meta_write_valid;
  wire[1:0] prober_io_meta_write_bits_data_coh_state;
  wire[19:0] prober_io_meta_write_bits_data_tag;
  wire prober_io_meta_write_bits_way_en;
  wire prober_io_meta_write_valid;
  wire meta_io_read_ready;
  wire[5:0] T264;
  wire[37:0] T265;
  wire[5:0] mshrs_io_meta_read_bits_idx;
  wire mshrs_io_meta_read_valid;
  wire[5:0] T266;
  wire[37:0] T267;
  wire[1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire[19:0] metaWriteArb_io_out_bits_data_tag;
  wire metaWriteArb_io_out_bits_way_en;
  wire[5:0] metaWriteArb_io_out_bits_idx;
  wire metaWriteArb_io_out_valid;
  wire[5:0] metaReadArb_io_out_bits_idx;
  reg  s1_req_phys;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire mshrs_io_replay_bits_phys;
  reg  s2_req_phys;
  wire T273;
  wire[30:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire s1_readwrite;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire s1_read;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire wbArb_io_in_1_ready;
  wire[2:0] FlowThroughSerializer_io_out_bits_payload_master_xact_id;
  wire[1:0] FlowThroughSerializer_io_out_bits_payload_client_xact_id;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_dst;
  wire[1:0] FlowThroughSerializer_io_out_bits_header_src;
  wire T288;
  wire metaWriteArb_io_in_0_ready;
  wire metaReadArb_io_in_1_ready;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] s2_replaced_way_en;
  reg  R292;
  wire T293;
  wire[1:0] T294;
  wire[1:0] T295;
  reg [1:0] s2_repl_meta_coh_state;
  wire[1:0] T296;
  wire[1:0] T297;
  wire[19:0] T298;
  reg [19:0] s2_repl_meta_tag;
  wire[19:0] T299;
  wire[19:0] T300;
  reg [7:0] s2_req_tag;
  wire[7:0] T301;
  reg [7:0] s1_req_tag;
  wire[7:0] T302;
  wire[7:0] T303;
  wire[7:0] T304;
  wire[7:0] mshrs_io_replay_bits_tag;
  reg  s2_req_kill;
  wire T305;
  reg  s1_req_kill;
  wire T306;
  wire T307;
  wire T308;
  wire mshrs_io_replay_bits_kill;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire mshrs_io_probe_rdy;
  wire wbArb_io_in_0_ready;
  wire metaWriteArb_io_in_1_ready;
  wire metaReadArb_io_in_2_ready;
  wire releaseArb_io_in_1_ready;
  wire[1:0] probe_bits_p_type;
  wire[2:0] probe_bits_master_xact_id;
  wire[25:0] probe_bits_addr;
  wire T332;
  wire T333;
  wire probe_valid;
  wire releaseArb_io_in_0_ready;
  wire readArb_io_in_2_ready;
  wire metaReadArb_io_in_3_ready;
  wire[2:0] wbArb_io_out_bits_r_type;
  wire[2:0] wbArb_io_out_bits_master_xact_id;
  wire[1:0] wbArb_io_out_bits_client_xact_id;
  wire wbArb_io_out_bits_way_en;
  wire[5:0] wbArb_io_out_bits_idx;
  wire[19:0] wbArb_io_out_bits_tag;
  wire wbArb_io_out_valid;
  wire[2:0] T334;
  wire[2:0] releaseArb_io_out_bits_r_type;
  wire[511:0] T335;
  wire[511:0] releaseArb_io_out_bits_data;
  wire[2:0] T336;
  wire[2:0] releaseArb_io_out_bits_master_xact_id;
  wire[1:0] T337;
  wire[1:0] releaseArb_io_out_bits_client_xact_id;
  wire[25:0] T338;
  wire[25:0] releaseArb_io_out_bits_addr;
  wire[1:0] T339;
  wire[1:0] T340;
  wire T341;
  wire releaseArb_io_out_valid;
  wire probe_ready;
  wire T342;
  wire T343;
  wire[2:0] mshrs_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] mshrs_io_mem_finish_bits_header_dst;
  wire[1:0] mshrs_io_mem_finish_bits_header_src;
  wire mshrs_io_mem_finish_valid;
  wire FlowThroughSerializer_io_in_ready;
  wire[3:0] T344;
  wire[3:0] mshrs_io_mem_req_bits_atomic_opcode;
  wire[2:0] T345;
  wire[2:0] mshrs_io_mem_req_bits_subword_addr;
  wire[5:0] T346;
  wire[5:0] mshrs_io_mem_req_bits_write_mask;
  wire[2:0] T347;
  wire[2:0] mshrs_io_mem_req_bits_a_type;
  wire[511:0] T348;
  wire[511:0] mshrs_io_mem_req_bits_data;
  wire[1:0] T349;
  wire[1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire[25:0] T350;
  wire[25:0] mshrs_io_mem_req_bits_addr;
  wire[1:0] T351;
  wire[1:0] T352;
  wire T353;
  wire mshrs_io_mem_req_valid;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire mshrs_io_fence_rdy;
  wire[29:0] dtlb_io_ptw_req_bits;
  wire dtlb_io_ptw_req_valid;
  wire T358;
  wire dtlb_io_resp_xcpt_st;
  wire T359;
  wire dtlb_io_resp_xcpt_ld;
  wire T360;
  wire misaligned;
  wire T361;
  wire T362;
  wire[2:0] T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[1:0] T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire s1_sc;
  wire[3:0] T381;
  wire[63:0] T382;
  wire[63:0] T383;
  wire[63:0] T384;
  wire[7:0] T385;
  wire[7:0] T386;
  wire[7:0] T387;
  wire[63:0] T388;
  wire[15:0] T389;
  wire[15:0] T390;
  wire[63:0] T391;
  wire[31:0] T392;
  wire[31:0] T393;
  wire[31:0] T394;
  wire T395;
  wire[31:0] T396;
  wire[31:0] T397;
  wire[31:0] T398;
  wire[31:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[15:0] T412;
  wire T413;
  wire[47:0] T414;
  wire[47:0] T415;
  wire[47:0] T416;
  wire[47:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire[7:0] T423;
  wire T424;
  wire[55:0] T425;
  wire[55:0] T426;
  wire[55:0] T427;
  wire[55:0] T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire dtlb_io_req_ready;
  wire T455;
  wire metaReadArb_io_in_4_ready;
  wire T456;
  wire readArb_io_in_3_ready;
  reg  block_miss;
  wire T457;
  wire T458;
  wire T459;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    s2_req_data = {2{$random}};
    s1_replay = {1{$random}};
    s1_req_cmd = {1{$random}};
    s2_req_cmd = {1{$random}};
    s1_clk_en = {1{$random}};
    s2_recycle_next = {1{$random}};
    s2_req_addr = {2{$random}};
    s1_req_addr = {2{$random}};
    s2_hit_state_state = {1{$random}};
    s2_tag_match_way = {1{$random}};
    R86 = {1{$random}};
    s2_valid = {1{$random}};
    s1_valid = {1{$random}};
    s1_req_data = {2{$random}};
    s1_recycled = {1{$random}};
    R109 = {2{$random}};
    R116 = {2{$random}};
    s2_store_bypass_data = {2{$random}};
    s4_req_data = {2{$random}};
    s3_req_data = {2{$random}};
    s3_valid = {1{$random}};
    lrsc_addr = {2{$random}};
    s2_nack_hit = {1{$random}};
    lrsc_count = {1{$random}};
    s3_req_cmd = {1{$random}};
    s3_req_addr = {2{$random}};
    s4_req_cmd = {1{$random}};
    s4_req_addr = {2{$random}};
    s4_valid = {1{$random}};
    s2_store_bypass = {1{$random}};
    s2_req_typ = {1{$random}};
    s1_req_typ = {1{$random}};
    s3_way = {1{$random}};
    s1_req_phys = {1{$random}};
    s2_req_phys = {1{$random}};
    R292 = {1{$random}};
    s2_repl_meta_coh_state = {1{$random}};
    s2_repl_meta_tag = {1{$random}};
    s2_req_tag = {1{$random}};
    s1_req_tag = {1{$random}};
    s2_req_kill = {1{$random}};
    s1_req_kill = {1{$random}};
    block_miss = {1{$random}};
  end
`endif

  assign T0 = writeArb_io_in_1_ready | T1;
  assign T1 = T2 ^ 1'h1;
  assign T2 = T4 | T3;
  assign T3 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h2;
  assign T4 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h1;
  assign T5 = io_mem_release_ready;
  assign T6 = T101 ? s1_req_data : T7;
  assign T7 = T11 ? T8 : s2_req_data;
  assign T8 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_req_bits_data;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign T11 = s1_clk_en & s1_write;
  assign s1_write = T95 | T12;
  assign T12 = T94 | T13;
  assign T13 = s1_req_cmd == 5'h4;
  assign T14 = s2_recycle ? s2_req_cmd : T15;
  assign T15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : T16;
  assign T16 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign T17 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign s2_recycle = T18;
  assign T18 = s2_recycle_ecc | s2_recycle_next;
  assign T19 = reset ? 1'h0 : T20;
  assign T20 = T93 ? T21 : s2_recycle_next;
  assign T21 = T92 & s2_recycle_ecc;
  assign s2_recycle_ecc = T44 & T22;
  assign T22 = T42 & T23;
  assign T23 = T24 - 1'h1;
  assign T24 = 1'h1 << T25;
  assign T25 = T26 + 1'h1;
  assign T26 = T27 - T27;
  assign T27 = s2_req_addr[2'h3:2'h3];
  assign T28 = s1_clk_en ? T29 : s2_req_addr;
  assign T29 = {12'h0, s1_addr};
  assign s1_addr = {dtlb_io_resp_ppn, T30};
  assign T30 = s1_req_addr[4'hc:1'h0];
  assign T31 = s2_recycle ? s2_req_addr : T32;
  assign T32 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : T33;
  assign T33 = prober_io_meta_read_valid ? T39 : T34;
  assign T34 = wb_io_meta_read_valid ? T36 : T35;
  assign T35 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign T36 = {12'h0, T37};
  assign T37 = T38 << 3'h6;
  assign T38 = {wb_io_meta_read_bits_tag, wb_io_meta_read_bits_idx};
  assign T39 = {12'h0, T40};
  assign T40 = T41 << 3'h6;
  assign T41 = {prober_io_meta_read_bits_tag, prober_io_meta_read_bits_idx};
  assign T42 = T43 >> T27;
  assign T43 = 2'h0;
  assign T44 = T84 & s2_hit;
  assign s2_hit = T56 & T45;
  assign T45 = s2_hit_state_state == T46;
  assign T46 = T47;
  assign T47 = T49 ? 2'h3 : s2_hit_state_state;
  assign T48 = s1_clk_en ? meta_io_resp_0_coh_state : s2_hit_state_state;
  assign T49 = T53 | T50;
  assign T50 = T52 | T51;
  assign T51 = s2_req_cmd == 5'h4;
  assign T52 = s2_req_cmd[2'h3:2'h3];
  assign T53 = T55 | T54;
  assign T54 = s2_req_cmd == 5'h7;
  assign T55 = s2_req_cmd == 5'h1;
  assign T56 = T77 & T57;
  assign T57 = T66 ? T63 : T58;
  assign T58 = T60 | T59;
  assign T59 = s2_hit_state_state == 2'h3;
  assign T60 = T62 | T61;
  assign T61 = s2_hit_state_state == 2'h2;
  assign T62 = s2_hit_state_state == 2'h1;
  assign T63 = T65 | T64;
  assign T64 = s2_hit_state_state == 2'h3;
  assign T65 = s2_hit_state_state == 2'h2;
  assign T66 = T68 | T67;
  assign T67 = s2_req_cmd == 5'h6;
  assign T68 = T70 | T69;
  assign T69 = s2_req_cmd == 5'h3;
  assign T70 = T74 | T71;
  assign T71 = T73 | T72;
  assign T72 = s2_req_cmd == 5'h4;
  assign T73 = s2_req_cmd[2'h3:2'h3];
  assign T74 = T76 | T75;
  assign T75 = s2_req_cmd == 5'h7;
  assign T76 = s2_req_cmd == 5'h1;
  assign T77 = s2_tag_match_way != 1'h0;
  assign T78 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign s1_tag_match_way = T79;
  assign T79 = T81 & T80;
  assign T80 = meta_io_resp_0_coh_state != 2'h0;
  assign T81 = s1_tag_eq_way;
  assign s1_tag_eq_way = T82;
  assign T82 = meta_io_resp_0_tag == T83;
  assign T83 = s1_addr >> 4'hc;
  assign T84 = s2_valid | s2_replay;
  assign s2_replay = R86 & T85;
  assign T85 = s2_req_cmd != 5'h5;
  assign T87 = reset ? 1'h0 : s1_replay;
  assign T88 = reset ? 1'h0 : s1_valid_masked;
  assign s1_valid_masked = s1_valid & T89;
  assign T89 = io_cpu_req_bits_kill ^ 1'h1;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = io_cpu_req_ready & io_cpu_req_valid;
  assign T92 = s1_valid | s1_replay;
  assign T93 = s1_valid | s1_replay;
  assign T94 = s1_req_cmd[2'h3:2'h3];
  assign T95 = T97 | T96;
  assign T96 = s1_req_cmd == 5'h7;
  assign T97 = s1_req_cmd == 5'h1;
  assign T98 = s2_recycle ? s2_req_data : T99;
  assign T99 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : T100;
  assign T100 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T101 = s1_clk_en & s1_recycled;
  assign T102 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T103 = s2_data_word[6'h3f:1'h0];
  assign s2_data_word = s2_store_bypass ? T120 : s2_data_word_prebypass;
  assign s2_data_word_prebypass = s2_data_uncorrected >> T104;
  assign T104 = {T27, 6'h0};
  assign s2_data_uncorrected = T105;
  assign T105 = {T119, T106};
  assign T106 = s2_data_muxed[6'h3f:1'h0];
  assign s2_data_muxed = T107;
  assign T107 = T108;
  assign T108 = {R116, R109};
  assign T110 = T111[6'h3f:1'h0];
  assign T111 = T114 ? T113 : T112;
  assign T112 = {64'h0, R109};
  assign T113 = data_io_resp_0 >> 1'h0;
  assign T114 = s1_clk_en & T115;
  assign T115 = s1_tag_eq_way;
  assign T117 = T114 ? T118 : R116;
  assign T118 = data_io_resp_0 >> 7'h40;
  assign T119 = s2_data_muxed[7'h7f:7'h40];
  assign T120 = {64'h0, s2_store_bypass_data};
  assign T121 = T217 ? T122 : s2_store_bypass_data;
  assign T122 = T201 ? amoalu_io_out : T123;
  assign T123 = T186 ? s3_req_data : s4_req_data;
  assign T124 = T142 ? s3_req_data : s4_req_data;
  assign T125 = T126[6'h3f:1'h0];
  assign T126 = T129 ? T139 : T127;
  assign T127 = {64'h0, T128};
  assign T128 = T129 ? s2_req_data : s3_req_data;
  assign T129 = T138 & T130;
  assign T130 = T131 | T22;
  assign T131 = T135 | T132;
  assign T132 = T134 | T133;
  assign T133 = s2_req_cmd == 5'h4;
  assign T134 = s2_req_cmd[2'h3:2'h3];
  assign T135 = T137 | T136;
  assign T136 = s2_req_cmd == 5'h7;
  assign T137 = s2_req_cmd == 5'h1;
  assign T138 = s2_valid | s2_replay;
  assign T139 = T22 ? s2_data_corrected : T140;
  assign T140 = {64'h0, amoalu_io_out};
  assign s2_data_corrected = T141;
  assign T141 = {T119, T106};
  assign T142 = s3_valid & metaReadArb_io_out_valid;
  assign T143 = reset ? 1'h0 : T144;
  assign T144 = T152 & T145;
  assign T145 = T149 | T146;
  assign T146 = T148 | T147;
  assign T147 = s2_req_cmd == 5'h4;
  assign T148 = s2_req_cmd[2'h3:2'h3];
  assign T149 = T151 | T150;
  assign T150 = s2_req_cmd == 5'h7;
  assign T151 = s2_req_cmd == 5'h1;
  assign T152 = T184 & T153;
  assign T153 = s2_sc_fail ^ 1'h1;
  assign s2_sc_fail = s2_sc & T154;
  assign T154 = s2_lrsc_addr_match ^ 1'h1;
  assign s2_lrsc_addr_match = T174 & T155;
  assign T155 = lrsc_addr == T156;
  assign T156 = s2_req_addr >> 3'h6;
  assign T157 = T159 ? T158 : lrsc_addr;
  assign T158 = s2_req_addr >> 3'h6;
  assign T159 = T160 & s2_lr;
  assign s2_lr = s2_req_cmd == 5'h6;
  assign T160 = T161 | s2_replay;
  assign T161 = s2_valid_masked & s2_hit;
  assign s2_valid_masked = T162;
  assign T162 = s2_valid & T163;
  assign T163 = s2_nack ^ 1'h1;
  assign s2_nack = T166 | s2_nack_miss;
  assign s2_nack_miss = T165 & T164;
  assign T164 = mshrs_io_req_ready ^ 1'h1;
  assign T165 = s2_hit ^ 1'h1;
  assign T166 = s2_nack_hit | s2_nack_victim;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T167 = T173 ? s1_nack : s2_nack_hit;
  assign s1_nack = T172 | T168;
  assign T168 = T170 & T169;
  assign T169 = prober_io_req_ready ^ 1'h1;
  assign T170 = T171 == prober_io_meta_write_bits_idx;
  assign T171 = s1_req_addr[4'hb:3'h6];
  assign T172 = T275 & dtlb_io_resp_miss;
  assign T173 = s1_valid | s1_replay;
  assign T174 = lrsc_count != 5'h0;
  assign T175 = reset ? 5'h0 : T176;
  assign T176 = io_cpu_ptw_sret ? 5'h0 : T177;
  assign T177 = T183 ? 5'h0 : T178;
  assign T178 = T181 ? 5'h1f : T179;
  assign T179 = T174 ? T180 : lrsc_count;
  assign T180 = lrsc_count - 5'h1;
  assign T181 = T159 & T182;
  assign T182 = T174 ^ 1'h1;
  assign T183 = T160 & s2_sc;
  assign s2_sc = s2_req_cmd == 5'h7;
  assign T184 = T185 | s2_replay;
  assign T185 = s2_valid_masked & s2_hit;
  assign T186 = T195 & T187;
  assign T187 = T192 | T188;
  assign T188 = T191 | T189;
  assign T189 = s3_req_cmd == 5'h4;
  assign T190 = T129 ? s2_req_cmd : s3_req_cmd;
  assign T191 = s3_req_cmd[2'h3:2'h3];
  assign T192 = T194 | T193;
  assign T193 = s3_req_cmd == 5'h7;
  assign T194 = s3_req_cmd == 5'h1;
  assign T195 = s3_valid & T196;
  assign T196 = T199 == T197;
  assign T197 = s3_req_addr >> 2'h3;
  assign T198 = T129 ? s2_req_addr : s3_req_addr;
  assign T199 = {12'h0, T200};
  assign T200 = s1_addr >> 2'h3;
  assign T201 = T209 & T202;
  assign T202 = T206 | T203;
  assign T203 = T205 | T204;
  assign T204 = s2_req_cmd == 5'h4;
  assign T205 = s2_req_cmd[2'h3:2'h3];
  assign T206 = T208 | T207;
  assign T207 = s2_req_cmd == 5'h7;
  assign T208 = s2_req_cmd == 5'h1;
  assign T209 = T214 & T210;
  assign T210 = T212 == T211;
  assign T211 = s2_req_addr >> 2'h3;
  assign T212 = {12'h0, T213};
  assign T213 = s1_addr >> 2'h3;
  assign T214 = T216 & T215;
  assign T215 = s2_sc_fail ^ 1'h1;
  assign T216 = s2_valid_masked | s2_replay;
  assign T217 = s1_clk_en & T218;
  assign T218 = T235 | T219;
  assign T219 = T228 & T220;
  assign T220 = T225 | T221;
  assign T221 = T224 | T222;
  assign T222 = s4_req_cmd == 5'h4;
  assign T223 = T142 ? s3_req_cmd : s4_req_cmd;
  assign T224 = s4_req_cmd[2'h3:2'h3];
  assign T225 = T227 | T226;
  assign T226 = s4_req_cmd == 5'h7;
  assign T227 = s4_req_cmd == 5'h1;
  assign T228 = s4_valid & T229;
  assign T229 = T232 == T230;
  assign T230 = s4_req_addr >> 2'h3;
  assign T231 = T142 ? s3_req_addr : s4_req_addr;
  assign T232 = {12'h0, T233};
  assign T233 = s1_addr >> 2'h3;
  assign T234 = reset ? 1'h0 : s3_valid;
  assign T235 = T201 | T186;
  assign T236 = T217 ? 1'h1 : T237;
  assign T237 = s1_clk_en ? 1'h0 : s2_store_bypass;
  assign T238 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign T239 = s2_recycle ? s2_req_typ : T240;
  assign T240 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : T241;
  assign T241 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign T242 = s2_req_cmd[2'h3:1'h0];
  assign T243 = s2_req_addr[3'h5:1'h0];
  assign T244 = {s3_req_data, s3_req_data};
  assign T245 = 1'h1 << T246;
  assign T246 = T247;
  assign T247 = s3_req_addr[2'h3:2'h3];
  assign T248 = s3_req_addr[4'hb:1'h0];
  assign T249 = T129 ? s2_tag_match_way : s3_way;
  assign T250 = FlowThroughSerializer_io_out_bits_payload_data[7'h7f:1'h0];
  assign T251 = FlowThroughSerializer_io_out_valid & T252;
  assign T252 = T254 | T253;
  assign T253 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h2;
  assign T254 = FlowThroughSerializer_io_out_bits_payload_g_type == 4'h1;
  assign T255 = T256 | T0;
  assign T256 = FlowThroughSerializer_io_out_valid ^ 1'h1;
  assign T257 = s2_req_addr[4'hb:1'h0];
  assign T258 = mshrs_io_replay_bits_addr[4'hb:1'h0];
  assign T259 = io_cpu_req_bits_addr[4'hb:1'h0];
  assign T260 = T261;
  assign T261 = {T263, T262};
  assign T262 = writeArb_io_out_bits_data[6'h3f:1'h0];
  assign T263 = writeArb_io_out_bits_data[7'h7f:7'h40];
  assign T264 = T265[3'h5:1'h0];
  assign T265 = s2_req_addr >> 3'h6;
  assign T266 = T267[3'h5:1'h0];
  assign T267 = io_cpu_req_bits_addr >> 3'h6;
  assign T268 = s2_recycle ? s2_req_phys : T269;
  assign T269 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : T270;
  assign T270 = prober_io_meta_read_valid ? 1'h1 : T271;
  assign T271 = wb_io_meta_read_valid ? 1'h1 : T272;
  assign T272 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign T273 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign T274 = s1_req_addr >> 4'hd;
  assign T275 = T277 & T276;
  assign T276 = s1_req_phys ^ 1'h1;
  assign T277 = s1_valid_masked & s1_readwrite;
  assign s1_readwrite = T281 | T278;
  assign T278 = T280 | T279;
  assign T279 = s1_req_cmd == 5'h3;
  assign T280 = s1_req_cmd == 5'h2;
  assign T281 = s1_read | s1_write;
  assign s1_read = T285 | T282;
  assign T282 = T284 | T283;
  assign T283 = s1_req_cmd == 5'h4;
  assign T284 = s1_req_cmd[2'h3:2'h3];
  assign T285 = T287 | T286;
  assign T286 = s1_req_cmd == 5'h6;
  assign T287 = s1_req_cmd == 5'h0;
  assign T288 = T0 & FlowThroughSerializer_io_out_valid;
  assign T289 = io_mem_acquire_ready;
  assign T290 = T291[1'h0:1'h0];
  assign T291 = T77 ? T294 : s2_replaced_way_en;
  assign s2_replaced_way_en = 1'h1 << R292;
  assign T293 = s1_clk_en ? 1'h0 : R292;
  assign T294 = {1'h0, s2_tag_match_way};
  assign T295 = T77 ? T297 : s2_repl_meta_coh_state;
  assign T296 = s1_clk_en ? meta_io_resp_0_coh_state : s2_repl_meta_coh_state;
  assign T297 = s2_hit_state_state;
  assign T298 = T77 ? T300 : s2_repl_meta_tag;
  assign T299 = s1_clk_en ? meta_io_resp_0_tag : s2_repl_meta_tag;
  assign T300 = s2_repl_meta_tag;
  assign T301 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign T302 = s2_recycle ? s2_req_tag : T303;
  assign T303 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : T304;
  assign T304 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign T305 = s1_clk_en ? s1_req_kill : s2_req_kill;
  assign T306 = s2_recycle ? s2_req_kill : T307;
  assign T307 = mshrs_io_replay_valid ? mshrs_io_replay_bits_kill : T308;
  assign T308 = io_cpu_req_valid ? io_cpu_req_bits_kill : s1_req_kill;
  assign T309 = s2_nack_hit ? 1'h0 : T310;
  assign T310 = T330 & T311;
  assign T311 = T319 | T312;
  assign T312 = T316 | T313;
  assign T313 = T315 | T314;
  assign T314 = s2_req_cmd == 5'h4;
  assign T315 = s2_req_cmd[2'h3:2'h3];
  assign T316 = T318 | T317;
  assign T317 = s2_req_cmd == 5'h7;
  assign T318 = s2_req_cmd == 5'h1;
  assign T319 = T327 | T320;
  assign T320 = T324 | T321;
  assign T321 = T323 | T322;
  assign T322 = s2_req_cmd == 5'h4;
  assign T323 = s2_req_cmd[2'h3:2'h3];
  assign T324 = T326 | T325;
  assign T325 = s2_req_cmd == 5'h6;
  assign T326 = s2_req_cmd == 5'h0;
  assign T327 = T329 | T328;
  assign T328 = s2_req_cmd == 5'h3;
  assign T329 = s2_req_cmd == 5'h2;
  assign T330 = s2_valid_masked & T331;
  assign T331 = s2_hit ^ 1'h1;
  assign probe_bits_p_type = io_mem_probe_bits_payload_p_type;
  assign probe_bits_master_xact_id = io_mem_probe_bits_payload_master_xact_id;
  assign probe_bits_addr = io_mem_probe_bits_payload_addr;
  assign T332 = probe_valid & T333;
  assign T333 = T174 ^ 1'h1;
  assign probe_valid = io_mem_probe_valid;
  assign io_mem_release_bits_payload_r_type = T334;
  assign T334 = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_payload_data = T335;
  assign T335 = releaseArb_io_out_bits_data;
  assign io_mem_release_bits_payload_master_xact_id = T336;
  assign T336 = releaseArb_io_out_bits_master_xact_id;
  assign io_mem_release_bits_payload_client_xact_id = T337;
  assign T337 = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_payload_addr = T338;
  assign T338 = releaseArb_io_out_bits_addr;
  assign io_mem_release_bits_header_dst = T339;
  assign T339 = 2'h0;
  assign io_mem_release_bits_header_src = T340;
  assign T340 = 2'h0;
  assign io_mem_release_valid = T341;
  assign T341 = releaseArb_io_out_valid;
  assign io_mem_probe_ready = probe_ready;
  assign probe_ready = T342;
  assign T342 = prober_io_req_ready & T343;
  assign T343 = T174 ^ 1'h1;
  assign io_mem_finish_bits_payload_master_xact_id = mshrs_io_mem_finish_bits_payload_master_xact_id;
  assign io_mem_finish_bits_header_dst = mshrs_io_mem_finish_bits_header_dst;
  assign io_mem_finish_bits_header_src = mshrs_io_mem_finish_bits_header_src;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_grant_ready = FlowThroughSerializer_io_in_ready;
  assign io_mem_acquire_bits_payload_atomic_opcode = T344;
  assign T344 = mshrs_io_mem_req_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = T345;
  assign T345 = mshrs_io_mem_req_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = T346;
  assign T346 = mshrs_io_mem_req_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = T347;
  assign T347 = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_payload_data = T348;
  assign T348 = mshrs_io_mem_req_bits_data;
  assign io_mem_acquire_bits_payload_client_xact_id = T349;
  assign T349 = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = T350;
  assign T350 = mshrs_io_mem_req_bits_addr;
  assign io_mem_acquire_bits_header_dst = T351;
  assign T351 = 2'h0;
  assign io_mem_acquire_bits_header_src = T352;
  assign T352 = 2'h0;
  assign io_mem_acquire_valid = T353;
  assign T353 = mshrs_io_mem_req_valid;
  assign io_cpu_ordered = T354;
  assign T354 = T356 & T355;
  assign T355 = s2_valid ^ 1'h1;
  assign T356 = mshrs_io_fence_rdy & T357;
  assign T357 = s1_valid ^ 1'h1;
  assign io_cpu_ptw_req_bits = dtlb_io_ptw_req_bits;
  assign io_cpu_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_cpu_xcpt_pf_st = T358;
  assign T358 = s1_write & dtlb_io_resp_xcpt_st;
  assign io_cpu_xcpt_pf_ld = T359;
  assign T359 = s1_read & dtlb_io_resp_xcpt_ld;
  assign io_cpu_xcpt_ma_st = T360;
  assign T360 = s1_write & misaligned;
  assign misaligned = T365 | T361;
  assign T361 = T364 & T362;
  assign T362 = T363 != 3'h0;
  assign T363 = s1_req_addr[2'h2:1'h0];
  assign T364 = s1_req_typ == 3'h3;
  assign T365 = T372 | T366;
  assign T366 = T369 & T367;
  assign T367 = T368 != 2'h0;
  assign T368 = s1_req_addr[1'h1:1'h0];
  assign T369 = T371 | T370;
  assign T370 = s1_req_typ == 3'h6;
  assign T371 = s1_req_typ == 3'h2;
  assign T372 = T375 & T373;
  assign T373 = T374 != 1'h0;
  assign T374 = s1_req_addr[1'h0:1'h0];
  assign T375 = T377 | T376;
  assign T376 = s1_req_typ == 3'h5;
  assign T377 = s1_req_typ == 3'h1;
  assign io_cpu_xcpt_ma_ld = T378;
  assign T378 = s1_read & misaligned;
  assign io_cpu_replay_next_bits = s1_req_tag;
  assign io_cpu_replay_next_valid = T379;
  assign T379 = s1_replay & T380;
  assign T380 = s1_read | s1_sc;
  assign s1_sc = s1_req_cmd == 5'h7;
  assign io_cpu_resp_bits_store_data = s2_req_data;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_cmd = T381;
  assign T381 = s2_req_cmd[2'h3:1'h0];
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data_subword = T382;
  assign T382 = T384 | T383;
  assign T383 = {63'h0, s2_sc_fail};
  assign T384 = {T425, T385};
  assign T385 = s2_sc ? 8'h0 : T386;
  assign T386 = T424 ? T423 : T387;
  assign T387 = T388[3'h7:1'h0];
  assign T388 = {T414, T389};
  assign T389 = T413 ? T412 : T390;
  assign T390 = T391[4'hf:1'h0];
  assign T391 = {T396, T392};
  assign T392 = T395 ? T394 : T393;
  assign T393 = s2_data_word[5'h1f:1'h0];
  assign T394 = s2_data_word[6'h3f:6'h20];
  assign T395 = s2_req_addr[2'h2:2'h2];
  assign T396 = T409 ? T398 : T397;
  assign T397 = s2_data_word[6'h3f:6'h20];
  assign T398 = 32'h0 - T399;
  assign T399 = {31'h0, T400};
  assign T400 = T402 & T401;
  assign T401 = T392[5'h1f:5'h1f];
  assign T402 = T404 | T403;
  assign T403 = s2_req_typ == 3'h3;
  assign T404 = T406 | T405;
  assign T405 = s2_req_typ == 3'h2;
  assign T406 = T408 | T407;
  assign T407 = s2_req_typ == 3'h1;
  assign T408 = s2_req_typ == 3'h0;
  assign T409 = T411 | T410;
  assign T410 = s2_req_typ == 3'h6;
  assign T411 = s2_req_typ == 3'h2;
  assign T412 = T391[5'h1f:5'h10];
  assign T413 = s2_req_addr[1'h1:1'h1];
  assign T414 = T420 ? T416 : T415;
  assign T415 = T391[6'h3f:5'h10];
  assign T416 = 48'h0 - T417;
  assign T417 = {47'h0, T418};
  assign T418 = T402 & T419;
  assign T419 = T389[4'hf:4'hf];
  assign T420 = T422 | T421;
  assign T421 = s2_req_typ == 3'h5;
  assign T422 = s2_req_typ == 3'h1;
  assign T423 = T388[4'hf:4'h8];
  assign T424 = s2_req_addr[1'h0:1'h0];
  assign T425 = T431 ? T427 : T426;
  assign T426 = T388[6'h3f:4'h8];
  assign T427 = 56'h0 - T428;
  assign T428 = {55'h0, T429};
  assign T429 = T402 & T430;
  assign T430 = T385[3'h7:3'h7];
  assign T431 = s2_sc | T432;
  assign T432 = T434 | T433;
  assign T433 = s2_req_typ == 3'h4;
  assign T434 = s2_req_typ == 3'h0;
  assign io_cpu_resp_bits_data = T391;
  assign io_cpu_resp_bits_has_data = T435;
  assign T435 = T436 | s2_sc;
  assign T436 = T440 | T437;
  assign T437 = T439 | T438;
  assign T438 = s2_req_cmd == 5'h4;
  assign T439 = s2_req_cmd[2'h3:2'h3];
  assign T440 = T442 | T441;
  assign T441 = s2_req_cmd == 5'h6;
  assign T442 = s2_req_cmd == 5'h0;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_replay = s2_replay;
  assign io_cpu_resp_bits_nack = T443;
  assign T443 = s2_valid & s2_nack;
  assign io_cpu_resp_valid = T444;
  assign T444 = T446 & T445;
  assign T445 = T22 ^ 1'h1;
  assign T446 = s2_replay | T447;
  assign T447 = s2_valid_masked & s2_hit;
  assign io_cpu_req_ready = T448;
  assign T448 = block_miss ? 1'h0 : T449;
  assign T449 = T456 ? 1'h0 : T450;
  assign T450 = T455 ? 1'h0 : T451;
  assign T451 = T452 == 1'h0;
  assign T452 = T454 & T453;
  assign T453 = io_cpu_req_bits_phys ^ 1'h1;
  assign T454 = dtlb_io_req_ready ^ 1'h1;
  assign T455 = metaReadArb_io_in_4_ready ^ 1'h1;
  assign T456 = readArb_io_in_3_ready ^ 1'h1;
  assign T457 = reset ? 1'h0 : T458;
  assign T458 = T459 & s2_nack_miss;
  assign T459 = s2_valid | block_miss;
  WritebackUnit wb(.clk(clk), .reset(reset),
       .io_req_ready( wb_io_req_ready ),
       .io_req_valid( wbArb_io_out_valid ),
       .io_req_bits_tag( wbArb_io_out_bits_tag ),
       .io_req_bits_idx( wbArb_io_out_bits_idx ),
       .io_req_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_req_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_req_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_req_bits_r_type( wbArb_io_out_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_3_ready ),
       .io_meta_read_valid( wb_io_meta_read_valid ),
       .io_meta_read_bits_idx( wb_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( wb_io_meta_read_bits_tag ),
       .io_data_req_ready( readArb_io_in_2_ready ),
       .io_data_req_valid( wb_io_data_req_valid ),
       .io_data_req_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_data_req_bits_addr( wb_io_data_req_bits_addr ),
       .io_data_resp( s2_data_corrected ),
       .io_release_ready( releaseArb_io_in_0_ready ),
       .io_release_valid( wb_io_release_valid ),
       .io_release_bits_addr( wb_io_release_bits_addr ),
       .io_release_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_release_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_release_bits_data( wb_io_release_bits_data ),
       .io_release_bits_r_type( wb_io_release_bits_r_type )
  );
  ProbeUnit prober(.clk(clk), .reset(reset),
       .io_req_ready( prober_io_req_ready ),
       .io_req_valid( T332 ),
       .io_req_bits_addr( probe_bits_addr ),
       .io_req_bits_master_xact_id( probe_bits_master_xact_id ),
       .io_req_bits_p_type( probe_bits_p_type ),
       //.io_req_bits_client_xact_id(  )
       .io_rep_ready( releaseArb_io_in_1_ready ),
       .io_rep_valid( prober_io_rep_valid ),
       .io_rep_bits_addr( prober_io_rep_bits_addr ),
       .io_rep_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_rep_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_rep_bits_data( prober_io_rep_bits_data ),
       .io_rep_bits_r_type( prober_io_rep_bits_r_type ),
       .io_meta_read_ready( metaReadArb_io_in_2_ready ),
       .io_meta_read_valid( prober_io_meta_read_valid ),
       .io_meta_read_bits_idx( prober_io_meta_read_bits_idx ),
       .io_meta_read_bits_tag( prober_io_meta_read_bits_tag ),
       .io_meta_write_ready( metaWriteArb_io_in_1_ready ),
       .io_meta_write_valid( prober_io_meta_write_valid ),
       .io_meta_write_bits_idx( prober_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_wb_req_ready( wbArb_io_in_0_ready ),
       .io_wb_req_valid( prober_io_wb_req_valid ),
       .io_wb_req_bits_tag( prober_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( prober_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_way_en( s2_tag_match_way ),
       .io_mshr_rdy( mshrs_io_probe_rdy ),
       .io_line_state_state( s2_hit_state_state )
  );
  `ifndef SYNTHESIS
    assign prober.io_req_bits_client_xact_id = {1{$random}};
  `endif
  MSHRFile mshrs(.clk(clk), .reset(reset),
       .io_req_ready( mshrs_io_req_ready ),
       .io_req_valid( T309 ),
       .io_req_bits_kill( s2_req_kill ),
       .io_req_bits_typ( s2_req_typ ),
       .io_req_bits_phys( s2_req_phys ),
       .io_req_bits_addr( s2_req_addr ),
       .io_req_bits_data( s2_req_data ),
       .io_req_bits_tag( s2_req_tag ),
       .io_req_bits_cmd( s2_req_cmd ),
       .io_req_bits_tag_match( T77 ),
       .io_req_bits_old_meta_tag( T298 ),
       .io_req_bits_old_meta_coh_state( T295 ),
       .io_req_bits_way_en( T290 ),
       .io_secondary_miss( mshrs_io_secondary_miss ),
       .io_mem_req_ready( T289 ),
       .io_mem_req_valid( mshrs_io_mem_req_valid ),
       .io_mem_req_bits_addr( mshrs_io_mem_req_bits_addr ),
       .io_mem_req_bits_client_xact_id( mshrs_io_mem_req_bits_client_xact_id ),
       .io_mem_req_bits_data( mshrs_io_mem_req_bits_data ),
       .io_mem_req_bits_a_type( mshrs_io_mem_req_bits_a_type ),
       .io_mem_req_bits_write_mask( mshrs_io_mem_req_bits_write_mask ),
       .io_mem_req_bits_subword_addr( mshrs_io_mem_req_bits_subword_addr ),
       .io_mem_req_bits_atomic_opcode( mshrs_io_mem_req_bits_atomic_opcode ),
       .io_mem_resp_way_en( mshrs_io_mem_resp_way_en ),
       .io_mem_resp_addr( mshrs_io_mem_resp_addr ),
       //.io_mem_resp_wmask(  )
       //.io_mem_resp_data(  )
       .io_meta_read_ready( metaReadArb_io_in_1_ready ),
       .io_meta_read_valid( mshrs_io_meta_read_valid ),
       .io_meta_read_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_meta_read_bits_tag(  )
       .io_meta_write_ready( metaWriteArb_io_in_0_ready ),
       .io_meta_write_valid( mshrs_io_meta_write_valid ),
       .io_meta_write_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_meta_write_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_meta_write_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_meta_write_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_replay_ready( readArb_io_in_1_ready ),
       .io_replay_valid( mshrs_io_replay_valid ),
       .io_replay_bits_kill( mshrs_io_replay_bits_kill ),
       .io_replay_bits_typ( mshrs_io_replay_bits_typ ),
       .io_replay_bits_phys( mshrs_io_replay_bits_phys ),
       .io_replay_bits_addr( mshrs_io_replay_bits_addr ),
       .io_replay_bits_data( mshrs_io_replay_bits_data ),
       .io_replay_bits_tag( mshrs_io_replay_bits_tag ),
       .io_replay_bits_cmd( mshrs_io_replay_bits_cmd ),
       //.io_replay_bits_sdq_id(  )
       .io_mem_grant_valid( T288 ),
       .io_mem_grant_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       .io_mem_grant_bits_header_dst( FlowThroughSerializer_io_out_bits_header_dst ),
       .io_mem_grant_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( FlowThroughSerializer_io_out_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type ),
       .io_mem_finish_ready( io_mem_finish_ready ),
       .io_mem_finish_valid( mshrs_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( mshrs_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( mshrs_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( mshrs_io_mem_finish_bits_payload_master_xact_id ),
       .io_wb_req_ready( wbArb_io_in_1_ready ),
       .io_wb_req_valid( mshrs_io_wb_req_valid ),
       .io_wb_req_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_wb_req_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_wb_req_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_wb_req_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_wb_req_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_wb_req_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_probe_rdy( mshrs_io_probe_rdy ),
       .io_fence_rdy( mshrs_io_fence_rdy )
  );
  TLB dtlb(.clk(clk), .reset(reset),
       .io_req_ready( dtlb_io_req_ready ),
       .io_req_valid( T275 ),
       .io_req_bits_asid( 7'h0 ),
       .io_req_bits_vpn( T274 ),
       .io_req_bits_passthrough( s1_req_phys ),
       .io_req_bits_instruction( 1'h0 ),
       .io_resp_miss( dtlb_io_resp_miss ),
       //.io_resp_hit_idx(  )
       .io_resp_ppn( dtlb_io_resp_ppn ),
       .io_resp_xcpt_ld( dtlb_io_resp_xcpt_ld ),
       .io_resp_xcpt_st( dtlb_io_resp_xcpt_st ),
       //.io_resp_xcpt_if(  )
       .io_ptw_req_ready( io_cpu_ptw_req_ready ),
       .io_ptw_req_valid( dtlb_io_ptw_req_valid ),
       .io_ptw_req_bits( dtlb_io_ptw_req_bits ),
       .io_ptw_resp_valid( io_cpu_ptw_resp_valid ),
       .io_ptw_resp_bits_error( io_cpu_ptw_resp_bits_error ),
       .io_ptw_resp_bits_ppn( io_cpu_ptw_resp_bits_ppn ),
       .io_ptw_resp_bits_perm( io_cpu_ptw_resp_bits_perm ),
       .io_ptw_status_ip( io_cpu_ptw_status_ip ),
       .io_ptw_status_im( io_cpu_ptw_status_im ),
       .io_ptw_status_zero( io_cpu_ptw_status_zero ),
       .io_ptw_status_er( io_cpu_ptw_status_er ),
       .io_ptw_status_vm( io_cpu_ptw_status_vm ),
       .io_ptw_status_s64( io_cpu_ptw_status_s64 ),
       .io_ptw_status_u64( io_cpu_ptw_status_u64 ),
       .io_ptw_status_ef( io_cpu_ptw_status_ef ),
       .io_ptw_status_pei( io_cpu_ptw_status_pei ),
       .io_ptw_status_ei( io_cpu_ptw_status_ei ),
       .io_ptw_status_ps( io_cpu_ptw_status_ps ),
       .io_ptw_status_s( io_cpu_ptw_status_s ),
       .io_ptw_invalidate( io_cpu_ptw_invalidate ),
       .io_ptw_sret( io_cpu_ptw_sret )
  );
  MetadataArray meta(.clk(clk), .reset(reset),
       .io_read_ready( meta_io_read_ready ),
       .io_read_valid( metaReadArb_io_out_valid ),
       .io_read_bits_idx( metaReadArb_io_out_bits_idx ),
       .io_write_ready( meta_io_write_ready ),
       .io_write_valid( metaWriteArb_io_out_valid ),
       .io_write_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_write_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_write_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_write_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state ),
       .io_resp_0_tag( meta_io_resp_0_tag ),
       .io_resp_0_coh_state( meta_io_resp_0_coh_state )
  );
  Arbiter_7 metaReadArb(
       .io_in_4_ready( metaReadArb_io_in_4_ready ),
       .io_in_4_valid( io_cpu_req_valid ),
       .io_in_4_bits_idx( T266 ),
       .io_in_3_ready( metaReadArb_io_in_3_ready ),
       .io_in_3_valid( wb_io_meta_read_valid ),
       .io_in_3_bits_idx( wb_io_meta_read_bits_idx ),
       .io_in_2_ready( metaReadArb_io_in_2_ready ),
       .io_in_2_valid( prober_io_meta_read_valid ),
       .io_in_2_bits_idx( prober_io_meta_read_bits_idx ),
       .io_in_1_ready( metaReadArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_meta_read_valid ),
       .io_in_1_bits_idx( mshrs_io_meta_read_bits_idx ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_idx( T264 ),
       .io_out_ready( meta_io_read_ready ),
       .io_out_valid( metaReadArb_io_out_valid ),
       .io_out_bits_idx( metaReadArb_io_out_bits_idx )
       //.io_chosen(  )
  );
  Arbiter_1 metaWriteArb(
       .io_in_1_ready( metaWriteArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_meta_write_valid ),
       .io_in_1_bits_idx( prober_io_meta_write_bits_idx ),
       .io_in_1_bits_way_en( prober_io_meta_write_bits_way_en ),
       .io_in_1_bits_data_tag( prober_io_meta_write_bits_data_tag ),
       .io_in_1_bits_data_coh_state( prober_io_meta_write_bits_data_coh_state ),
       .io_in_0_ready( metaWriteArb_io_in_0_ready ),
       .io_in_0_valid( mshrs_io_meta_write_valid ),
       .io_in_0_bits_idx( mshrs_io_meta_write_bits_idx ),
       .io_in_0_bits_way_en( mshrs_io_meta_write_bits_way_en ),
       .io_in_0_bits_data_tag( mshrs_io_meta_write_bits_data_tag ),
       .io_in_0_bits_data_coh_state( mshrs_io_meta_write_bits_data_coh_state ),
       .io_out_ready( meta_io_write_ready ),
       .io_out_valid( metaWriteArb_io_out_valid ),
       .io_out_bits_idx( metaWriteArb_io_out_bits_idx ),
       .io_out_bits_way_en( metaWriteArb_io_out_bits_way_en ),
       .io_out_bits_data_tag( metaWriteArb_io_out_bits_data_tag ),
       .io_out_bits_data_coh_state( metaWriteArb_io_out_bits_data_coh_state )
       //.io_chosen(  )
  );
  DataArray data(.clk(clk),
       //.io_read_ready(  )
       .io_read_valid( readArb_io_out_valid ),
       .io_read_bits_way_en( readArb_io_out_bits_way_en ),
       .io_read_bits_addr( readArb_io_out_bits_addr ),
       .io_write_ready( data_io_write_ready ),
       .io_write_valid( writeArb_io_out_valid ),
       .io_write_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_write_bits_addr( writeArb_io_out_bits_addr ),
       .io_write_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_write_bits_data( T260 ),
       .io_resp_0( data_io_resp_0 )
  );
  Arbiter_8 readArb(
       .io_in_3_ready( readArb_io_in_3_ready ),
       .io_in_3_valid( io_cpu_req_valid ),
       .io_in_3_bits_way_en( 1'h1 ),
       .io_in_3_bits_addr( T259 ),
       .io_in_2_ready( readArb_io_in_2_ready ),
       .io_in_2_valid( wb_io_data_req_valid ),
       .io_in_2_bits_way_en( wb_io_data_req_bits_way_en ),
       .io_in_2_bits_addr( wb_io_data_req_bits_addr ),
       .io_in_1_ready( readArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_replay_valid ),
       .io_in_1_bits_way_en( 1'h1 ),
       .io_in_1_bits_addr( T258 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s2_recycle ),
       .io_in_0_bits_way_en( 1'h1 ),
       .io_in_0_bits_addr( T257 ),
       .io_out_ready( T255 ),
       .io_out_valid( readArb_io_out_valid ),
       .io_out_bits_way_en( readArb_io_out_bits_way_en ),
       .io_out_bits_addr( readArb_io_out_bits_addr )
       //.io_chosen(  )
  );
  Arbiter_9 writeArb(
       .io_in_1_ready( writeArb_io_in_1_ready ),
       .io_in_1_valid( T251 ),
       .io_in_1_bits_way_en( mshrs_io_mem_resp_way_en ),
       .io_in_1_bits_addr( mshrs_io_mem_resp_addr ),
       .io_in_1_bits_wmask( 2'h3 ),
       .io_in_1_bits_data( T250 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( s3_valid ),
       .io_in_0_bits_way_en( s3_way ),
       .io_in_0_bits_addr( T248 ),
       .io_in_0_bits_wmask( T245 ),
       .io_in_0_bits_data( T244 ),
       .io_out_ready( data_io_write_ready ),
       .io_out_valid( writeArb_io_out_valid ),
       .io_out_bits_way_en( writeArb_io_out_bits_way_en ),
       .io_out_bits_addr( writeArb_io_out_bits_addr ),
       .io_out_bits_wmask( writeArb_io_out_bits_wmask ),
       .io_out_bits_data( writeArb_io_out_bits_data )
       //.io_chosen(  )
  );
  AMOALU amoalu(
       .io_addr( T243 ),
       .io_cmd( T242 ),
       .io_typ( s2_req_typ ),
       .io_lhs( T103 ),
       .io_rhs( s2_req_data ),
       .io_out( amoalu_io_out )
  );
  Arbiter_10 releaseArb(
       .io_in_1_ready( releaseArb_io_in_1_ready ),
       .io_in_1_valid( prober_io_rep_valid ),
       .io_in_1_bits_addr( prober_io_rep_bits_addr ),
       .io_in_1_bits_client_xact_id( prober_io_rep_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( prober_io_rep_bits_master_xact_id ),
       .io_in_1_bits_data( prober_io_rep_bits_data ),
       .io_in_1_bits_r_type( prober_io_rep_bits_r_type ),
       .io_in_0_ready( releaseArb_io_in_0_ready ),
       .io_in_0_valid( wb_io_release_valid ),
       .io_in_0_bits_addr( wb_io_release_bits_addr ),
       .io_in_0_bits_client_xact_id( wb_io_release_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( wb_io_release_bits_master_xact_id ),
       .io_in_0_bits_data( wb_io_release_bits_data ),
       .io_in_0_bits_r_type( wb_io_release_bits_r_type ),
       .io_out_ready( T5 ),
       .io_out_valid( releaseArb_io_out_valid ),
       .io_out_bits_addr( releaseArb_io_out_bits_addr ),
       .io_out_bits_client_xact_id( releaseArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( releaseArb_io_out_bits_master_xact_id ),
       .io_out_bits_data( releaseArb_io_out_bits_data ),
       .io_out_bits_r_type( releaseArb_io_out_bits_r_type )
       //.io_chosen(  )
  );
  FlowThroughSerializer_1 FlowThroughSerializer(.clk(clk), .reset(reset),
       .io_in_ready( FlowThroughSerializer_io_in_ready ),
       .io_in_valid( io_mem_grant_valid ),
       .io_in_bits_header_src( io_mem_grant_bits_header_src ),
       .io_in_bits_header_dst( io_mem_grant_bits_header_dst ),
       .io_in_bits_payload_data( io_mem_grant_bits_payload_data ),
       .io_in_bits_payload_client_xact_id( io_mem_grant_bits_payload_client_xact_id ),
       .io_in_bits_payload_master_xact_id( io_mem_grant_bits_payload_master_xact_id ),
       .io_in_bits_payload_g_type( io_mem_grant_bits_payload_g_type ),
       .io_out_ready( T0 ),
       .io_out_valid( FlowThroughSerializer_io_out_valid ),
       .io_out_bits_header_src( FlowThroughSerializer_io_out_bits_header_src ),
       .io_out_bits_header_dst( FlowThroughSerializer_io_out_bits_header_dst ),
       .io_out_bits_payload_data( FlowThroughSerializer_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( FlowThroughSerializer_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( FlowThroughSerializer_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( FlowThroughSerializer_io_out_bits_payload_g_type )
       //.io_cnt(  )
       //.io_done(  )
  );
  Arbiter_4 wbArb(
       .io_in_1_ready( wbArb_io_in_1_ready ),
       .io_in_1_valid( mshrs_io_wb_req_valid ),
       .io_in_1_bits_tag( mshrs_io_wb_req_bits_tag ),
       .io_in_1_bits_idx( mshrs_io_wb_req_bits_idx ),
       .io_in_1_bits_way_en( mshrs_io_wb_req_bits_way_en ),
       .io_in_1_bits_client_xact_id( mshrs_io_wb_req_bits_client_xact_id ),
       .io_in_1_bits_master_xact_id( mshrs_io_wb_req_bits_master_xact_id ),
       .io_in_1_bits_r_type( mshrs_io_wb_req_bits_r_type ),
       .io_in_0_ready( wbArb_io_in_0_ready ),
       .io_in_0_valid( prober_io_wb_req_valid ),
       .io_in_0_bits_tag( prober_io_wb_req_bits_tag ),
       .io_in_0_bits_idx( prober_io_wb_req_bits_idx ),
       .io_in_0_bits_way_en( prober_io_wb_req_bits_way_en ),
       .io_in_0_bits_client_xact_id( prober_io_wb_req_bits_client_xact_id ),
       .io_in_0_bits_master_xact_id( prober_io_wb_req_bits_master_xact_id ),
       .io_in_0_bits_r_type( prober_io_wb_req_bits_r_type ),
       .io_out_ready( wb_io_req_ready ),
       .io_out_valid( wbArb_io_out_valid ),
       .io_out_bits_tag( wbArb_io_out_bits_tag ),
       .io_out_bits_idx( wbArb_io_out_bits_idx ),
       .io_out_bits_way_en( wbArb_io_out_bits_way_en ),
       .io_out_bits_client_xact_id( wbArb_io_out_bits_client_xact_id ),
       .io_out_bits_master_xact_id( wbArb_io_out_bits_master_xact_id ),
       .io_out_bits_r_type( wbArb_io_out_bits_r_type )
       //.io_chosen(  )
  );

  always @(posedge clk) begin
    if(T101) begin
      s2_req_data <= s1_req_data;
    end else if(T11) begin
      s2_req_data <= T8;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T10;
    end
    if(s2_recycle) begin
      s1_req_cmd <= s2_req_cmd;
    end else if(mshrs_io_replay_valid) begin
      s1_req_cmd <= mshrs_io_replay_bits_cmd;
    end else if(io_cpu_req_valid) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if(s1_clk_en) begin
      s2_req_cmd <= s1_req_cmd;
    end
    s1_clk_en <= metaReadArb_io_out_valid;
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else if(T93) begin
      s2_recycle_next <= T21;
    end
    if(s1_clk_en) begin
      s2_req_addr <= T29;
    end
    if(s2_recycle) begin
      s1_req_addr <= s2_req_addr;
    end else if(mshrs_io_replay_valid) begin
      s1_req_addr <= mshrs_io_replay_bits_addr;
    end else if(prober_io_meta_read_valid) begin
      s1_req_addr <= T39;
    end else if(wb_io_meta_read_valid) begin
      s1_req_addr <= T36;
    end else if(io_cpu_req_valid) begin
      s1_req_addr <= io_cpu_req_bits_addr;
    end
    if(s1_clk_en) begin
      s2_hit_state_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_tag_match_way <= s1_tag_match_way;
    end
    if(reset) begin
      R86 <= 1'h0;
    end else begin
      R86 <= s1_replay;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T91;
    end
    if(s2_recycle) begin
      s1_req_data <= s2_req_data;
    end else if(mshrs_io_replay_valid) begin
      s1_req_data <= mshrs_io_replay_bits_data;
    end else if(io_cpu_req_valid) begin
      s1_req_data <= io_cpu_req_bits_data;
    end
    if(s1_clk_en) begin
      s1_recycled <= s2_recycle;
    end
    R109 <= T110;
    if(T114) begin
      R116 <= T118;
    end
    if(T217) begin
      s2_store_bypass_data <= T122;
    end
    if(T142) begin
      s4_req_data <= s3_req_data;
    end
    s3_req_data <= T125;
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T144;
    end
    if(T159) begin
      lrsc_addr <= T158;
    end
    if(T173) begin
      s2_nack_hit <= s1_nack;
    end
    if(reset) begin
      lrsc_count <= 5'h0;
    end else if(io_cpu_ptw_sret) begin
      lrsc_count <= 5'h0;
    end else if(T183) begin
      lrsc_count <= 5'h0;
    end else if(T181) begin
      lrsc_count <= 5'h1f;
    end else if(T174) begin
      lrsc_count <= T180;
    end
    if(T129) begin
      s3_req_cmd <= s2_req_cmd;
    end
    if(T129) begin
      s3_req_addr <= s2_req_addr;
    end
    if(T142) begin
      s4_req_cmd <= s3_req_cmd;
    end
    if(T142) begin
      s4_req_addr <= s3_req_addr;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(T217) begin
      s2_store_bypass <= 1'h1;
    end else if(s1_clk_en) begin
      s2_store_bypass <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_req_typ <= s1_req_typ;
    end
    if(s2_recycle) begin
      s1_req_typ <= s2_req_typ;
    end else if(mshrs_io_replay_valid) begin
      s1_req_typ <= mshrs_io_replay_bits_typ;
    end else if(io_cpu_req_valid) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if(T129) begin
      s3_way <= s2_tag_match_way;
    end
    if(s2_recycle) begin
      s1_req_phys <= s2_req_phys;
    end else if(mshrs_io_replay_valid) begin
      s1_req_phys <= mshrs_io_replay_bits_phys;
    end else if(prober_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(wb_io_meta_read_valid) begin
      s1_req_phys <= 1'h1;
    end else if(io_cpu_req_valid) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    if(s1_clk_en) begin
      s2_req_phys <= s1_req_phys;
    end
    if(s1_clk_en) begin
      R292 <= 1'h0;
    end
    if(s1_clk_en) begin
      s2_repl_meta_coh_state <= meta_io_resp_0_coh_state;
    end
    if(s1_clk_en) begin
      s2_repl_meta_tag <= meta_io_resp_0_tag;
    end
    if(s1_clk_en) begin
      s2_req_tag <= s1_req_tag;
    end
    if(s2_recycle) begin
      s1_req_tag <= s2_req_tag;
    end else if(mshrs_io_replay_valid) begin
      s1_req_tag <= mshrs_io_replay_bits_tag;
    end else if(io_cpu_req_valid) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if(s1_clk_en) begin
      s2_req_kill <= s1_req_kill;
    end
    if(s2_recycle) begin
      s1_req_kill <= s2_req_kill;
    end else if(mshrs_io_replay_valid) begin
      s1_req_kill <= mshrs_io_replay_bits_kill;
    end else if(io_cpu_req_valid) begin
      s1_req_kill <= io_cpu_req_bits_kill;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T458;
    end
  end
endmodule

module RRArbiter_0(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [29:0] io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [29:0] io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output[29:0] io_out_bits,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[29:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits = T9;
  assign T9 = T10 ? io_in_1_bits : io_in_0_bits;
  assign T10 = T0;
  assign io_out_valid = T11;
  assign T11 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T12;
  assign T12 = T13 & io_out_ready;
  assign T13 = T20 | T14;
  assign T14 = T15 ^ 1'h1;
  assign T15 = T18 | T16;
  assign T16 = io_in_1_valid & T17;
  assign T17 = R5 < 1'h1;
  assign T18 = io_in_0_valid & T19;
  assign T19 = R5 < 1'h0;
  assign T20 = R5 < 1'h0;
  assign io_in_1_ready = T21;
  assign T21 = T22 & io_out_ready;
  assign T22 = T26 | T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = T25 | io_in_0_valid;
  assign T25 = T18 | T16;
  assign T26 = T28 & T27;
  assign T27 = R5 < 1'h1;
  assign T28 = T18 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module PTW(input clk, input reset,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input [29:0] io_requestor_1_req_bits,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_error,
    output[18:0] io_requestor_1_resp_bits_ppn,
    output[5:0] io_requestor_1_resp_bits_perm,
    output[7:0] io_requestor_1_status_ip,
    output[7:0] io_requestor_1_status_im,
    output[6:0] io_requestor_1_status_zero,
    output io_requestor_1_status_er,
    output io_requestor_1_status_vm,
    output io_requestor_1_status_s64,
    output io_requestor_1_status_u64,
    output io_requestor_1_status_ef,
    output io_requestor_1_status_pei,
    output io_requestor_1_status_ei,
    output io_requestor_1_status_ps,
    output io_requestor_1_status_s,
    output io_requestor_1_invalidate,
    output io_requestor_1_sret,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input [29:0] io_requestor_0_req_bits,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_error,
    output[18:0] io_requestor_0_resp_bits_ppn,
    output[5:0] io_requestor_0_resp_bits_perm,
    output[7:0] io_requestor_0_status_ip,
    output[7:0] io_requestor_0_status_im,
    output[6:0] io_requestor_0_status_zero,
    output io_requestor_0_status_er,
    output io_requestor_0_status_vm,
    output io_requestor_0_status_s64,
    output io_requestor_0_status_u64,
    output io_requestor_0_status_ef,
    output io_requestor_0_status_pei,
    output io_requestor_0_status_ei,
    output io_requestor_0_status_ps,
    output io_requestor_0_status_s,
    output io_requestor_0_invalidate,
    output io_requestor_0_sret,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    //output[63:0] io_mem_req_bits_data
    //output[7:0] io_mem_req_bits_tag
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    //input  io_mem_ptw_req_valid
    //input [29:0] io_mem_ptw_req_bits
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered,
    input [31:0] io_dpath_ptbr,
    input  io_dpath_invalidate,
    input  io_dpath_sret,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s
);

  wire T0;
  reg [2:0] state;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire T10;
  wire arb_io_out_valid;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg [1:0] count;
  wire[1:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire T29;
  wire T30;
  wire[43:0] T31;
  wire[31:0] T32;
  wire[28:0] T33;
  wire[28:0] T34;
  wire[9:0] T35;
  wire[9:0] T36;
  wire[9:0] T37;
  wire[9:0] T38;
  reg [29:0] r_req_vpn;
  wire[29:0] T39;
  wire[29:0] arb_io_out_bits;
  wire T40;
  wire[9:0] T41;
  wire[19:0] T42;
  wire T43;
  wire[1:0] T44;
  wire[9:0] T45;
  wire[29:0] T46;
  wire T47;
  wire[18:0] T48;
  reg [63:0] r_pte;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  wire[31:0] T52;
  wire[12:0] T53;
  wire[18:0] T54;
  wire T55;
  wire[5:0] T56;
  wire[18:0] T57;
  wire[30:0] T58;
  wire[30:0] T59;
  wire[30:0] T60;
  wire[30:0] T61;
  wire[19:0] T62;
  wire[10:0] T63;
  wire[30:0] r_resp_ppn;
  wire[30:0] T64;
  wire[9:0] T65;
  wire[20:0] T66;
  wire T67;
  wire[1:0] T68;
  wire T69;
  wire resp_err;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  r_req_dest;
  wire T74;
  wire arb_io_chosen;
  wire resp_val;
  wire T75;
  wire T76;
  wire arb_io_in_0_ready;
  wire[5:0] T77;
  wire[18:0] T78;
  wire[30:0] T79;
  wire T80;
  wire T81;
  wire arb_io_in_1_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    count = {1{$random}};
    r_req_vpn = {1{$random}};
    r_pte = {2{$random}};
    r_req_dest = {1{$random}};
  end
`endif

  assign T0 = state == 3'h0;
  assign T1 = reset ? 3'h0 : T2;
  assign T2 = T30 ? 3'h0 : T3;
  assign T3 = T29 ? 3'h0 : T4;
  assign T4 = T22 ? 3'h1 : T5;
  assign T5 = T17 ? 3'h3 : T6;
  assign T6 = T16 ? 3'h4 : T7;
  assign T7 = T14 ? 3'h1 : T8;
  assign T8 = T12 ? 3'h2 : T9;
  assign T9 = T10 ? 3'h1 : state;
  assign T10 = T11 & arb_io_out_valid;
  assign T11 = 3'h0 == state;
  assign T12 = T13 & io_mem_req_ready;
  assign T13 = 3'h1 == state;
  assign T14 = T15 & io_mem_resp_bits_nack;
  assign T15 = 3'h2 == state;
  assign T16 = T15 & io_mem_resp_valid;
  assign T17 = T20 & T18;
  assign T18 = T19 ^ 1'h1;
  assign T19 = io_mem_resp_bits_data[1'h1:1'h1];
  assign T20 = T16 & T21;
  assign T21 = io_mem_resp_bits_data[1'h0:1'h0];
  assign T22 = T20 & T23;
  assign T23 = T28 & T24;
  assign T24 = count < 2'h2;
  assign T25 = T22 ? T27 : T26;
  assign T26 = T11 ? 2'h0 : count;
  assign T27 = count + 2'h1;
  assign T28 = T18 ^ 1'h1;
  assign T29 = 3'h3 == state;
  assign T30 = 3'h4 == state;
  assign io_mem_req_bits_cmd = 5'h0;
  assign io_mem_req_bits_addr = T31;
  assign T31 = {12'h0, T32};
  assign T32 = T33 << 2'h3;
  assign T33 = T34;
  assign T34 = {T48, T35};
  assign T35 = T47 ? T45 : T36;
  assign T36 = T43 ? T41 : T37;
  assign T37 = T38[4'h9:1'h0];
  assign T38 = r_req_vpn >> 5'h14;
  assign T39 = T40 ? arb_io_out_bits : r_req_vpn;
  assign T40 = T0 & arb_io_out_valid;
  assign T41 = T42[4'h9:1'h0];
  assign T42 = r_req_vpn >> 4'ha;
  assign T43 = T44[1'h0:1'h0];
  assign T44 = count;
  assign T45 = T46[4'h9:1'h0];
  assign T46 = r_req_vpn >> 1'h0;
  assign T47 = T44[1'h1:1'h1];
  assign T48 = r_pte[5'h1f:4'hd];
  assign T49 = io_mem_resp_valid ? io_mem_resp_bits_data : T50;
  assign T50 = T40 ? T51 : r_pte;
  assign T51 = {32'h0, T52};
  assign T52 = {T54, T53};
  assign T53 = io_mem_resp_bits_data[4'hc:1'h0];
  assign T54 = io_dpath_ptbr[5'h1f:4'hd];
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_kill = 1'h0;
  assign io_mem_req_valid = T55;
  assign T55 = state == 3'h1;
  assign io_requestor_0_sret = io_dpath_sret;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_s = io_dpath_status_s;
  assign io_requestor_0_status_ps = io_dpath_status_ps;
  assign io_requestor_0_status_ei = io_dpath_status_ei;
  assign io_requestor_0_status_pei = io_dpath_status_pei;
  assign io_requestor_0_status_ef = io_dpath_status_ef;
  assign io_requestor_0_status_u64 = io_dpath_status_u64;
  assign io_requestor_0_status_s64 = io_dpath_status_s64;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_er = io_dpath_status_er;
  assign io_requestor_0_status_zero = io_dpath_status_zero;
  assign io_requestor_0_status_im = io_dpath_status_im;
  assign io_requestor_0_status_ip = io_dpath_status_ip;
  assign io_requestor_0_resp_bits_perm = T56;
  assign T56 = r_pte[4'h8:2'h3];
  assign io_requestor_0_resp_bits_ppn = T57;
  assign T57 = T58[5'h12:1'h0];
  assign T58 = T59;
  assign T59 = T69 ? r_resp_ppn : T60;
  assign T60 = T67 ? T64 : T61;
  assign T61 = {T63, T62};
  assign T62 = r_req_vpn[5'h13:1'h0];
  assign T63 = r_resp_ppn >> 5'h14;
  assign r_resp_ppn = io_mem_req_bits_addr >> 4'hd;
  assign T64 = {T66, T65};
  assign T65 = r_req_vpn[4'h9:1'h0];
  assign T66 = r_resp_ppn >> 4'ha;
  assign T67 = T68[1'h0:1'h0];
  assign T68 = count;
  assign T69 = T68[1'h1:1'h1];
  assign io_requestor_0_resp_bits_error = resp_err;
  assign resp_err = T71 | T70;
  assign T70 = state == 3'h2;
  assign T71 = state == 3'h4;
  assign io_requestor_0_resp_valid = T72;
  assign T72 = resp_val & T73;
  assign T73 = r_req_dest == 1'h0;
  assign T74 = T40 ? arb_io_chosen : r_req_dest;
  assign resp_val = T76 | T75;
  assign T75 = state == 3'h4;
  assign T76 = state == 3'h3;
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_1_sret = io_dpath_sret;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_s = io_dpath_status_s;
  assign io_requestor_1_status_ps = io_dpath_status_ps;
  assign io_requestor_1_status_ei = io_dpath_status_ei;
  assign io_requestor_1_status_pei = io_dpath_status_pei;
  assign io_requestor_1_status_ef = io_dpath_status_ef;
  assign io_requestor_1_status_u64 = io_dpath_status_u64;
  assign io_requestor_1_status_s64 = io_dpath_status_s64;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_er = io_dpath_status_er;
  assign io_requestor_1_status_zero = io_dpath_status_zero;
  assign io_requestor_1_status_im = io_dpath_status_im;
  assign io_requestor_1_status_ip = io_dpath_status_ip;
  assign io_requestor_1_resp_bits_perm = T77;
  assign T77 = r_pte[4'h8:2'h3];
  assign io_requestor_1_resp_bits_ppn = T78;
  assign T78 = T79[5'h12:1'h0];
  assign T79 = T59;
  assign io_requestor_1_resp_bits_error = resp_err;
  assign io_requestor_1_resp_valid = T80;
  assign T80 = resp_val & T81;
  assign T81 = r_req_dest == 1'h1;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  RRArbiter_0 arb(.clk(clk), .reset(reset),
       .io_in_1_ready( arb_io_in_1_ready ),
       .io_in_1_valid( io_requestor_1_req_valid ),
       .io_in_1_bits( io_requestor_1_req_bits ),
       .io_in_0_ready( arb_io_in_0_ready ),
       .io_in_0_valid( io_requestor_0_req_valid ),
       .io_in_0_bits( io_requestor_0_req_bits ),
       .io_out_ready( T0 ),
       .io_out_valid( arb_io_out_valid ),
       .io_out_bits( arb_io_out_bits ),
       .io_chosen( arb_io_chosen )
  );

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T30) begin
      state <= 3'h0;
    end else if(T29) begin
      state <= 3'h0;
    end else if(T22) begin
      state <= 3'h1;
    end else if(T17) begin
      state <= 3'h3;
    end else if(T16) begin
      state <= 3'h4;
    end else if(T14) begin
      state <= 3'h1;
    end else if(T12) begin
      state <= 3'h2;
    end else if(T10) begin
      state <= 3'h1;
    end
    if(T22) begin
      count <= T27;
    end else if(T11) begin
      count <= 2'h0;
    end
    if(T40) begin
      r_req_vpn <= arb_io_out_bits;
    end
    if(io_mem_resp_valid) begin
      r_pte <= io_mem_resp_bits_data;
    end else if(T40) begin
      r_pte <= T51;
    end
    if(T40) begin
      r_req_dest <= arb_io_chosen;
    end
  end
endmodule

module Control(input clk, input reset,
    output[2:0] io_dpath_sel_pc,
    output io_dpath_killd,
    output io_dpath_ren_1,
    output io_dpath_ren_0,
    output[2:0] io_dpath_sel_alu2,
    output[1:0] io_dpath_sel_alu1,
    output[2:0] io_dpath_sel_imm,
    output io_dpath_fn_dw,
    output[3:0] io_dpath_fn_alu,
    output io_dpath_div_mul_val,
    output io_dpath_div_mul_kill,
    //output io_dpath_div_val
    //output io_dpath_div_kill
    output[2:0] io_dpath_csr,
    output io_dpath_sret,
    output io_dpath_mem_load,
    output io_dpath_wb_load,
    output io_dpath_ex_fp_val,
    output io_dpath_mem_fp_val,
    output io_dpath_ex_wen,
    output io_dpath_ex_valid,
    output io_dpath_mem_jalr,
    output io_dpath_mem_branch,
    output io_dpath_mem_wen,
    output io_dpath_wb_wen,
    output[2:0] io_dpath_ex_mem_type,
    output io_dpath_ex_rs2_val,
    output io_dpath_ex_rocc_val,
    output io_dpath_mem_rocc_val,
    output io_dpath_bypass_1,
    output io_dpath_bypass_0,
    output[1:0] io_dpath_bypass_src_1,
    output[1:0] io_dpath_bypass_src_0,
    output io_dpath_ll_ready,
    output io_dpath_retire,
    output io_dpath_exception,
    output[63:0] io_dpath_cause,
    output io_dpath_badvaddr_wen,
    input [31:0] io_dpath_inst,
    //input  io_dpath_jalr_eq
    input  io_dpath_mem_br_taken,
    input  io_dpath_mem_misprediction,
    input  io_dpath_div_mul_rdy,
    input  io_dpath_ll_wen,
    input [4:0] io_dpath_ll_waddr,
    input [4:0] io_dpath_ex_waddr,
    input  io_dpath_mem_rs1_ra,
    input [4:0] io_dpath_mem_waddr,
    input [4:0] io_dpath_wb_waddr,
    input [7:0] io_dpath_status_ip,
    input [7:0] io_dpath_status_im,
    input [6:0] io_dpath_status_zero,
    input  io_dpath_status_er,
    input  io_dpath_status_vm,
    input  io_dpath_status_s64,
    input  io_dpath_status_u64,
    input  io_dpath_status_ef,
    input  io_dpath_status_pei,
    input  io_dpath_status_ei,
    input  io_dpath_status_ps,
    input  io_dpath_status_s,
    input  io_dpath_fp_sboard_clr,
    input [4:0] io_dpath_fp_sboard_clra,
    input  io_dpath_csr_replay,
    output io_imem_req_valid,
    //output[43:0] io_imem_req_bits_pc
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    //output[42:0] io_imem_btb_update_bits_pc
    //output[42:0] io_imem_btb_update_bits_target
    //output[42:0] io_imem_btb_update_bits_returnAddr
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    //output[43:0] io_dmem_req_bits_addr
    //output[63:0] io_dmem_req_bits_data
    //output[7:0] io_dmem_req_bits_tag
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output io_fpu_valid,
    input  io_fpu_fcsr_rdy,
    input  io_fpu_nack_mem,
    input  io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input  io_fpu_dec_ldst,
    input  io_fpu_dec_wen,
    input  io_fpu_dec_ren1,
    input  io_fpu_dec_ren2,
    input  io_fpu_dec_ren3,
    input  io_fpu_dec_swap23,
    input  io_fpu_dec_single,
    input  io_fpu_dec_fromint,
    input  io_fpu_dec_toint,
    input  io_fpu_dec_fastpipe,
    input  io_fpu_dec_fma,
    input  io_fpu_dec_round,
    input  io_fpu_sboard_set,
    input  io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire T0;
  reg  wb_reg_xcpt;
  wire T1;
  wire T2;
  wire take_pc_wb;
  wire T3;
  reg  wb_reg_sret;
  wire T4;
  wire T5;
  wire T6;
  reg  mem_reg_replay;
  wire T7;
  wire replay_ex;
  wire replay_ex_other;
  reg  mem_reg_replay_next;
  wire T8;
  reg  ex_reg_replay_next;
  wire T9;
  wire T10;
  wire id_csr_flush;
  wire T11;
  wire T12;
  wire T13;
  wire[11:0] T14;
  wire[11:0] T15;
  wire T16;
  wire[11:0] T17;
  wire T18;
  wire id_csr_wen;
  wire T19;
  wire T20;
  wire T21;
  wire[1:0] T22;
  wire T23;
  wire[31:0] T24;
  wire T25;
  wire[31:0] T26;
  wire T27;
  wire T28;
  wire[4:0] T29;
  wire T30;
  wire T31;
  wire[31:0] T32;
  wire ctrl_killd;
  wire T33;
  wire ctrl_draind;
  wire id_interrupt;
  wire id_interrupt_unmasked;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire ctrl_stalld;
  wire id_do_fence;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[31:0] T70;
  wire T71;
  wire T72;
  wire[31:0] T73;
  wire T74;
  wire T75;
  wire[31:0] T76;
  wire T77;
  wire T78;
  wire[31:0] T79;
  wire T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire[31:0] T87;
  reg  id_reg_fence;
  wire T88;
  wire T89;
  wire T90;
  wire id_mem_busy;
  reg  ex_reg_mem_val;
  wire T91;
  wire T92;
  wire T93;
  wire id_fence_next;
  wire T94;
  wire T95;
  wire T96;
  wire[31:0] T97;
  wire T98;
  wire[31:0] T99;
  wire T100;
  wire T101;
  wire[31:0] T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire id_stall_fpu;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire[4:0] T116;
  wire T117;
  reg [31:0] R118;
  wire[31:0] T119;
  wire[31:0] T120;
  wire[31:0] T121;
  wire[31:0] T122;
  wire[31:0] T123;
  wire[31:0] T124;
  wire[31:0] T125;
  wire T126;
  wire T127;
  wire replay_wb;
  wire T128;
  wire T129;
  reg  wb_reg_rocc_val;
  wire T130;
  reg  mem_reg_rocc_val;
  wire T131;
  reg  ex_reg_rocc_val;
  wire T132;
  wire T133;
  wire ctrl_killx;
  wire T134;
  wire take_pc_mem_wb;
  wire take_pc_mem;
  wire T135;
  reg  mem_reg_jal;
  wire T136;
  reg  ex_reg_jal;
  wire T137;
  wire T138;
  wire[31:0] T139;
  wire T140;
  reg  mem_reg_jalr;
  wire T141;
  reg  ex_reg_jalr;
  wire T142;
  wire T143;
  wire[31:0] T144;
  reg  mem_reg_branch;
  wire T145;
  reg  ex_reg_branch;
  wire T146;
  wire T147;
  wire[31:0] T148;
  wire ctrl_killm;
  wire T149;
  wire fpu_kill_mem;
  reg  mem_reg_fp_val;
  wire T150;
  reg  ex_reg_fp_val;
  wire T151;
  wire T152;
  wire T153;
  wire[31:0] T154;
  wire T155;
  wire[31:0] T156;
  wire T157;
  wire mem_xcpt;
  wire T158;
  reg  mem_reg_mem_val;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  reg  mem_reg_xcpt;
  wire T167;
  wire ex_xcpt;
  wire T168;
  wire T169;
  reg  ex_reg_xcpt;
  wire T170;
  wire id_xcpt;
  wire T171;
  wire[31:0] T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire id_csr_fp;
  wire T177;
  wire[11:0] T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire[31:0] T183;
  wire T184;
  wire id_csr_privileged;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire[1:0] T190;
  wire T191;
  wire T192;
  wire[1:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire[1:0] T198;
  wire T199;
  wire T200;
  wire[1:0] T201;
  wire T202;
  wire T203;
  wire[1:0] T204;
  wire T205;
  wire T206;
  wire id_csr_invalid;
  wire T207;
  reg  T208;
  wire T210;
  wire T211;
  wire T212;
  wire[31:0] T213;
  wire T214;
  wire T215;
  wire[31:0] T216;
  wire T217;
  wire T218;
  wire[31:0] T219;
  wire T220;
  wire T221;
  wire[31:0] T222;
  wire T223;
  wire T224;
  wire[31:0] T225;
  wire T226;
  wire T227;
  wire[31:0] T228;
  wire T229;
  wire T230;
  wire[31:0] T231;
  wire T232;
  wire T233;
  wire[31:0] T234;
  wire T235;
  wire T236;
  wire[31:0] T237;
  wire T238;
  wire T239;
  wire[31:0] T240;
  wire T241;
  wire T242;
  wire[31:0] T243;
  wire T244;
  wire T245;
  wire[31:0] T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire[31:0] T251;
  wire T252;
  wire T253;
  wire[31:0] T254;
  wire T255;
  wire T256;
  wire[31:0] T257;
  wire T258;
  wire T259;
  wire[31:0] T260;
  wire T261;
  wire T262;
  wire[31:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[31:0] T267;
  wire T268;
  wire T269;
  wire T270;
  wire[31:0] T271;
  wire T272;
  wire T273;
  wire[31:0] T274;
  wire T275;
  wire T276;
  wire[31:0] T277;
  wire T278;
  wire T279;
  wire[31:0] T280;
  wire T281;
  wire T282;
  wire[31:0] T283;
  wire T284;
  wire T285;
  wire[31:0] T286;
  wire T287;
  wire T288;
  wire[31:0] T289;
  wire T290;
  wire T291;
  wire[31:0] T292;
  wire T293;
  wire T294;
  wire[31:0] T295;
  wire T296;
  wire T297;
  wire[31:0] T298;
  wire T299;
  wire T300;
  wire[31:0] T301;
  wire T302;
  wire T303;
  wire[31:0] T304;
  wire T305;
  wire T306;
  wire[31:0] T307;
  wire T308;
  wire T309;
  wire[31:0] T310;
  wire T311;
  wire T312;
  reg  ex_reg_xcpt_interrupt;
  wire T313;
  wire T314;
  wire T315;
  reg  mem_reg_xcpt_interrupt;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire killm_common;
  wire T320;
  reg  mem_reg_valid;
  wire T321;
  reg  ex_reg_valid;
  wire T322;
  wire T323;
  wire T324;
  wire dcache_kill_mem;
  reg  mem_reg_wen;
  wire T325;
  reg  ex_reg_wen;
  wire T326;
  wire T327;
  wire T328;
  wire[31:0] T329;
  wire T330;
  wire T331;
  wire[31:0] T332;
  wire T333;
  wire T334;
  wire[31:0] T335;
  wire T336;
  wire T337;
  wire[31:0] T338;
  wire T339;
  wire T340;
  wire[31:0] T341;
  wire T342;
  wire T343;
  wire[31:0] T344;
  wire T345;
  wire[31:0] T346;
  wire replay_wb_common;
  wire T347;
  reg  wb_reg_replay;
  wire T348;
  wire T349;
  wire replay_mem;
  wire T350;
  wire T351;
  wire T352;
  reg  wb_reg_fp_wen;
  wire T353;
  reg  mem_reg_fp_wen;
  wire T354;
  reg  ex_reg_fp_wen;
  wire T355;
  wire T356;
  wire wb_dcache_miss;
  wire T357;
  reg  wb_reg_mem_val;
  wire T358;
  wire[31:0] T359;
  wire[31:0] T360;
  wire[31:0] T361;
  wire[31:0] T362;
  wire T363;
  wire[31:0] T364;
  wire[31:0] T365;
  wire[31:0] T366;
  wire[31:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire[4:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire[4:0] T392;
  wire[4:0] T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire id_sboard_hazard;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire[4:0] T402;
  wire[4:0] T403;
  wire T404;
  wire[31:0] T405;
  wire[31:0] T406;
  wire[31:0] T407;
  wire[31:0] T408;
  reg [31:0] R409;
  wire[31:0] T410;
  wire[31:0] T411;
  wire[31:0] T412;
  wire[31:0] T413;
  wire[31:0] T414;
  wire[31:0] T415;
  wire T416;
  wire wb_set_sboard;
  wire T417;
  reg  wb_reg_div_mul_val;
  wire T418;
  reg  mem_reg_div_mul_val;
  wire T419;
  reg  ex_reg_div_mul_val;
  wire T420;
  wire T421;
  wire T422;
  wire[31:0] T423;
  wire T424;
  wire[31:0] T425;
  wire T426;
  wire id_wen_not0;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire[4:0] T433;
  wire[4:0] T434;
  wire T435;
  wire id_renx2_not0;
  wire T436;
  wire T437;
  wire T438;
  wire[31:0] T439;
  wire T440;
  wire T441;
  wire[31:0] T442;
  wire T443;
  wire[31:0] T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire[4:0] T449;
  wire[4:0] T450;
  wire T451;
  wire id_renx1_not0;
  wire T452;
  wire T453;
  wire T454;
  wire[31:0] T455;
  wire T456;
  wire T457;
  wire[31:0] T458;
  wire T459;
  wire T460;
  wire[31:0] T461;
  wire T462;
  wire T463;
  wire[31:0] T464;
  wire T465;
  wire T466;
  wire[31:0] T467;
  wire T468;
  wire[31:0] T469;
  wire T470;
  wire id_wb_hazard;
  wire T471;
  wire T472;
  reg  wb_reg_fp_val;
  wire T473;
  wire fp_data_hazard_wb;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire data_hazard_wb;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  reg  wb_reg_wen;
  wire T494;
  wire T495;
  wire id_mem_hazard;
  wire T496;
  wire fp_data_hazard_mem;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  reg  mem_reg_slow_bypass;
  wire T514;
  wire ex_slow_bypass;
  wire T515;
  wire T516;
  reg [2:0] ex_reg_mem_type;
  wire[2:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire[1:0] T520;
  wire T521;
  wire[31:0] T522;
  wire T523;
  wire[31:0] T524;
  wire T525;
  wire[31:0] T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  reg [4:0] ex_reg_mem_cmd;
  wire[4:0] T534;
  wire[4:0] T535;
  wire[3:0] T536;
  wire[2:0] T537;
  wire[1:0] T538;
  wire T539;
  wire T540;
  wire[31:0] T541;
  wire T542;
  wire T543;
  wire[31:0] T544;
  wire T545;
  wire[31:0] T546;
  wire T547;
  wire T548;
  wire[31:0] T549;
  wire T550;
  wire[31:0] T551;
  wire T552;
  wire T553;
  wire[31:0] T554;
  wire T555;
  wire T556;
  wire[31:0] T557;
  wire T558;
  wire[31:0] T559;
  wire T560;
  wire T561;
  reg [1:0] mem_reg_csr;
  wire[1:0] T562;
  reg [1:0] ex_reg_csr;
  wire[1:0] T563;
  wire data_hazard_mem;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire id_ex_hazard;
  wire T572;
  wire T573;
  wire fp_data_hazard_ex;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire data_hazard_ex;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  reg  ex_reg_load_use;
  wire T603;
  wire id_load_use;
  wire T604;
  wire T605;
  wire replay_ex_structural;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  reg  mem_reg_sret;
  wire T611;
  reg  ex_reg_sret;
  wire T612;
  wire T613;
  wire wb_rocc_val;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  reg  wb_reg_flush_inst;
  wire T618;
  reg  mem_reg_flush_inst;
  wire T619;
  reg  ex_reg_flush_inst;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  reg [1:0] mem_reg_btb_resp_bht_value;
  wire[1:0] T627;
  reg [1:0] ex_reg_btb_resp_bht_value;
  wire[1:0] T628;
  wire T629;
  wire T630;
  reg  ex_reg_btb_hit;
  wire T631;
  reg [3:0] mem_reg_btb_resp_bht_index;
  wire[3:0] T632;
  reg [3:0] ex_reg_btb_resp_bht_index;
  wire[3:0] T633;
  reg [2:0] mem_reg_btb_resp_entry;
  wire[2:0] T634;
  reg [2:0] ex_reg_btb_resp_entry;
  wire[2:0] T635;
  reg [42:0] mem_reg_btb_resp_target;
  wire[42:0] T636;
  reg [42:0] ex_reg_btb_resp_target;
  wire[42:0] T637;
  reg  mem_reg_btb_resp_taken;
  wire T638;
  reg  ex_reg_btb_resp_taken;
  wire T639;
  reg  mem_reg_btb_hit;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  reg [63:0] wb_reg_cause;
  wire[63:0] T645;
  wire[63:0] mem_cause;
  wire[63:0] T646;
  wire[3:0] T647;
  wire[3:0] T648;
  wire[3:0] T649;
  reg [63:0] mem_reg_cause;
  wire[63:0] T650;
  wire[63:0] ex_cause;
  reg [63:0] ex_reg_cause;
  wire[63:0] T651;
  wire[63:0] id_cause;
  wire[63:0] T652;
  wire[3:0] T653;
  wire[3:0] T654;
  wire[3:0] T655;
  wire[3:0] T656;
  wire[3:0] T657;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[63:0] id_interrupt_cause;
  wire[63:0] T660;
  wire[63:0] T661;
  wire[63:0] T662;
  wire[63:0] T663;
  wire[63:0] T664;
  wire[63:0] T665;
  wire T666;
  wire T667;
  reg  wb_reg_valid;
  wire T668;
  wire T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire[1:0] T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire[1:0] T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire[2:0] T711;
  reg [1:0] wb_reg_csr;
  wire[1:0] T712;
  wire T713;
  wire[3:0] T714;
  wire[3:0] T715;
  wire[2:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire[31:0] T720;
  wire T721;
  wire T722;
  wire[31:0] T723;
  wire T724;
  wire[31:0] T725;
  wire T726;
  wire T727;
  wire[31:0] T728;
  wire T729;
  wire T730;
  wire[31:0] T731;
  wire T732;
  wire T733;
  wire[31:0] T734;
  wire T735;
  wire T736;
  wire[31:0] T737;
  wire T738;
  wire[31:0] T739;
  wire T740;
  wire T741;
  wire[31:0] T742;
  wire T743;
  wire T744;
  wire[31:0] T745;
  wire T746;
  wire T747;
  wire[31:0] T748;
  wire T749;
  wire[31:0] T750;
  wire T751;
  wire T752;
  wire[31:0] T753;
  wire T754;
  wire T755;
  wire T756;
  wire[31:0] T757;
  wire T758;
  wire[31:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire[31:0] T763;
  wire T764;
  wire[31:0] T765;
  wire[2:0] T766;
  wire[2:0] T767;
  wire[1:0] T768;
  wire T769;
  wire T770;
  wire[31:0] T771;
  wire T772;
  wire[31:0] T773;
  wire T774;
  wire T775;
  wire[31:0] T776;
  wire T777;
  wire T778;
  wire[31:0] T779;
  wire T780;
  wire T781;
  wire[31:0] T782;
  wire T783;
  wire[31:0] T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire T787;
  wire T788;
  wire[31:0] T789;
  wire T790;
  wire T791;
  wire[31:0] T792;
  wire T793;
  wire T794;
  wire T795;
  wire[31:0] T796;
  wire T797;
  wire[31:0] T798;
  wire T799;
  wire T800;
  wire[31:0] T801;
  wire T802;
  wire[31:0] T803;
  wire[2:0] T804;
  wire[1:0] T805;
  wire[1:0] T806;
  wire T807;
  wire T808;
  wire[31:0] T809;
  wire T810;
  wire T811;
  wire T812;
  wire[31:0] T813;
  wire T814;
  wire T815;
  wire[31:0] T816;
  wire T817;
  wire[31:0] T818;
  wire T819;
  wire T820;
  wire[31:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[31:0] T825;
  wire T826;
  wire T827;
  wire T828;
  wire[2:0] T829;
  wire[1:0] T830;
  wire[1:0] T831;
  wire[1:0] T832;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_xcpt = {1{$random}};
    wb_reg_sret = {1{$random}};
    mem_reg_replay = {1{$random}};
    mem_reg_replay_next = {1{$random}};
    ex_reg_replay_next = {1{$random}};
    id_reg_fence = {1{$random}};
    ex_reg_mem_val = {1{$random}};
    R118 = {1{$random}};
    wb_reg_rocc_val = {1{$random}};
    mem_reg_rocc_val = {1{$random}};
    ex_reg_rocc_val = {1{$random}};
    mem_reg_jal = {1{$random}};
    ex_reg_jal = {1{$random}};
    mem_reg_jalr = {1{$random}};
    ex_reg_jalr = {1{$random}};
    mem_reg_branch = {1{$random}};
    ex_reg_branch = {1{$random}};
    mem_reg_fp_val = {1{$random}};
    ex_reg_fp_val = {1{$random}};
    mem_reg_mem_val = {1{$random}};
    mem_reg_xcpt = {1{$random}};
    ex_reg_xcpt = {1{$random}};
    ex_reg_xcpt_interrupt = {1{$random}};
    mem_reg_xcpt_interrupt = {1{$random}};
    mem_reg_valid = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_reg_wen = {1{$random}};
    ex_reg_wen = {1{$random}};
    wb_reg_replay = {1{$random}};
    wb_reg_fp_wen = {1{$random}};
    mem_reg_fp_wen = {1{$random}};
    ex_reg_fp_wen = {1{$random}};
    wb_reg_mem_val = {1{$random}};
    R409 = {1{$random}};
    wb_reg_div_mul_val = {1{$random}};
    mem_reg_div_mul_val = {1{$random}};
    ex_reg_div_mul_val = {1{$random}};
    wb_reg_fp_val = {1{$random}};
    wb_reg_wen = {1{$random}};
    mem_reg_slow_bypass = {1{$random}};
    ex_reg_mem_type = {1{$random}};
    ex_reg_mem_cmd = {1{$random}};
    mem_reg_csr = {1{$random}};
    ex_reg_csr = {1{$random}};
    ex_reg_load_use = {1{$random}};
    mem_reg_sret = {1{$random}};
    ex_reg_sret = {1{$random}};
    wb_reg_flush_inst = {1{$random}};
    mem_reg_flush_inst = {1{$random}};
    ex_reg_flush_inst = {1{$random}};
    mem_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_resp_bht_value = {1{$random}};
    ex_reg_btb_hit = {1{$random}};
    mem_reg_btb_resp_bht_index = {1{$random}};
    ex_reg_btb_resp_bht_index = {1{$random}};
    mem_reg_btb_resp_entry = {1{$random}};
    ex_reg_btb_resp_entry = {1{$random}};
    mem_reg_btb_resp_target = {2{$random}};
    ex_reg_btb_resp_target = {2{$random}};
    mem_reg_btb_resp_taken = {1{$random}};
    ex_reg_btb_resp_taken = {1{$random}};
    mem_reg_btb_hit = {1{$random}};
    wb_reg_cause = {2{$random}};
    mem_reg_cause = {2{$random}};
    ex_reg_cause = {2{$random}};
    wb_reg_valid = {1{$random}};
    wb_reg_csr = {1{$random}};
  end
`endif

  assign io_rocc_exception = T0;
  assign T0 = wb_reg_xcpt & io_dpath_status_er;
  assign T1 = mem_xcpt & T2;
  assign T2 = take_pc_wb ^ 1'h1;
  assign take_pc_wb = T3;
  assign T3 = T613 | wb_reg_sret;
  assign T4 = ctrl_killm ? 1'h0 : T5;
  assign T5 = mem_reg_sret & T6;
  assign T6 = mem_reg_replay ^ 1'h1;
  assign T7 = T610 & replay_ex;
  assign replay_ex = replay_ex_structural | replay_ex_other;
  assign replay_ex_other = T602 | mem_reg_replay_next;
  assign T8 = ctrl_killx ? 1'h0 : ex_reg_replay_next;
  assign T9 = ctrl_killd ? 1'h0 : T10;
  assign T10 = T31 | id_csr_flush;
  assign id_csr_flush = T18 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T16 | T13;
  assign T13 = T14 == 12'h400;
  assign T14 = T15 & 12'hc0d;
  assign T15 = io_dpath_inst[5'h1f:5'h14];
  assign T16 = T17 == 12'h400;
  assign T17 = T15 & 12'hc0e;
  assign T18 = T30 & id_csr_wen;
  assign id_csr_wen = T28 | T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T27 | T21;
  assign T21 = 2'h3 == T22;
  assign T22 = {T25, T23};
  assign T23 = T24 == 32'h1070;
  assign T24 = io_dpath_inst & 32'h1070;
  assign T25 = T26 == 32'h2070;
  assign T26 = io_dpath_inst & 32'h2070;
  assign T27 = 2'h2 == T22;
  assign T28 = T29 != 5'h0;
  assign T29 = io_dpath_inst[5'h13:4'hf];
  assign T30 = T22 != 2'h0;
  assign T31 = T32 == 32'h1008;
  assign T32 = io_dpath_inst & 32'h3058;
  assign ctrl_killd = T33;
  assign T33 = T64 | ctrl_draind;
  assign ctrl_draind = id_interrupt | ex_reg_replay_next;
  assign id_interrupt = io_dpath_status_ei & id_interrupt_unmasked;
  assign id_interrupt_unmasked = T37 | T34;
  assign T34 = T36 & T35;
  assign T35 = io_dpath_status_ip[3'h7:3'h7];
  assign T36 = io_dpath_status_im[3'h7:3'h7];
  assign T37 = T41 | T38;
  assign T38 = T40 & T39;
  assign T39 = io_dpath_status_ip[3'h6:3'h6];
  assign T40 = io_dpath_status_im[3'h6:3'h6];
  assign T41 = T45 | T42;
  assign T42 = T44 & T43;
  assign T43 = io_dpath_status_ip[3'h5:3'h5];
  assign T44 = io_dpath_status_im[3'h5:3'h5];
  assign T45 = T49 | T46;
  assign T46 = T48 & T47;
  assign T47 = io_dpath_status_ip[3'h4:3'h4];
  assign T48 = io_dpath_status_im[3'h4:3'h4];
  assign T49 = T53 | T50;
  assign T50 = T52 & T51;
  assign T51 = io_dpath_status_ip[2'h3:2'h3];
  assign T52 = io_dpath_status_im[2'h3:2'h3];
  assign T53 = T57 | T54;
  assign T54 = T56 & T55;
  assign T55 = io_dpath_status_ip[2'h2:2'h2];
  assign T56 = io_dpath_status_im[2'h2:2'h2];
  assign T57 = T61 | T58;
  assign T58 = T60 & T59;
  assign T59 = io_dpath_status_ip[1'h1:1'h1];
  assign T60 = io_dpath_status_im[1'h1:1'h1];
  assign T61 = T63 & T62;
  assign T62 = io_dpath_status_ip[1'h0:1'h0];
  assign T63 = io_dpath_status_im[1'h0:1'h0];
  assign T64 = T600 | ctrl_stalld;
  assign ctrl_stalld = T105 | id_do_fence;
  assign id_do_fence = id_mem_busy & T65;
  assign T65 = T66 | id_csr_flush;
  assign T66 = T100 | T67;
  assign T67 = id_reg_fence & T68;
  assign T68 = T71 | T69;
  assign T69 = T70 == 32'h1000202f;
  assign T70 = io_dpath_inst & 32'hf9f0607f;
  assign T71 = T74 | T72;
  assign T72 = T73 == 32'h800202f;
  assign T73 = io_dpath_inst & 32'he800607f;
  assign T74 = T77 | T75;
  assign T75 = T76 == 32'h202f;
  assign T76 = io_dpath_inst & 32'h1800607f;
  assign T77 = T80 | T78;
  assign T78 = T79 == 32'h2003;
  assign T79 = io_dpath_inst & 32'h605b;
  assign T80 = T83 | T81;
  assign T81 = T82 == 32'h3;
  assign T82 = io_dpath_inst & 32'h107f;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h3;
  assign T85 = io_dpath_inst & 32'h207f;
  assign T86 = T87 == 32'h3;
  assign T87 = io_dpath_inst & 32'h405f;
  assign T88 = reset ? 1'h0 : T89;
  assign T89 = id_fence_next | T90;
  assign T90 = id_reg_fence & id_mem_busy;
  assign id_mem_busy = T93 | ex_reg_mem_val;
  assign T91 = ctrl_killd ? 1'h0 : T92;
  assign T92 = T68;
  assign T93 = io_dmem_ordered ^ 1'h1;
  assign id_fence_next = T98 | T94;
  assign T94 = T96 & T95;
  assign T95 = io_dpath_inst[5'h19:5'h19];
  assign T96 = T97 == 32'h2008;
  assign T97 = io_dpath_inst & 32'h6048;
  assign T98 = T99 == 32'h8;
  assign T99 = io_dpath_inst & 32'h3058;
  assign T100 = T103 | T101;
  assign T101 = T102 == 32'h100f;
  assign T102 = io_dpath_inst & 32'h707f;
  assign T103 = T96 & T104;
  assign T104 = io_dpath_inst[5'h1a:5'h1a];
  assign T105 = T108 | T106;
  assign T106 = T68 & T107;
  assign T107 = io_dmem_req_ready ^ 1'h1;
  assign T108 = T397 | T109;
  assign T109 = T152 & id_stall_fpu;
  assign id_stall_fpu = T369 | T110;
  assign T110 = io_fpu_dec_wen & T111;
  assign T111 = T117 & T112;
  assign T112 = T113 - 1'h1;
  assign T113 = 1'h1 << T114;
  assign T114 = T115 + 5'h1;
  assign T115 = T116 - T116;
  assign T116 = io_dpath_inst[4'hb:3'h7];
  assign T117 = R118 >> T116;
  assign T119 = reset ? 32'h0 : T120;
  assign T120 = T368 ? T364 : T121;
  assign T121 = T363 ? T359 : T122;
  assign T122 = T126 ? T123 : R118;
  assign T123 = R118 | T124;
  assign T124 = T126 ? T125 : 32'h0;
  assign T125 = 1'h1 << io_dpath_wb_waddr;
  assign T126 = T351 & T127;
  assign T127 = replay_wb ^ 1'h1;
  assign replay_wb = replay_wb_common | T128;
  assign T128 = wb_reg_rocc_val & T129;
  assign T129 = io_rocc_cmd_ready ^ 1'h1;
  assign T130 = ctrl_killm ? 1'h0 : mem_reg_rocc_val;
  assign T131 = ctrl_killx ? 1'h0 : ex_reg_rocc_val;
  assign T132 = ctrl_killd ? 1'h0 : T133;
  assign T133 = 1'h0;
  assign ctrl_killx = T134;
  assign T134 = take_pc_mem_wb | replay_ex;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign take_pc_mem = io_dpath_mem_misprediction & T135;
  assign T135 = T140 | mem_reg_jal;
  assign T136 = ctrl_killx ? 1'h0 : ex_reg_jal;
  assign T137 = ctrl_killd ? 1'h0 : T138;
  assign T138 = T139 == 32'h68;
  assign T139 = io_dpath_inst & 32'h68;
  assign T140 = mem_reg_branch | mem_reg_jalr;
  assign T141 = ctrl_killx ? 1'h0 : ex_reg_jalr;
  assign T142 = ctrl_killd ? 1'h0 : T143;
  assign T143 = T144 == 32'h24;
  assign T144 = io_dpath_inst & 32'h203c;
  assign T145 = ctrl_killx ? 1'h0 : ex_reg_branch;
  assign T146 = ctrl_killd ? 1'h0 : T147;
  assign T147 = T148 == 32'h60;
  assign T148 = io_dpath_inst & 32'h74;
  assign ctrl_killm = T149;
  assign T149 = T157 | fpu_kill_mem;
  assign fpu_kill_mem = mem_reg_fp_val & io_fpu_nack_mem;
  assign T150 = ctrl_killx ? 1'h0 : ex_reg_fp_val;
  assign T151 = ctrl_killd ? 1'h0 : T152;
  assign T152 = T155 | T153;
  assign T153 = T154 == 32'h40;
  assign T154 = io_dpath_inst & 32'h60;
  assign T155 = T156 == 32'h4;
  assign T156 = io_dpath_inst & 32'h5c;
  assign T157 = killm_common | mem_xcpt;
  assign mem_xcpt = T160 | T158;
  assign T158 = mem_reg_mem_val & io_dmem_xcpt_pf_st;
  assign T159 = ctrl_killx ? 1'h0 : ex_reg_mem_val;
  assign T160 = T162 | T161;
  assign T161 = mem_reg_mem_val & io_dmem_xcpt_pf_ld;
  assign T162 = T164 | T163;
  assign T163 = mem_reg_mem_val & io_dmem_xcpt_ma_st;
  assign T164 = T166 | T165;
  assign T165 = mem_reg_mem_val & io_dmem_xcpt_ma_ld;
  assign T166 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T167 = ctrl_killx ? 1'h0 : ex_xcpt;
  assign ex_xcpt = T169 | T168;
  assign T168 = ex_reg_fp_val & io_fpu_illegal_rm;
  assign T169 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T170 = ctrl_killd ? 1'h0 : id_xcpt;
  assign id_xcpt = T173 | T171;
  assign T171 = T172 == 32'h70;
  assign T172 = io_dpath_inst & 32'h80003070;
  assign T173 = T179 | T174;
  assign T174 = T176 & T175;
  assign T175 = io_dpath_status_ef ^ 1'h1;
  assign T176 = T152 | id_csr_fp;
  assign id_csr_fp = T30 & T177;
  assign T177 = T178 == 12'h0;
  assign T178 = T15 & 12'h480;
  assign T179 = T184 | T180;
  assign T180 = T182 & T181;
  assign T181 = io_dpath_status_s ^ 1'h1;
  assign T182 = T183 == 32'h80000050;
  assign T183 = io_dpath_inst & 32'he0003050;
  assign T184 = T205 | id_csr_privileged;
  assign id_csr_privileged = T30 & T185;
  assign T185 = T191 | T186;
  assign T186 = T187 & id_csr_wen;
  assign T187 = T189 & T188;
  assign T188 = io_dpath_status_s ^ 1'h1;
  assign T189 = T190 == 2'h1;
  assign T190 = T15[4'h9:4'h8];
  assign T191 = T194 | T192;
  assign T192 = 2'h2 <= T193;
  assign T193 = T15[4'h9:4'h8];
  assign T194 = T199 | T195;
  assign T195 = T197 & T196;
  assign T196 = io_dpath_status_s ^ 1'h1;
  assign T197 = T198 == 2'h1;
  assign T198 = T15[4'hb:4'ha];
  assign T199 = T202 | T200;
  assign T200 = T201 == 2'h2;
  assign T201 = T15[4'hb:4'ha];
  assign T202 = T203 & id_csr_wen;
  assign T203 = T204 == 2'h3;
  assign T204 = T15[4'hb:4'ha];
  assign T205 = T311 | T206;
  assign T206 = T210 | id_csr_invalid;
  assign id_csr_invalid = T30 & T207;
  assign T207 = T208 ^ 1'h1;
  always @(*) case (T15)
    0: T208 = 1'h0;
    1: T208 = 1'h1;
    2: T208 = 1'h1;
    3: T208 = 1'h1;
    4: T208 = 1'h0;
    5: T208 = 1'h0;
    6: T208 = 1'h0;
    7: T208 = 1'h0;
    8: T208 = 1'h0;
    9: T208 = 1'h0;
    10: T208 = 1'h0;
    11: T208 = 1'h0;
    12: T208 = 1'h0;
    13: T208 = 1'h0;
    14: T208 = 1'h0;
    15: T208 = 1'h0;
    16: T208 = 1'h0;
    17: T208 = 1'h0;
    18: T208 = 1'h0;
    19: T208 = 1'h0;
    20: T208 = 1'h0;
    21: T208 = 1'h0;
    22: T208 = 1'h0;
    23: T208 = 1'h0;
    24: T208 = 1'h0;
    25: T208 = 1'h0;
    26: T208 = 1'h0;
    27: T208 = 1'h0;
    28: T208 = 1'h0;
    29: T208 = 1'h0;
    30: T208 = 1'h0;
    31: T208 = 1'h0;
    32: T208 = 1'h0;
    33: T208 = 1'h0;
    34: T208 = 1'h0;
    35: T208 = 1'h0;
    36: T208 = 1'h0;
    37: T208 = 1'h0;
    38: T208 = 1'h0;
    39: T208 = 1'h0;
    40: T208 = 1'h0;
    41: T208 = 1'h0;
    42: T208 = 1'h0;
    43: T208 = 1'h0;
    44: T208 = 1'h0;
    45: T208 = 1'h0;
    46: T208 = 1'h0;
    47: T208 = 1'h0;
    48: T208 = 1'h0;
    49: T208 = 1'h0;
    50: T208 = 1'h0;
    51: T208 = 1'h0;
    52: T208 = 1'h0;
    53: T208 = 1'h0;
    54: T208 = 1'h0;
    55: T208 = 1'h0;
    56: T208 = 1'h0;
    57: T208 = 1'h0;
    58: T208 = 1'h0;
    59: T208 = 1'h0;
    60: T208 = 1'h0;
    61: T208 = 1'h0;
    62: T208 = 1'h0;
    63: T208 = 1'h0;
    64: T208 = 1'h0;
    65: T208 = 1'h0;
    66: T208 = 1'h0;
    67: T208 = 1'h0;
    68: T208 = 1'h0;
    69: T208 = 1'h0;
    70: T208 = 1'h0;
    71: T208 = 1'h0;
    72: T208 = 1'h0;
    73: T208 = 1'h0;
    74: T208 = 1'h0;
    75: T208 = 1'h0;
    76: T208 = 1'h0;
    77: T208 = 1'h0;
    78: T208 = 1'h0;
    79: T208 = 1'h0;
    80: T208 = 1'h0;
    81: T208 = 1'h0;
    82: T208 = 1'h0;
    83: T208 = 1'h0;
    84: T208 = 1'h0;
    85: T208 = 1'h0;
    86: T208 = 1'h0;
    87: T208 = 1'h0;
    88: T208 = 1'h0;
    89: T208 = 1'h0;
    90: T208 = 1'h0;
    91: T208 = 1'h0;
    92: T208 = 1'h0;
    93: T208 = 1'h0;
    94: T208 = 1'h0;
    95: T208 = 1'h0;
    96: T208 = 1'h0;
    97: T208 = 1'h0;
    98: T208 = 1'h0;
    99: T208 = 1'h0;
    100: T208 = 1'h0;
    101: T208 = 1'h0;
    102: T208 = 1'h0;
    103: T208 = 1'h0;
    104: T208 = 1'h0;
    105: T208 = 1'h0;
    106: T208 = 1'h0;
    107: T208 = 1'h0;
    108: T208 = 1'h0;
    109: T208 = 1'h0;
    110: T208 = 1'h0;
    111: T208 = 1'h0;
    112: T208 = 1'h0;
    113: T208 = 1'h0;
    114: T208 = 1'h0;
    115: T208 = 1'h0;
    116: T208 = 1'h0;
    117: T208 = 1'h0;
    118: T208 = 1'h0;
    119: T208 = 1'h0;
    120: T208 = 1'h0;
    121: T208 = 1'h0;
    122: T208 = 1'h0;
    123: T208 = 1'h0;
    124: T208 = 1'h0;
    125: T208 = 1'h0;
    126: T208 = 1'h0;
    127: T208 = 1'h0;
    128: T208 = 1'h0;
    129: T208 = 1'h0;
    130: T208 = 1'h0;
    131: T208 = 1'h0;
    132: T208 = 1'h0;
    133: T208 = 1'h0;
    134: T208 = 1'h0;
    135: T208 = 1'h0;
    136: T208 = 1'h0;
    137: T208 = 1'h0;
    138: T208 = 1'h0;
    139: T208 = 1'h0;
    140: T208 = 1'h0;
    141: T208 = 1'h0;
    142: T208 = 1'h0;
    143: T208 = 1'h0;
    144: T208 = 1'h0;
    145: T208 = 1'h0;
    146: T208 = 1'h0;
    147: T208 = 1'h0;
    148: T208 = 1'h0;
    149: T208 = 1'h0;
    150: T208 = 1'h0;
    151: T208 = 1'h0;
    152: T208 = 1'h0;
    153: T208 = 1'h0;
    154: T208 = 1'h0;
    155: T208 = 1'h0;
    156: T208 = 1'h0;
    157: T208 = 1'h0;
    158: T208 = 1'h0;
    159: T208 = 1'h0;
    160: T208 = 1'h0;
    161: T208 = 1'h0;
    162: T208 = 1'h0;
    163: T208 = 1'h0;
    164: T208 = 1'h0;
    165: T208 = 1'h0;
    166: T208 = 1'h0;
    167: T208 = 1'h0;
    168: T208 = 1'h0;
    169: T208 = 1'h0;
    170: T208 = 1'h0;
    171: T208 = 1'h0;
    172: T208 = 1'h0;
    173: T208 = 1'h0;
    174: T208 = 1'h0;
    175: T208 = 1'h0;
    176: T208 = 1'h0;
    177: T208 = 1'h0;
    178: T208 = 1'h0;
    179: T208 = 1'h0;
    180: T208 = 1'h0;
    181: T208 = 1'h0;
    182: T208 = 1'h0;
    183: T208 = 1'h0;
    184: T208 = 1'h0;
    185: T208 = 1'h0;
    186: T208 = 1'h0;
    187: T208 = 1'h0;
    188: T208 = 1'h0;
    189: T208 = 1'h0;
    190: T208 = 1'h0;
    191: T208 = 1'h0;
    192: T208 = 1'h1;
    193: T208 = 1'h0;
    194: T208 = 1'h0;
    195: T208 = 1'h0;
    196: T208 = 1'h0;
    197: T208 = 1'h0;
    198: T208 = 1'h0;
    199: T208 = 1'h0;
    200: T208 = 1'h0;
    201: T208 = 1'h0;
    202: T208 = 1'h0;
    203: T208 = 1'h0;
    204: T208 = 1'h0;
    205: T208 = 1'h0;
    206: T208 = 1'h0;
    207: T208 = 1'h0;
    208: T208 = 1'h0;
    209: T208 = 1'h0;
    210: T208 = 1'h0;
    211: T208 = 1'h0;
    212: T208 = 1'h0;
    213: T208 = 1'h0;
    214: T208 = 1'h0;
    215: T208 = 1'h0;
    216: T208 = 1'h0;
    217: T208 = 1'h0;
    218: T208 = 1'h0;
    219: T208 = 1'h0;
    220: T208 = 1'h0;
    221: T208 = 1'h0;
    222: T208 = 1'h0;
    223: T208 = 1'h0;
    224: T208 = 1'h0;
    225: T208 = 1'h0;
    226: T208 = 1'h0;
    227: T208 = 1'h0;
    228: T208 = 1'h0;
    229: T208 = 1'h0;
    230: T208 = 1'h0;
    231: T208 = 1'h0;
    232: T208 = 1'h0;
    233: T208 = 1'h0;
    234: T208 = 1'h0;
    235: T208 = 1'h0;
    236: T208 = 1'h0;
    237: T208 = 1'h0;
    238: T208 = 1'h0;
    239: T208 = 1'h0;
    240: T208 = 1'h0;
    241: T208 = 1'h0;
    242: T208 = 1'h0;
    243: T208 = 1'h0;
    244: T208 = 1'h0;
    245: T208 = 1'h0;
    246: T208 = 1'h0;
    247: T208 = 1'h0;
    248: T208 = 1'h0;
    249: T208 = 1'h0;
    250: T208 = 1'h0;
    251: T208 = 1'h0;
    252: T208 = 1'h0;
    253: T208 = 1'h0;
    254: T208 = 1'h0;
    255: T208 = 1'h0;
    256: T208 = 1'h0;
    257: T208 = 1'h0;
    258: T208 = 1'h0;
    259: T208 = 1'h0;
    260: T208 = 1'h0;
    261: T208 = 1'h0;
    262: T208 = 1'h0;
    263: T208 = 1'h0;
    264: T208 = 1'h0;
    265: T208 = 1'h0;
    266: T208 = 1'h0;
    267: T208 = 1'h0;
    268: T208 = 1'h0;
    269: T208 = 1'h0;
    270: T208 = 1'h0;
    271: T208 = 1'h0;
    272: T208 = 1'h0;
    273: T208 = 1'h0;
    274: T208 = 1'h0;
    275: T208 = 1'h0;
    276: T208 = 1'h0;
    277: T208 = 1'h0;
    278: T208 = 1'h0;
    279: T208 = 1'h0;
    280: T208 = 1'h0;
    281: T208 = 1'h0;
    282: T208 = 1'h0;
    283: T208 = 1'h0;
    284: T208 = 1'h0;
    285: T208 = 1'h0;
    286: T208 = 1'h0;
    287: T208 = 1'h0;
    288: T208 = 1'h0;
    289: T208 = 1'h0;
    290: T208 = 1'h0;
    291: T208 = 1'h0;
    292: T208 = 1'h0;
    293: T208 = 1'h0;
    294: T208 = 1'h0;
    295: T208 = 1'h0;
    296: T208 = 1'h0;
    297: T208 = 1'h0;
    298: T208 = 1'h0;
    299: T208 = 1'h0;
    300: T208 = 1'h0;
    301: T208 = 1'h0;
    302: T208 = 1'h0;
    303: T208 = 1'h0;
    304: T208 = 1'h0;
    305: T208 = 1'h0;
    306: T208 = 1'h0;
    307: T208 = 1'h0;
    308: T208 = 1'h0;
    309: T208 = 1'h0;
    310: T208 = 1'h0;
    311: T208 = 1'h0;
    312: T208 = 1'h0;
    313: T208 = 1'h0;
    314: T208 = 1'h0;
    315: T208 = 1'h0;
    316: T208 = 1'h0;
    317: T208 = 1'h0;
    318: T208 = 1'h0;
    319: T208 = 1'h0;
    320: T208 = 1'h0;
    321: T208 = 1'h0;
    322: T208 = 1'h0;
    323: T208 = 1'h0;
    324: T208 = 1'h0;
    325: T208 = 1'h0;
    326: T208 = 1'h0;
    327: T208 = 1'h0;
    328: T208 = 1'h0;
    329: T208 = 1'h0;
    330: T208 = 1'h0;
    331: T208 = 1'h0;
    332: T208 = 1'h0;
    333: T208 = 1'h0;
    334: T208 = 1'h0;
    335: T208 = 1'h0;
    336: T208 = 1'h0;
    337: T208 = 1'h0;
    338: T208 = 1'h0;
    339: T208 = 1'h0;
    340: T208 = 1'h0;
    341: T208 = 1'h0;
    342: T208 = 1'h0;
    343: T208 = 1'h0;
    344: T208 = 1'h0;
    345: T208 = 1'h0;
    346: T208 = 1'h0;
    347: T208 = 1'h0;
    348: T208 = 1'h0;
    349: T208 = 1'h0;
    350: T208 = 1'h0;
    351: T208 = 1'h0;
    352: T208 = 1'h0;
    353: T208 = 1'h0;
    354: T208 = 1'h0;
    355: T208 = 1'h0;
    356: T208 = 1'h0;
    357: T208 = 1'h0;
    358: T208 = 1'h0;
    359: T208 = 1'h0;
    360: T208 = 1'h0;
    361: T208 = 1'h0;
    362: T208 = 1'h0;
    363: T208 = 1'h0;
    364: T208 = 1'h0;
    365: T208 = 1'h0;
    366: T208 = 1'h0;
    367: T208 = 1'h0;
    368: T208 = 1'h0;
    369: T208 = 1'h0;
    370: T208 = 1'h0;
    371: T208 = 1'h0;
    372: T208 = 1'h0;
    373: T208 = 1'h0;
    374: T208 = 1'h0;
    375: T208 = 1'h0;
    376: T208 = 1'h0;
    377: T208 = 1'h0;
    378: T208 = 1'h0;
    379: T208 = 1'h0;
    380: T208 = 1'h0;
    381: T208 = 1'h0;
    382: T208 = 1'h0;
    383: T208 = 1'h0;
    384: T208 = 1'h0;
    385: T208 = 1'h0;
    386: T208 = 1'h0;
    387: T208 = 1'h0;
    388: T208 = 1'h0;
    389: T208 = 1'h0;
    390: T208 = 1'h0;
    391: T208 = 1'h0;
    392: T208 = 1'h0;
    393: T208 = 1'h0;
    394: T208 = 1'h0;
    395: T208 = 1'h0;
    396: T208 = 1'h0;
    397: T208 = 1'h0;
    398: T208 = 1'h0;
    399: T208 = 1'h0;
    400: T208 = 1'h0;
    401: T208 = 1'h0;
    402: T208 = 1'h0;
    403: T208 = 1'h0;
    404: T208 = 1'h0;
    405: T208 = 1'h0;
    406: T208 = 1'h0;
    407: T208 = 1'h0;
    408: T208 = 1'h0;
    409: T208 = 1'h0;
    410: T208 = 1'h0;
    411: T208 = 1'h0;
    412: T208 = 1'h0;
    413: T208 = 1'h0;
    414: T208 = 1'h0;
    415: T208 = 1'h0;
    416: T208 = 1'h0;
    417: T208 = 1'h0;
    418: T208 = 1'h0;
    419: T208 = 1'h0;
    420: T208 = 1'h0;
    421: T208 = 1'h0;
    422: T208 = 1'h0;
    423: T208 = 1'h0;
    424: T208 = 1'h0;
    425: T208 = 1'h0;
    426: T208 = 1'h0;
    427: T208 = 1'h0;
    428: T208 = 1'h0;
    429: T208 = 1'h0;
    430: T208 = 1'h0;
    431: T208 = 1'h0;
    432: T208 = 1'h0;
    433: T208 = 1'h0;
    434: T208 = 1'h0;
    435: T208 = 1'h0;
    436: T208 = 1'h0;
    437: T208 = 1'h0;
    438: T208 = 1'h0;
    439: T208 = 1'h0;
    440: T208 = 1'h0;
    441: T208 = 1'h0;
    442: T208 = 1'h0;
    443: T208 = 1'h0;
    444: T208 = 1'h0;
    445: T208 = 1'h0;
    446: T208 = 1'h0;
    447: T208 = 1'h0;
    448: T208 = 1'h0;
    449: T208 = 1'h0;
    450: T208 = 1'h0;
    451: T208 = 1'h0;
    452: T208 = 1'h0;
    453: T208 = 1'h0;
    454: T208 = 1'h0;
    455: T208 = 1'h0;
    456: T208 = 1'h0;
    457: T208 = 1'h0;
    458: T208 = 1'h0;
    459: T208 = 1'h0;
    460: T208 = 1'h0;
    461: T208 = 1'h0;
    462: T208 = 1'h0;
    463: T208 = 1'h0;
    464: T208 = 1'h0;
    465: T208 = 1'h0;
    466: T208 = 1'h0;
    467: T208 = 1'h0;
    468: T208 = 1'h0;
    469: T208 = 1'h0;
    470: T208 = 1'h0;
    471: T208 = 1'h0;
    472: T208 = 1'h0;
    473: T208 = 1'h0;
    474: T208 = 1'h0;
    475: T208 = 1'h0;
    476: T208 = 1'h0;
    477: T208 = 1'h0;
    478: T208 = 1'h0;
    479: T208 = 1'h0;
    480: T208 = 1'h0;
    481: T208 = 1'h0;
    482: T208 = 1'h0;
    483: T208 = 1'h0;
    484: T208 = 1'h0;
    485: T208 = 1'h0;
    486: T208 = 1'h0;
    487: T208 = 1'h0;
    488: T208 = 1'h0;
    489: T208 = 1'h0;
    490: T208 = 1'h0;
    491: T208 = 1'h0;
    492: T208 = 1'h0;
    493: T208 = 1'h0;
    494: T208 = 1'h0;
    495: T208 = 1'h0;
    496: T208 = 1'h0;
    497: T208 = 1'h0;
    498: T208 = 1'h0;
    499: T208 = 1'h0;
    500: T208 = 1'h0;
    501: T208 = 1'h0;
    502: T208 = 1'h0;
    503: T208 = 1'h0;
    504: T208 = 1'h0;
    505: T208 = 1'h0;
    506: T208 = 1'h0;
    507: T208 = 1'h0;
    508: T208 = 1'h0;
    509: T208 = 1'h0;
    510: T208 = 1'h0;
    511: T208 = 1'h0;
    512: T208 = 1'h0;
    513: T208 = 1'h0;
    514: T208 = 1'h0;
    515: T208 = 1'h0;
    516: T208 = 1'h0;
    517: T208 = 1'h0;
    518: T208 = 1'h0;
    519: T208 = 1'h0;
    520: T208 = 1'h0;
    521: T208 = 1'h0;
    522: T208 = 1'h0;
    523: T208 = 1'h0;
    524: T208 = 1'h0;
    525: T208 = 1'h0;
    526: T208 = 1'h0;
    527: T208 = 1'h0;
    528: T208 = 1'h0;
    529: T208 = 1'h0;
    530: T208 = 1'h0;
    531: T208 = 1'h0;
    532: T208 = 1'h0;
    533: T208 = 1'h0;
    534: T208 = 1'h0;
    535: T208 = 1'h0;
    536: T208 = 1'h0;
    537: T208 = 1'h0;
    538: T208 = 1'h0;
    539: T208 = 1'h0;
    540: T208 = 1'h0;
    541: T208 = 1'h0;
    542: T208 = 1'h0;
    543: T208 = 1'h0;
    544: T208 = 1'h0;
    545: T208 = 1'h0;
    546: T208 = 1'h0;
    547: T208 = 1'h0;
    548: T208 = 1'h0;
    549: T208 = 1'h0;
    550: T208 = 1'h0;
    551: T208 = 1'h0;
    552: T208 = 1'h0;
    553: T208 = 1'h0;
    554: T208 = 1'h0;
    555: T208 = 1'h0;
    556: T208 = 1'h0;
    557: T208 = 1'h0;
    558: T208 = 1'h0;
    559: T208 = 1'h0;
    560: T208 = 1'h0;
    561: T208 = 1'h0;
    562: T208 = 1'h0;
    563: T208 = 1'h0;
    564: T208 = 1'h0;
    565: T208 = 1'h0;
    566: T208 = 1'h0;
    567: T208 = 1'h0;
    568: T208 = 1'h0;
    569: T208 = 1'h0;
    570: T208 = 1'h0;
    571: T208 = 1'h0;
    572: T208 = 1'h0;
    573: T208 = 1'h0;
    574: T208 = 1'h0;
    575: T208 = 1'h0;
    576: T208 = 1'h0;
    577: T208 = 1'h0;
    578: T208 = 1'h0;
    579: T208 = 1'h0;
    580: T208 = 1'h0;
    581: T208 = 1'h0;
    582: T208 = 1'h0;
    583: T208 = 1'h0;
    584: T208 = 1'h0;
    585: T208 = 1'h0;
    586: T208 = 1'h0;
    587: T208 = 1'h0;
    588: T208 = 1'h0;
    589: T208 = 1'h0;
    590: T208 = 1'h0;
    591: T208 = 1'h0;
    592: T208 = 1'h0;
    593: T208 = 1'h0;
    594: T208 = 1'h0;
    595: T208 = 1'h0;
    596: T208 = 1'h0;
    597: T208 = 1'h0;
    598: T208 = 1'h0;
    599: T208 = 1'h0;
    600: T208 = 1'h0;
    601: T208 = 1'h0;
    602: T208 = 1'h0;
    603: T208 = 1'h0;
    604: T208 = 1'h0;
    605: T208 = 1'h0;
    606: T208 = 1'h0;
    607: T208 = 1'h0;
    608: T208 = 1'h0;
    609: T208 = 1'h0;
    610: T208 = 1'h0;
    611: T208 = 1'h0;
    612: T208 = 1'h0;
    613: T208 = 1'h0;
    614: T208 = 1'h0;
    615: T208 = 1'h0;
    616: T208 = 1'h0;
    617: T208 = 1'h0;
    618: T208 = 1'h0;
    619: T208 = 1'h0;
    620: T208 = 1'h0;
    621: T208 = 1'h0;
    622: T208 = 1'h0;
    623: T208 = 1'h0;
    624: T208 = 1'h0;
    625: T208 = 1'h0;
    626: T208 = 1'h0;
    627: T208 = 1'h0;
    628: T208 = 1'h0;
    629: T208 = 1'h0;
    630: T208 = 1'h0;
    631: T208 = 1'h0;
    632: T208 = 1'h0;
    633: T208 = 1'h0;
    634: T208 = 1'h0;
    635: T208 = 1'h0;
    636: T208 = 1'h0;
    637: T208 = 1'h0;
    638: T208 = 1'h0;
    639: T208 = 1'h0;
    640: T208 = 1'h0;
    641: T208 = 1'h0;
    642: T208 = 1'h0;
    643: T208 = 1'h0;
    644: T208 = 1'h0;
    645: T208 = 1'h0;
    646: T208 = 1'h0;
    647: T208 = 1'h0;
    648: T208 = 1'h0;
    649: T208 = 1'h0;
    650: T208 = 1'h0;
    651: T208 = 1'h0;
    652: T208 = 1'h0;
    653: T208 = 1'h0;
    654: T208 = 1'h0;
    655: T208 = 1'h0;
    656: T208 = 1'h0;
    657: T208 = 1'h0;
    658: T208 = 1'h0;
    659: T208 = 1'h0;
    660: T208 = 1'h0;
    661: T208 = 1'h0;
    662: T208 = 1'h0;
    663: T208 = 1'h0;
    664: T208 = 1'h0;
    665: T208 = 1'h0;
    666: T208 = 1'h0;
    667: T208 = 1'h0;
    668: T208 = 1'h0;
    669: T208 = 1'h0;
    670: T208 = 1'h0;
    671: T208 = 1'h0;
    672: T208 = 1'h0;
    673: T208 = 1'h0;
    674: T208 = 1'h0;
    675: T208 = 1'h0;
    676: T208 = 1'h0;
    677: T208 = 1'h0;
    678: T208 = 1'h0;
    679: T208 = 1'h0;
    680: T208 = 1'h0;
    681: T208 = 1'h0;
    682: T208 = 1'h0;
    683: T208 = 1'h0;
    684: T208 = 1'h0;
    685: T208 = 1'h0;
    686: T208 = 1'h0;
    687: T208 = 1'h0;
    688: T208 = 1'h0;
    689: T208 = 1'h0;
    690: T208 = 1'h0;
    691: T208 = 1'h0;
    692: T208 = 1'h0;
    693: T208 = 1'h0;
    694: T208 = 1'h0;
    695: T208 = 1'h0;
    696: T208 = 1'h0;
    697: T208 = 1'h0;
    698: T208 = 1'h0;
    699: T208 = 1'h0;
    700: T208 = 1'h0;
    701: T208 = 1'h0;
    702: T208 = 1'h0;
    703: T208 = 1'h0;
    704: T208 = 1'h0;
    705: T208 = 1'h0;
    706: T208 = 1'h0;
    707: T208 = 1'h0;
    708: T208 = 1'h0;
    709: T208 = 1'h0;
    710: T208 = 1'h0;
    711: T208 = 1'h0;
    712: T208 = 1'h0;
    713: T208 = 1'h0;
    714: T208 = 1'h0;
    715: T208 = 1'h0;
    716: T208 = 1'h0;
    717: T208 = 1'h0;
    718: T208 = 1'h0;
    719: T208 = 1'h0;
    720: T208 = 1'h0;
    721: T208 = 1'h0;
    722: T208 = 1'h0;
    723: T208 = 1'h0;
    724: T208 = 1'h0;
    725: T208 = 1'h0;
    726: T208 = 1'h0;
    727: T208 = 1'h0;
    728: T208 = 1'h0;
    729: T208 = 1'h0;
    730: T208 = 1'h0;
    731: T208 = 1'h0;
    732: T208 = 1'h0;
    733: T208 = 1'h0;
    734: T208 = 1'h0;
    735: T208 = 1'h0;
    736: T208 = 1'h0;
    737: T208 = 1'h0;
    738: T208 = 1'h0;
    739: T208 = 1'h0;
    740: T208 = 1'h0;
    741: T208 = 1'h0;
    742: T208 = 1'h0;
    743: T208 = 1'h0;
    744: T208 = 1'h0;
    745: T208 = 1'h0;
    746: T208 = 1'h0;
    747: T208 = 1'h0;
    748: T208 = 1'h0;
    749: T208 = 1'h0;
    750: T208 = 1'h0;
    751: T208 = 1'h0;
    752: T208 = 1'h0;
    753: T208 = 1'h0;
    754: T208 = 1'h0;
    755: T208 = 1'h0;
    756: T208 = 1'h0;
    757: T208 = 1'h0;
    758: T208 = 1'h0;
    759: T208 = 1'h0;
    760: T208 = 1'h0;
    761: T208 = 1'h0;
    762: T208 = 1'h0;
    763: T208 = 1'h0;
    764: T208 = 1'h0;
    765: T208 = 1'h0;
    766: T208 = 1'h0;
    767: T208 = 1'h0;
    768: T208 = 1'h0;
    769: T208 = 1'h0;
    770: T208 = 1'h0;
    771: T208 = 1'h0;
    772: T208 = 1'h0;
    773: T208 = 1'h0;
    774: T208 = 1'h0;
    775: T208 = 1'h0;
    776: T208 = 1'h0;
    777: T208 = 1'h0;
    778: T208 = 1'h0;
    779: T208 = 1'h0;
    780: T208 = 1'h0;
    781: T208 = 1'h0;
    782: T208 = 1'h0;
    783: T208 = 1'h0;
    784: T208 = 1'h0;
    785: T208 = 1'h0;
    786: T208 = 1'h0;
    787: T208 = 1'h0;
    788: T208 = 1'h0;
    789: T208 = 1'h0;
    790: T208 = 1'h0;
    791: T208 = 1'h0;
    792: T208 = 1'h0;
    793: T208 = 1'h0;
    794: T208 = 1'h0;
    795: T208 = 1'h0;
    796: T208 = 1'h0;
    797: T208 = 1'h0;
    798: T208 = 1'h0;
    799: T208 = 1'h0;
    800: T208 = 1'h0;
    801: T208 = 1'h0;
    802: T208 = 1'h0;
    803: T208 = 1'h0;
    804: T208 = 1'h0;
    805: T208 = 1'h0;
    806: T208 = 1'h0;
    807: T208 = 1'h0;
    808: T208 = 1'h0;
    809: T208 = 1'h0;
    810: T208 = 1'h0;
    811: T208 = 1'h0;
    812: T208 = 1'h0;
    813: T208 = 1'h0;
    814: T208 = 1'h0;
    815: T208 = 1'h0;
    816: T208 = 1'h0;
    817: T208 = 1'h0;
    818: T208 = 1'h0;
    819: T208 = 1'h0;
    820: T208 = 1'h0;
    821: T208 = 1'h0;
    822: T208 = 1'h0;
    823: T208 = 1'h0;
    824: T208 = 1'h0;
    825: T208 = 1'h0;
    826: T208 = 1'h0;
    827: T208 = 1'h0;
    828: T208 = 1'h0;
    829: T208 = 1'h0;
    830: T208 = 1'h0;
    831: T208 = 1'h0;
    832: T208 = 1'h0;
    833: T208 = 1'h0;
    834: T208 = 1'h0;
    835: T208 = 1'h0;
    836: T208 = 1'h0;
    837: T208 = 1'h0;
    838: T208 = 1'h0;
    839: T208 = 1'h0;
    840: T208 = 1'h0;
    841: T208 = 1'h0;
    842: T208 = 1'h0;
    843: T208 = 1'h0;
    844: T208 = 1'h0;
    845: T208 = 1'h0;
    846: T208 = 1'h0;
    847: T208 = 1'h0;
    848: T208 = 1'h0;
    849: T208 = 1'h0;
    850: T208 = 1'h0;
    851: T208 = 1'h0;
    852: T208 = 1'h0;
    853: T208 = 1'h0;
    854: T208 = 1'h0;
    855: T208 = 1'h0;
    856: T208 = 1'h0;
    857: T208 = 1'h0;
    858: T208 = 1'h0;
    859: T208 = 1'h0;
    860: T208 = 1'h0;
    861: T208 = 1'h0;
    862: T208 = 1'h0;
    863: T208 = 1'h0;
    864: T208 = 1'h0;
    865: T208 = 1'h0;
    866: T208 = 1'h0;
    867: T208 = 1'h0;
    868: T208 = 1'h0;
    869: T208 = 1'h0;
    870: T208 = 1'h0;
    871: T208 = 1'h0;
    872: T208 = 1'h0;
    873: T208 = 1'h0;
    874: T208 = 1'h0;
    875: T208 = 1'h0;
    876: T208 = 1'h0;
    877: T208 = 1'h0;
    878: T208 = 1'h0;
    879: T208 = 1'h0;
    880: T208 = 1'h0;
    881: T208 = 1'h0;
    882: T208 = 1'h0;
    883: T208 = 1'h0;
    884: T208 = 1'h0;
    885: T208 = 1'h0;
    886: T208 = 1'h0;
    887: T208 = 1'h0;
    888: T208 = 1'h0;
    889: T208 = 1'h0;
    890: T208 = 1'h0;
    891: T208 = 1'h0;
    892: T208 = 1'h0;
    893: T208 = 1'h0;
    894: T208 = 1'h0;
    895: T208 = 1'h0;
    896: T208 = 1'h0;
    897: T208 = 1'h0;
    898: T208 = 1'h0;
    899: T208 = 1'h0;
    900: T208 = 1'h0;
    901: T208 = 1'h0;
    902: T208 = 1'h0;
    903: T208 = 1'h0;
    904: T208 = 1'h0;
    905: T208 = 1'h0;
    906: T208 = 1'h0;
    907: T208 = 1'h0;
    908: T208 = 1'h0;
    909: T208 = 1'h0;
    910: T208 = 1'h0;
    911: T208 = 1'h0;
    912: T208 = 1'h0;
    913: T208 = 1'h0;
    914: T208 = 1'h0;
    915: T208 = 1'h0;
    916: T208 = 1'h0;
    917: T208 = 1'h0;
    918: T208 = 1'h0;
    919: T208 = 1'h0;
    920: T208 = 1'h0;
    921: T208 = 1'h0;
    922: T208 = 1'h0;
    923: T208 = 1'h0;
    924: T208 = 1'h0;
    925: T208 = 1'h0;
    926: T208 = 1'h0;
    927: T208 = 1'h0;
    928: T208 = 1'h0;
    929: T208 = 1'h0;
    930: T208 = 1'h0;
    931: T208 = 1'h0;
    932: T208 = 1'h0;
    933: T208 = 1'h0;
    934: T208 = 1'h0;
    935: T208 = 1'h0;
    936: T208 = 1'h0;
    937: T208 = 1'h0;
    938: T208 = 1'h0;
    939: T208 = 1'h0;
    940: T208 = 1'h0;
    941: T208 = 1'h0;
    942: T208 = 1'h0;
    943: T208 = 1'h0;
    944: T208 = 1'h0;
    945: T208 = 1'h0;
    946: T208 = 1'h0;
    947: T208 = 1'h0;
    948: T208 = 1'h0;
    949: T208 = 1'h0;
    950: T208 = 1'h0;
    951: T208 = 1'h0;
    952: T208 = 1'h0;
    953: T208 = 1'h0;
    954: T208 = 1'h0;
    955: T208 = 1'h0;
    956: T208 = 1'h0;
    957: T208 = 1'h0;
    958: T208 = 1'h0;
    959: T208 = 1'h0;
    960: T208 = 1'h0;
    961: T208 = 1'h0;
    962: T208 = 1'h0;
    963: T208 = 1'h0;
    964: T208 = 1'h0;
    965: T208 = 1'h0;
    966: T208 = 1'h0;
    967: T208 = 1'h0;
    968: T208 = 1'h0;
    969: T208 = 1'h0;
    970: T208 = 1'h0;
    971: T208 = 1'h0;
    972: T208 = 1'h0;
    973: T208 = 1'h0;
    974: T208 = 1'h0;
    975: T208 = 1'h0;
    976: T208 = 1'h0;
    977: T208 = 1'h0;
    978: T208 = 1'h0;
    979: T208 = 1'h0;
    980: T208 = 1'h0;
    981: T208 = 1'h0;
    982: T208 = 1'h0;
    983: T208 = 1'h0;
    984: T208 = 1'h0;
    985: T208 = 1'h0;
    986: T208 = 1'h0;
    987: T208 = 1'h0;
    988: T208 = 1'h0;
    989: T208 = 1'h0;
    990: T208 = 1'h0;
    991: T208 = 1'h0;
    992: T208 = 1'h0;
    993: T208 = 1'h0;
    994: T208 = 1'h0;
    995: T208 = 1'h0;
    996: T208 = 1'h0;
    997: T208 = 1'h0;
    998: T208 = 1'h0;
    999: T208 = 1'h0;
    1000: T208 = 1'h0;
    1001: T208 = 1'h0;
    1002: T208 = 1'h0;
    1003: T208 = 1'h0;
    1004: T208 = 1'h0;
    1005: T208 = 1'h0;
    1006: T208 = 1'h0;
    1007: T208 = 1'h0;
    1008: T208 = 1'h0;
    1009: T208 = 1'h0;
    1010: T208 = 1'h0;
    1011: T208 = 1'h0;
    1012: T208 = 1'h0;
    1013: T208 = 1'h0;
    1014: T208 = 1'h0;
    1015: T208 = 1'h0;
    1016: T208 = 1'h0;
    1017: T208 = 1'h0;
    1018: T208 = 1'h0;
    1019: T208 = 1'h0;
    1020: T208 = 1'h0;
    1021: T208 = 1'h0;
    1022: T208 = 1'h0;
    1023: T208 = 1'h0;
    1024: T208 = 1'h0;
    1025: T208 = 1'h0;
    1026: T208 = 1'h0;
    1027: T208 = 1'h0;
    1028: T208 = 1'h0;
    1029: T208 = 1'h0;
    1030: T208 = 1'h0;
    1031: T208 = 1'h0;
    1032: T208 = 1'h0;
    1033: T208 = 1'h0;
    1034: T208 = 1'h0;
    1035: T208 = 1'h0;
    1036: T208 = 1'h0;
    1037: T208 = 1'h0;
    1038: T208 = 1'h0;
    1039: T208 = 1'h0;
    1040: T208 = 1'h0;
    1041: T208 = 1'h0;
    1042: T208 = 1'h0;
    1043: T208 = 1'h0;
    1044: T208 = 1'h0;
    1045: T208 = 1'h0;
    1046: T208 = 1'h0;
    1047: T208 = 1'h0;
    1048: T208 = 1'h0;
    1049: T208 = 1'h0;
    1050: T208 = 1'h0;
    1051: T208 = 1'h0;
    1052: T208 = 1'h0;
    1053: T208 = 1'h0;
    1054: T208 = 1'h0;
    1055: T208 = 1'h0;
    1056: T208 = 1'h0;
    1057: T208 = 1'h0;
    1058: T208 = 1'h0;
    1059: T208 = 1'h0;
    1060: T208 = 1'h0;
    1061: T208 = 1'h0;
    1062: T208 = 1'h0;
    1063: T208 = 1'h0;
    1064: T208 = 1'h0;
    1065: T208 = 1'h0;
    1066: T208 = 1'h0;
    1067: T208 = 1'h0;
    1068: T208 = 1'h0;
    1069: T208 = 1'h0;
    1070: T208 = 1'h0;
    1071: T208 = 1'h0;
    1072: T208 = 1'h0;
    1073: T208 = 1'h0;
    1074: T208 = 1'h0;
    1075: T208 = 1'h0;
    1076: T208 = 1'h0;
    1077: T208 = 1'h0;
    1078: T208 = 1'h0;
    1079: T208 = 1'h0;
    1080: T208 = 1'h0;
    1081: T208 = 1'h0;
    1082: T208 = 1'h0;
    1083: T208 = 1'h0;
    1084: T208 = 1'h0;
    1085: T208 = 1'h0;
    1086: T208 = 1'h0;
    1087: T208 = 1'h0;
    1088: T208 = 1'h0;
    1089: T208 = 1'h0;
    1090: T208 = 1'h0;
    1091: T208 = 1'h0;
    1092: T208 = 1'h0;
    1093: T208 = 1'h0;
    1094: T208 = 1'h0;
    1095: T208 = 1'h0;
    1096: T208 = 1'h0;
    1097: T208 = 1'h0;
    1098: T208 = 1'h0;
    1099: T208 = 1'h0;
    1100: T208 = 1'h0;
    1101: T208 = 1'h0;
    1102: T208 = 1'h0;
    1103: T208 = 1'h0;
    1104: T208 = 1'h0;
    1105: T208 = 1'h0;
    1106: T208 = 1'h0;
    1107: T208 = 1'h0;
    1108: T208 = 1'h0;
    1109: T208 = 1'h0;
    1110: T208 = 1'h0;
    1111: T208 = 1'h0;
    1112: T208 = 1'h0;
    1113: T208 = 1'h0;
    1114: T208 = 1'h0;
    1115: T208 = 1'h0;
    1116: T208 = 1'h0;
    1117: T208 = 1'h0;
    1118: T208 = 1'h0;
    1119: T208 = 1'h0;
    1120: T208 = 1'h0;
    1121: T208 = 1'h0;
    1122: T208 = 1'h0;
    1123: T208 = 1'h0;
    1124: T208 = 1'h0;
    1125: T208 = 1'h0;
    1126: T208 = 1'h0;
    1127: T208 = 1'h0;
    1128: T208 = 1'h0;
    1129: T208 = 1'h0;
    1130: T208 = 1'h0;
    1131: T208 = 1'h0;
    1132: T208 = 1'h0;
    1133: T208 = 1'h0;
    1134: T208 = 1'h0;
    1135: T208 = 1'h0;
    1136: T208 = 1'h0;
    1137: T208 = 1'h0;
    1138: T208 = 1'h0;
    1139: T208 = 1'h0;
    1140: T208 = 1'h0;
    1141: T208 = 1'h0;
    1142: T208 = 1'h0;
    1143: T208 = 1'h0;
    1144: T208 = 1'h0;
    1145: T208 = 1'h0;
    1146: T208 = 1'h0;
    1147: T208 = 1'h0;
    1148: T208 = 1'h0;
    1149: T208 = 1'h0;
    1150: T208 = 1'h0;
    1151: T208 = 1'h0;
    1152: T208 = 1'h0;
    1153: T208 = 1'h0;
    1154: T208 = 1'h0;
    1155: T208 = 1'h0;
    1156: T208 = 1'h0;
    1157: T208 = 1'h0;
    1158: T208 = 1'h0;
    1159: T208 = 1'h0;
    1160: T208 = 1'h0;
    1161: T208 = 1'h0;
    1162: T208 = 1'h0;
    1163: T208 = 1'h0;
    1164: T208 = 1'h0;
    1165: T208 = 1'h0;
    1166: T208 = 1'h0;
    1167: T208 = 1'h0;
    1168: T208 = 1'h0;
    1169: T208 = 1'h0;
    1170: T208 = 1'h0;
    1171: T208 = 1'h0;
    1172: T208 = 1'h0;
    1173: T208 = 1'h0;
    1174: T208 = 1'h0;
    1175: T208 = 1'h0;
    1176: T208 = 1'h0;
    1177: T208 = 1'h0;
    1178: T208 = 1'h0;
    1179: T208 = 1'h0;
    1180: T208 = 1'h0;
    1181: T208 = 1'h0;
    1182: T208 = 1'h0;
    1183: T208 = 1'h0;
    1184: T208 = 1'h0;
    1185: T208 = 1'h0;
    1186: T208 = 1'h0;
    1187: T208 = 1'h0;
    1188: T208 = 1'h0;
    1189: T208 = 1'h0;
    1190: T208 = 1'h0;
    1191: T208 = 1'h0;
    1192: T208 = 1'h0;
    1193: T208 = 1'h0;
    1194: T208 = 1'h0;
    1195: T208 = 1'h0;
    1196: T208 = 1'h0;
    1197: T208 = 1'h0;
    1198: T208 = 1'h0;
    1199: T208 = 1'h0;
    1200: T208 = 1'h0;
    1201: T208 = 1'h0;
    1202: T208 = 1'h0;
    1203: T208 = 1'h0;
    1204: T208 = 1'h0;
    1205: T208 = 1'h0;
    1206: T208 = 1'h0;
    1207: T208 = 1'h0;
    1208: T208 = 1'h0;
    1209: T208 = 1'h0;
    1210: T208 = 1'h0;
    1211: T208 = 1'h0;
    1212: T208 = 1'h0;
    1213: T208 = 1'h0;
    1214: T208 = 1'h0;
    1215: T208 = 1'h0;
    1216: T208 = 1'h0;
    1217: T208 = 1'h0;
    1218: T208 = 1'h0;
    1219: T208 = 1'h0;
    1220: T208 = 1'h0;
    1221: T208 = 1'h0;
    1222: T208 = 1'h0;
    1223: T208 = 1'h0;
    1224: T208 = 1'h0;
    1225: T208 = 1'h0;
    1226: T208 = 1'h0;
    1227: T208 = 1'h0;
    1228: T208 = 1'h0;
    1229: T208 = 1'h0;
    1230: T208 = 1'h0;
    1231: T208 = 1'h0;
    1232: T208 = 1'h0;
    1233: T208 = 1'h0;
    1234: T208 = 1'h0;
    1235: T208 = 1'h0;
    1236: T208 = 1'h0;
    1237: T208 = 1'h0;
    1238: T208 = 1'h0;
    1239: T208 = 1'h0;
    1240: T208 = 1'h0;
    1241: T208 = 1'h0;
    1242: T208 = 1'h0;
    1243: T208 = 1'h0;
    1244: T208 = 1'h0;
    1245: T208 = 1'h0;
    1246: T208 = 1'h0;
    1247: T208 = 1'h0;
    1248: T208 = 1'h0;
    1249: T208 = 1'h0;
    1250: T208 = 1'h0;
    1251: T208 = 1'h0;
    1252: T208 = 1'h0;
    1253: T208 = 1'h0;
    1254: T208 = 1'h0;
    1255: T208 = 1'h0;
    1256: T208 = 1'h0;
    1257: T208 = 1'h0;
    1258: T208 = 1'h0;
    1259: T208 = 1'h0;
    1260: T208 = 1'h0;
    1261: T208 = 1'h0;
    1262: T208 = 1'h0;
    1263: T208 = 1'h0;
    1264: T208 = 1'h0;
    1265: T208 = 1'h0;
    1266: T208 = 1'h0;
    1267: T208 = 1'h0;
    1268: T208 = 1'h0;
    1269: T208 = 1'h0;
    1270: T208 = 1'h0;
    1271: T208 = 1'h0;
    1272: T208 = 1'h0;
    1273: T208 = 1'h0;
    1274: T208 = 1'h0;
    1275: T208 = 1'h0;
    1276: T208 = 1'h0;
    1277: T208 = 1'h0;
    1278: T208 = 1'h0;
    1279: T208 = 1'h0;
    1280: T208 = 1'h1;
    1281: T208 = 1'h1;
    1282: T208 = 1'h1;
    1283: T208 = 1'h1;
    1284: T208 = 1'h1;
    1285: T208 = 1'h1;
    1286: T208 = 1'h1;
    1287: T208 = 1'h1;
    1288: T208 = 1'h1;
    1289: T208 = 1'h1;
    1290: T208 = 1'h1;
    1291: T208 = 1'h1;
    1292: T208 = 1'h1;
    1293: T208 = 1'h1;
    1294: T208 = 1'h1;
    1295: T208 = 1'h1;
    1296: T208 = 1'h0;
    1297: T208 = 1'h0;
    1298: T208 = 1'h0;
    1299: T208 = 1'h0;
    1300: T208 = 1'h0;
    1301: T208 = 1'h0;
    1302: T208 = 1'h0;
    1303: T208 = 1'h0;
    1304: T208 = 1'h0;
    1305: T208 = 1'h0;
    1306: T208 = 1'h0;
    1307: T208 = 1'h0;
    1308: T208 = 1'h0;
    1309: T208 = 1'h1;
    1310: T208 = 1'h1;
    1311: T208 = 1'h1;
    1312: T208 = 1'h0;
    1313: T208 = 1'h0;
    1314: T208 = 1'h0;
    1315: T208 = 1'h0;
    1316: T208 = 1'h0;
    1317: T208 = 1'h0;
    1318: T208 = 1'h0;
    1319: T208 = 1'h0;
    1320: T208 = 1'h0;
    1321: T208 = 1'h0;
    1322: T208 = 1'h0;
    1323: T208 = 1'h0;
    1324: T208 = 1'h0;
    1325: T208 = 1'h0;
    1326: T208 = 1'h0;
    1327: T208 = 1'h0;
    1328: T208 = 1'h0;
    1329: T208 = 1'h0;
    1330: T208 = 1'h0;
    1331: T208 = 1'h0;
    1332: T208 = 1'h0;
    1333: T208 = 1'h0;
    1334: T208 = 1'h0;
    1335: T208 = 1'h0;
    1336: T208 = 1'h0;
    1337: T208 = 1'h0;
    1338: T208 = 1'h0;
    1339: T208 = 1'h0;
    1340: T208 = 1'h0;
    1341: T208 = 1'h0;
    1342: T208 = 1'h0;
    1343: T208 = 1'h0;
    1344: T208 = 1'h0;
    1345: T208 = 1'h0;
    1346: T208 = 1'h0;
    1347: T208 = 1'h0;
    1348: T208 = 1'h0;
    1349: T208 = 1'h0;
    1350: T208 = 1'h0;
    1351: T208 = 1'h0;
    1352: T208 = 1'h0;
    1353: T208 = 1'h0;
    1354: T208 = 1'h0;
    1355: T208 = 1'h0;
    1356: T208 = 1'h0;
    1357: T208 = 1'h0;
    1358: T208 = 1'h0;
    1359: T208 = 1'h0;
    1360: T208 = 1'h0;
    1361: T208 = 1'h0;
    1362: T208 = 1'h0;
    1363: T208 = 1'h0;
    1364: T208 = 1'h0;
    1365: T208 = 1'h0;
    1366: T208 = 1'h0;
    1367: T208 = 1'h0;
    1368: T208 = 1'h0;
    1369: T208 = 1'h0;
    1370: T208 = 1'h0;
    1371: T208 = 1'h0;
    1372: T208 = 1'h0;
    1373: T208 = 1'h0;
    1374: T208 = 1'h0;
    1375: T208 = 1'h0;
    1376: T208 = 1'h0;
    1377: T208 = 1'h0;
    1378: T208 = 1'h0;
    1379: T208 = 1'h0;
    1380: T208 = 1'h0;
    1381: T208 = 1'h0;
    1382: T208 = 1'h0;
    1383: T208 = 1'h0;
    1384: T208 = 1'h0;
    1385: T208 = 1'h0;
    1386: T208 = 1'h0;
    1387: T208 = 1'h0;
    1388: T208 = 1'h0;
    1389: T208 = 1'h0;
    1390: T208 = 1'h0;
    1391: T208 = 1'h0;
    1392: T208 = 1'h0;
    1393: T208 = 1'h0;
    1394: T208 = 1'h0;
    1395: T208 = 1'h0;
    1396: T208 = 1'h0;
    1397: T208 = 1'h0;
    1398: T208 = 1'h0;
    1399: T208 = 1'h0;
    1400: T208 = 1'h0;
    1401: T208 = 1'h0;
    1402: T208 = 1'h0;
    1403: T208 = 1'h0;
    1404: T208 = 1'h0;
    1405: T208 = 1'h0;
    1406: T208 = 1'h0;
    1407: T208 = 1'h0;
    1408: T208 = 1'h0;
    1409: T208 = 1'h0;
    1410: T208 = 1'h0;
    1411: T208 = 1'h0;
    1412: T208 = 1'h0;
    1413: T208 = 1'h0;
    1414: T208 = 1'h0;
    1415: T208 = 1'h0;
    1416: T208 = 1'h0;
    1417: T208 = 1'h0;
    1418: T208 = 1'h0;
    1419: T208 = 1'h0;
    1420: T208 = 1'h0;
    1421: T208 = 1'h0;
    1422: T208 = 1'h0;
    1423: T208 = 1'h0;
    1424: T208 = 1'h0;
    1425: T208 = 1'h0;
    1426: T208 = 1'h0;
    1427: T208 = 1'h0;
    1428: T208 = 1'h0;
    1429: T208 = 1'h0;
    1430: T208 = 1'h0;
    1431: T208 = 1'h0;
    1432: T208 = 1'h0;
    1433: T208 = 1'h0;
    1434: T208 = 1'h0;
    1435: T208 = 1'h0;
    1436: T208 = 1'h0;
    1437: T208 = 1'h0;
    1438: T208 = 1'h0;
    1439: T208 = 1'h0;
    1440: T208 = 1'h0;
    1441: T208 = 1'h0;
    1442: T208 = 1'h0;
    1443: T208 = 1'h0;
    1444: T208 = 1'h0;
    1445: T208 = 1'h0;
    1446: T208 = 1'h0;
    1447: T208 = 1'h0;
    1448: T208 = 1'h0;
    1449: T208 = 1'h0;
    1450: T208 = 1'h0;
    1451: T208 = 1'h0;
    1452: T208 = 1'h0;
    1453: T208 = 1'h0;
    1454: T208 = 1'h0;
    1455: T208 = 1'h0;
    1456: T208 = 1'h0;
    1457: T208 = 1'h0;
    1458: T208 = 1'h0;
    1459: T208 = 1'h0;
    1460: T208 = 1'h0;
    1461: T208 = 1'h0;
    1462: T208 = 1'h0;
    1463: T208 = 1'h0;
    1464: T208 = 1'h0;
    1465: T208 = 1'h0;
    1466: T208 = 1'h0;
    1467: T208 = 1'h0;
    1468: T208 = 1'h0;
    1469: T208 = 1'h0;
    1470: T208 = 1'h0;
    1471: T208 = 1'h0;
    1472: T208 = 1'h0;
    1473: T208 = 1'h0;
    1474: T208 = 1'h0;
    1475: T208 = 1'h0;
    1476: T208 = 1'h0;
    1477: T208 = 1'h0;
    1478: T208 = 1'h0;
    1479: T208 = 1'h0;
    1480: T208 = 1'h0;
    1481: T208 = 1'h0;
    1482: T208 = 1'h0;
    1483: T208 = 1'h0;
    1484: T208 = 1'h0;
    1485: T208 = 1'h0;
    1486: T208 = 1'h0;
    1487: T208 = 1'h0;
    1488: T208 = 1'h0;
    1489: T208 = 1'h0;
    1490: T208 = 1'h0;
    1491: T208 = 1'h0;
    1492: T208 = 1'h0;
    1493: T208 = 1'h0;
    1494: T208 = 1'h0;
    1495: T208 = 1'h0;
    1496: T208 = 1'h0;
    1497: T208 = 1'h0;
    1498: T208 = 1'h0;
    1499: T208 = 1'h0;
    1500: T208 = 1'h0;
    1501: T208 = 1'h0;
    1502: T208 = 1'h0;
    1503: T208 = 1'h0;
    1504: T208 = 1'h0;
    1505: T208 = 1'h0;
    1506: T208 = 1'h0;
    1507: T208 = 1'h0;
    1508: T208 = 1'h0;
    1509: T208 = 1'h0;
    1510: T208 = 1'h0;
    1511: T208 = 1'h0;
    1512: T208 = 1'h0;
    1513: T208 = 1'h0;
    1514: T208 = 1'h0;
    1515: T208 = 1'h0;
    1516: T208 = 1'h0;
    1517: T208 = 1'h0;
    1518: T208 = 1'h0;
    1519: T208 = 1'h0;
    1520: T208 = 1'h0;
    1521: T208 = 1'h0;
    1522: T208 = 1'h0;
    1523: T208 = 1'h0;
    1524: T208 = 1'h0;
    1525: T208 = 1'h0;
    1526: T208 = 1'h0;
    1527: T208 = 1'h0;
    1528: T208 = 1'h0;
    1529: T208 = 1'h0;
    1530: T208 = 1'h0;
    1531: T208 = 1'h0;
    1532: T208 = 1'h0;
    1533: T208 = 1'h0;
    1534: T208 = 1'h0;
    1535: T208 = 1'h0;
    1536: T208 = 1'h0;
    1537: T208 = 1'h0;
    1538: T208 = 1'h0;
    1539: T208 = 1'h0;
    1540: T208 = 1'h0;
    1541: T208 = 1'h0;
    1542: T208 = 1'h0;
    1543: T208 = 1'h0;
    1544: T208 = 1'h0;
    1545: T208 = 1'h0;
    1546: T208 = 1'h0;
    1547: T208 = 1'h0;
    1548: T208 = 1'h0;
    1549: T208 = 1'h0;
    1550: T208 = 1'h0;
    1551: T208 = 1'h0;
    1552: T208 = 1'h0;
    1553: T208 = 1'h0;
    1554: T208 = 1'h0;
    1555: T208 = 1'h0;
    1556: T208 = 1'h0;
    1557: T208 = 1'h0;
    1558: T208 = 1'h0;
    1559: T208 = 1'h0;
    1560: T208 = 1'h0;
    1561: T208 = 1'h0;
    1562: T208 = 1'h0;
    1563: T208 = 1'h0;
    1564: T208 = 1'h0;
    1565: T208 = 1'h0;
    1566: T208 = 1'h0;
    1567: T208 = 1'h0;
    1568: T208 = 1'h0;
    1569: T208 = 1'h0;
    1570: T208 = 1'h0;
    1571: T208 = 1'h0;
    1572: T208 = 1'h0;
    1573: T208 = 1'h0;
    1574: T208 = 1'h0;
    1575: T208 = 1'h0;
    1576: T208 = 1'h0;
    1577: T208 = 1'h0;
    1578: T208 = 1'h0;
    1579: T208 = 1'h0;
    1580: T208 = 1'h0;
    1581: T208 = 1'h0;
    1582: T208 = 1'h0;
    1583: T208 = 1'h0;
    1584: T208 = 1'h0;
    1585: T208 = 1'h0;
    1586: T208 = 1'h0;
    1587: T208 = 1'h0;
    1588: T208 = 1'h0;
    1589: T208 = 1'h0;
    1590: T208 = 1'h0;
    1591: T208 = 1'h0;
    1592: T208 = 1'h0;
    1593: T208 = 1'h0;
    1594: T208 = 1'h0;
    1595: T208 = 1'h0;
    1596: T208 = 1'h0;
    1597: T208 = 1'h0;
    1598: T208 = 1'h0;
    1599: T208 = 1'h0;
    1600: T208 = 1'h0;
    1601: T208 = 1'h0;
    1602: T208 = 1'h0;
    1603: T208 = 1'h0;
    1604: T208 = 1'h0;
    1605: T208 = 1'h0;
    1606: T208 = 1'h0;
    1607: T208 = 1'h0;
    1608: T208 = 1'h0;
    1609: T208 = 1'h0;
    1610: T208 = 1'h0;
    1611: T208 = 1'h0;
    1612: T208 = 1'h0;
    1613: T208 = 1'h0;
    1614: T208 = 1'h0;
    1615: T208 = 1'h0;
    1616: T208 = 1'h0;
    1617: T208 = 1'h0;
    1618: T208 = 1'h0;
    1619: T208 = 1'h0;
    1620: T208 = 1'h0;
    1621: T208 = 1'h0;
    1622: T208 = 1'h0;
    1623: T208 = 1'h0;
    1624: T208 = 1'h0;
    1625: T208 = 1'h0;
    1626: T208 = 1'h0;
    1627: T208 = 1'h0;
    1628: T208 = 1'h0;
    1629: T208 = 1'h0;
    1630: T208 = 1'h0;
    1631: T208 = 1'h0;
    1632: T208 = 1'h0;
    1633: T208 = 1'h0;
    1634: T208 = 1'h0;
    1635: T208 = 1'h0;
    1636: T208 = 1'h0;
    1637: T208 = 1'h0;
    1638: T208 = 1'h0;
    1639: T208 = 1'h0;
    1640: T208 = 1'h0;
    1641: T208 = 1'h0;
    1642: T208 = 1'h0;
    1643: T208 = 1'h0;
    1644: T208 = 1'h0;
    1645: T208 = 1'h0;
    1646: T208 = 1'h0;
    1647: T208 = 1'h0;
    1648: T208 = 1'h0;
    1649: T208 = 1'h0;
    1650: T208 = 1'h0;
    1651: T208 = 1'h0;
    1652: T208 = 1'h0;
    1653: T208 = 1'h0;
    1654: T208 = 1'h0;
    1655: T208 = 1'h0;
    1656: T208 = 1'h0;
    1657: T208 = 1'h0;
    1658: T208 = 1'h0;
    1659: T208 = 1'h0;
    1660: T208 = 1'h0;
    1661: T208 = 1'h0;
    1662: T208 = 1'h0;
    1663: T208 = 1'h0;
    1664: T208 = 1'h0;
    1665: T208 = 1'h0;
    1666: T208 = 1'h0;
    1667: T208 = 1'h0;
    1668: T208 = 1'h0;
    1669: T208 = 1'h0;
    1670: T208 = 1'h0;
    1671: T208 = 1'h0;
    1672: T208 = 1'h0;
    1673: T208 = 1'h0;
    1674: T208 = 1'h0;
    1675: T208 = 1'h0;
    1676: T208 = 1'h0;
    1677: T208 = 1'h0;
    1678: T208 = 1'h0;
    1679: T208 = 1'h0;
    1680: T208 = 1'h0;
    1681: T208 = 1'h0;
    1682: T208 = 1'h0;
    1683: T208 = 1'h0;
    1684: T208 = 1'h0;
    1685: T208 = 1'h0;
    1686: T208 = 1'h0;
    1687: T208 = 1'h0;
    1688: T208 = 1'h0;
    1689: T208 = 1'h0;
    1690: T208 = 1'h0;
    1691: T208 = 1'h0;
    1692: T208 = 1'h0;
    1693: T208 = 1'h0;
    1694: T208 = 1'h0;
    1695: T208 = 1'h0;
    1696: T208 = 1'h0;
    1697: T208 = 1'h0;
    1698: T208 = 1'h0;
    1699: T208 = 1'h0;
    1700: T208 = 1'h0;
    1701: T208 = 1'h0;
    1702: T208 = 1'h0;
    1703: T208 = 1'h0;
    1704: T208 = 1'h0;
    1705: T208 = 1'h0;
    1706: T208 = 1'h0;
    1707: T208 = 1'h0;
    1708: T208 = 1'h0;
    1709: T208 = 1'h0;
    1710: T208 = 1'h0;
    1711: T208 = 1'h0;
    1712: T208 = 1'h0;
    1713: T208 = 1'h0;
    1714: T208 = 1'h0;
    1715: T208 = 1'h0;
    1716: T208 = 1'h0;
    1717: T208 = 1'h0;
    1718: T208 = 1'h0;
    1719: T208 = 1'h0;
    1720: T208 = 1'h0;
    1721: T208 = 1'h0;
    1722: T208 = 1'h0;
    1723: T208 = 1'h0;
    1724: T208 = 1'h0;
    1725: T208 = 1'h0;
    1726: T208 = 1'h0;
    1727: T208 = 1'h0;
    1728: T208 = 1'h0;
    1729: T208 = 1'h0;
    1730: T208 = 1'h0;
    1731: T208 = 1'h0;
    1732: T208 = 1'h0;
    1733: T208 = 1'h0;
    1734: T208 = 1'h0;
    1735: T208 = 1'h0;
    1736: T208 = 1'h0;
    1737: T208 = 1'h0;
    1738: T208 = 1'h0;
    1739: T208 = 1'h0;
    1740: T208 = 1'h0;
    1741: T208 = 1'h0;
    1742: T208 = 1'h0;
    1743: T208 = 1'h0;
    1744: T208 = 1'h0;
    1745: T208 = 1'h0;
    1746: T208 = 1'h0;
    1747: T208 = 1'h0;
    1748: T208 = 1'h0;
    1749: T208 = 1'h0;
    1750: T208 = 1'h0;
    1751: T208 = 1'h0;
    1752: T208 = 1'h0;
    1753: T208 = 1'h0;
    1754: T208 = 1'h0;
    1755: T208 = 1'h0;
    1756: T208 = 1'h0;
    1757: T208 = 1'h0;
    1758: T208 = 1'h0;
    1759: T208 = 1'h0;
    1760: T208 = 1'h0;
    1761: T208 = 1'h0;
    1762: T208 = 1'h0;
    1763: T208 = 1'h0;
    1764: T208 = 1'h0;
    1765: T208 = 1'h0;
    1766: T208 = 1'h0;
    1767: T208 = 1'h0;
    1768: T208 = 1'h0;
    1769: T208 = 1'h0;
    1770: T208 = 1'h0;
    1771: T208 = 1'h0;
    1772: T208 = 1'h0;
    1773: T208 = 1'h0;
    1774: T208 = 1'h0;
    1775: T208 = 1'h0;
    1776: T208 = 1'h0;
    1777: T208 = 1'h0;
    1778: T208 = 1'h0;
    1779: T208 = 1'h0;
    1780: T208 = 1'h0;
    1781: T208 = 1'h0;
    1782: T208 = 1'h0;
    1783: T208 = 1'h0;
    1784: T208 = 1'h0;
    1785: T208 = 1'h0;
    1786: T208 = 1'h0;
    1787: T208 = 1'h0;
    1788: T208 = 1'h0;
    1789: T208 = 1'h0;
    1790: T208 = 1'h0;
    1791: T208 = 1'h0;
    1792: T208 = 1'h0;
    1793: T208 = 1'h0;
    1794: T208 = 1'h0;
    1795: T208 = 1'h0;
    1796: T208 = 1'h0;
    1797: T208 = 1'h0;
    1798: T208 = 1'h0;
    1799: T208 = 1'h0;
    1800: T208 = 1'h0;
    1801: T208 = 1'h0;
    1802: T208 = 1'h0;
    1803: T208 = 1'h0;
    1804: T208 = 1'h0;
    1805: T208 = 1'h0;
    1806: T208 = 1'h0;
    1807: T208 = 1'h0;
    1808: T208 = 1'h0;
    1809: T208 = 1'h0;
    1810: T208 = 1'h0;
    1811: T208 = 1'h0;
    1812: T208 = 1'h0;
    1813: T208 = 1'h0;
    1814: T208 = 1'h0;
    1815: T208 = 1'h0;
    1816: T208 = 1'h0;
    1817: T208 = 1'h0;
    1818: T208 = 1'h0;
    1819: T208 = 1'h0;
    1820: T208 = 1'h0;
    1821: T208 = 1'h0;
    1822: T208 = 1'h0;
    1823: T208 = 1'h0;
    1824: T208 = 1'h0;
    1825: T208 = 1'h0;
    1826: T208 = 1'h0;
    1827: T208 = 1'h0;
    1828: T208 = 1'h0;
    1829: T208 = 1'h0;
    1830: T208 = 1'h0;
    1831: T208 = 1'h0;
    1832: T208 = 1'h0;
    1833: T208 = 1'h0;
    1834: T208 = 1'h0;
    1835: T208 = 1'h0;
    1836: T208 = 1'h0;
    1837: T208 = 1'h0;
    1838: T208 = 1'h0;
    1839: T208 = 1'h0;
    1840: T208 = 1'h0;
    1841: T208 = 1'h0;
    1842: T208 = 1'h0;
    1843: T208 = 1'h0;
    1844: T208 = 1'h0;
    1845: T208 = 1'h0;
    1846: T208 = 1'h0;
    1847: T208 = 1'h0;
    1848: T208 = 1'h0;
    1849: T208 = 1'h0;
    1850: T208 = 1'h0;
    1851: T208 = 1'h0;
    1852: T208 = 1'h0;
    1853: T208 = 1'h0;
    1854: T208 = 1'h0;
    1855: T208 = 1'h0;
    1856: T208 = 1'h0;
    1857: T208 = 1'h0;
    1858: T208 = 1'h0;
    1859: T208 = 1'h0;
    1860: T208 = 1'h0;
    1861: T208 = 1'h0;
    1862: T208 = 1'h0;
    1863: T208 = 1'h0;
    1864: T208 = 1'h0;
    1865: T208 = 1'h0;
    1866: T208 = 1'h0;
    1867: T208 = 1'h0;
    1868: T208 = 1'h0;
    1869: T208 = 1'h0;
    1870: T208 = 1'h0;
    1871: T208 = 1'h0;
    1872: T208 = 1'h0;
    1873: T208 = 1'h0;
    1874: T208 = 1'h0;
    1875: T208 = 1'h0;
    1876: T208 = 1'h0;
    1877: T208 = 1'h0;
    1878: T208 = 1'h0;
    1879: T208 = 1'h0;
    1880: T208 = 1'h0;
    1881: T208 = 1'h0;
    1882: T208 = 1'h0;
    1883: T208 = 1'h0;
    1884: T208 = 1'h0;
    1885: T208 = 1'h0;
    1886: T208 = 1'h0;
    1887: T208 = 1'h0;
    1888: T208 = 1'h0;
    1889: T208 = 1'h0;
    1890: T208 = 1'h0;
    1891: T208 = 1'h0;
    1892: T208 = 1'h0;
    1893: T208 = 1'h0;
    1894: T208 = 1'h0;
    1895: T208 = 1'h0;
    1896: T208 = 1'h0;
    1897: T208 = 1'h0;
    1898: T208 = 1'h0;
    1899: T208 = 1'h0;
    1900: T208 = 1'h0;
    1901: T208 = 1'h0;
    1902: T208 = 1'h0;
    1903: T208 = 1'h0;
    1904: T208 = 1'h0;
    1905: T208 = 1'h0;
    1906: T208 = 1'h0;
    1907: T208 = 1'h0;
    1908: T208 = 1'h0;
    1909: T208 = 1'h0;
    1910: T208 = 1'h0;
    1911: T208 = 1'h0;
    1912: T208 = 1'h0;
    1913: T208 = 1'h0;
    1914: T208 = 1'h0;
    1915: T208 = 1'h0;
    1916: T208 = 1'h0;
    1917: T208 = 1'h0;
    1918: T208 = 1'h0;
    1919: T208 = 1'h0;
    1920: T208 = 1'h0;
    1921: T208 = 1'h0;
    1922: T208 = 1'h0;
    1923: T208 = 1'h0;
    1924: T208 = 1'h0;
    1925: T208 = 1'h0;
    1926: T208 = 1'h0;
    1927: T208 = 1'h0;
    1928: T208 = 1'h0;
    1929: T208 = 1'h0;
    1930: T208 = 1'h0;
    1931: T208 = 1'h0;
    1932: T208 = 1'h0;
    1933: T208 = 1'h0;
    1934: T208 = 1'h0;
    1935: T208 = 1'h0;
    1936: T208 = 1'h0;
    1937: T208 = 1'h0;
    1938: T208 = 1'h0;
    1939: T208 = 1'h0;
    1940: T208 = 1'h0;
    1941: T208 = 1'h0;
    1942: T208 = 1'h0;
    1943: T208 = 1'h0;
    1944: T208 = 1'h0;
    1945: T208 = 1'h0;
    1946: T208 = 1'h0;
    1947: T208 = 1'h0;
    1948: T208 = 1'h0;
    1949: T208 = 1'h0;
    1950: T208 = 1'h0;
    1951: T208 = 1'h0;
    1952: T208 = 1'h0;
    1953: T208 = 1'h0;
    1954: T208 = 1'h0;
    1955: T208 = 1'h0;
    1956: T208 = 1'h0;
    1957: T208 = 1'h0;
    1958: T208 = 1'h0;
    1959: T208 = 1'h0;
    1960: T208 = 1'h0;
    1961: T208 = 1'h0;
    1962: T208 = 1'h0;
    1963: T208 = 1'h0;
    1964: T208 = 1'h0;
    1965: T208 = 1'h0;
    1966: T208 = 1'h0;
    1967: T208 = 1'h0;
    1968: T208 = 1'h0;
    1969: T208 = 1'h0;
    1970: T208 = 1'h0;
    1971: T208 = 1'h0;
    1972: T208 = 1'h0;
    1973: T208 = 1'h0;
    1974: T208 = 1'h0;
    1975: T208 = 1'h0;
    1976: T208 = 1'h0;
    1977: T208 = 1'h0;
    1978: T208 = 1'h0;
    1979: T208 = 1'h0;
    1980: T208 = 1'h0;
    1981: T208 = 1'h0;
    1982: T208 = 1'h0;
    1983: T208 = 1'h0;
    1984: T208 = 1'h0;
    1985: T208 = 1'h0;
    1986: T208 = 1'h0;
    1987: T208 = 1'h0;
    1988: T208 = 1'h0;
    1989: T208 = 1'h0;
    1990: T208 = 1'h0;
    1991: T208 = 1'h0;
    1992: T208 = 1'h0;
    1993: T208 = 1'h0;
    1994: T208 = 1'h0;
    1995: T208 = 1'h0;
    1996: T208 = 1'h0;
    1997: T208 = 1'h0;
    1998: T208 = 1'h0;
    1999: T208 = 1'h0;
    2000: T208 = 1'h0;
    2001: T208 = 1'h0;
    2002: T208 = 1'h0;
    2003: T208 = 1'h0;
    2004: T208 = 1'h0;
    2005: T208 = 1'h0;
    2006: T208 = 1'h0;
    2007: T208 = 1'h0;
    2008: T208 = 1'h0;
    2009: T208 = 1'h0;
    2010: T208 = 1'h0;
    2011: T208 = 1'h0;
    2012: T208 = 1'h0;
    2013: T208 = 1'h0;
    2014: T208 = 1'h0;
    2015: T208 = 1'h0;
    2016: T208 = 1'h0;
    2017: T208 = 1'h0;
    2018: T208 = 1'h0;
    2019: T208 = 1'h0;
    2020: T208 = 1'h0;
    2021: T208 = 1'h0;
    2022: T208 = 1'h0;
    2023: T208 = 1'h0;
    2024: T208 = 1'h0;
    2025: T208 = 1'h0;
    2026: T208 = 1'h0;
    2027: T208 = 1'h0;
    2028: T208 = 1'h0;
    2029: T208 = 1'h0;
    2030: T208 = 1'h0;
    2031: T208 = 1'h0;
    2032: T208 = 1'h0;
    2033: T208 = 1'h0;
    2034: T208 = 1'h0;
    2035: T208 = 1'h0;
    2036: T208 = 1'h0;
    2037: T208 = 1'h0;
    2038: T208 = 1'h0;
    2039: T208 = 1'h0;
    2040: T208 = 1'h0;
    2041: T208 = 1'h0;
    2042: T208 = 1'h0;
    2043: T208 = 1'h0;
    2044: T208 = 1'h0;
    2045: T208 = 1'h0;
    2046: T208 = 1'h0;
    2047: T208 = 1'h0;
    2048: T208 = 1'h0;
    2049: T208 = 1'h0;
    2050: T208 = 1'h0;
    2051: T208 = 1'h0;
    2052: T208 = 1'h0;
    2053: T208 = 1'h0;
    2054: T208 = 1'h0;
    2055: T208 = 1'h0;
    2056: T208 = 1'h0;
    2057: T208 = 1'h0;
    2058: T208 = 1'h0;
    2059: T208 = 1'h0;
    2060: T208 = 1'h0;
    2061: T208 = 1'h0;
    2062: T208 = 1'h0;
    2063: T208 = 1'h0;
    2064: T208 = 1'h0;
    2065: T208 = 1'h0;
    2066: T208 = 1'h0;
    2067: T208 = 1'h0;
    2068: T208 = 1'h0;
    2069: T208 = 1'h0;
    2070: T208 = 1'h0;
    2071: T208 = 1'h0;
    2072: T208 = 1'h0;
    2073: T208 = 1'h0;
    2074: T208 = 1'h0;
    2075: T208 = 1'h0;
    2076: T208 = 1'h0;
    2077: T208 = 1'h0;
    2078: T208 = 1'h0;
    2079: T208 = 1'h0;
    2080: T208 = 1'h0;
    2081: T208 = 1'h0;
    2082: T208 = 1'h0;
    2083: T208 = 1'h0;
    2084: T208 = 1'h0;
    2085: T208 = 1'h0;
    2086: T208 = 1'h0;
    2087: T208 = 1'h0;
    2088: T208 = 1'h0;
    2089: T208 = 1'h0;
    2090: T208 = 1'h0;
    2091: T208 = 1'h0;
    2092: T208 = 1'h0;
    2093: T208 = 1'h0;
    2094: T208 = 1'h0;
    2095: T208 = 1'h0;
    2096: T208 = 1'h0;
    2097: T208 = 1'h0;
    2098: T208 = 1'h0;
    2099: T208 = 1'h0;
    2100: T208 = 1'h0;
    2101: T208 = 1'h0;
    2102: T208 = 1'h0;
    2103: T208 = 1'h0;
    2104: T208 = 1'h0;
    2105: T208 = 1'h0;
    2106: T208 = 1'h0;
    2107: T208 = 1'h0;
    2108: T208 = 1'h0;
    2109: T208 = 1'h0;
    2110: T208 = 1'h0;
    2111: T208 = 1'h0;
    2112: T208 = 1'h0;
    2113: T208 = 1'h0;
    2114: T208 = 1'h0;
    2115: T208 = 1'h0;
    2116: T208 = 1'h0;
    2117: T208 = 1'h0;
    2118: T208 = 1'h0;
    2119: T208 = 1'h0;
    2120: T208 = 1'h0;
    2121: T208 = 1'h0;
    2122: T208 = 1'h0;
    2123: T208 = 1'h0;
    2124: T208 = 1'h0;
    2125: T208 = 1'h0;
    2126: T208 = 1'h0;
    2127: T208 = 1'h0;
    2128: T208 = 1'h0;
    2129: T208 = 1'h0;
    2130: T208 = 1'h0;
    2131: T208 = 1'h0;
    2132: T208 = 1'h0;
    2133: T208 = 1'h0;
    2134: T208 = 1'h0;
    2135: T208 = 1'h0;
    2136: T208 = 1'h0;
    2137: T208 = 1'h0;
    2138: T208 = 1'h0;
    2139: T208 = 1'h0;
    2140: T208 = 1'h0;
    2141: T208 = 1'h0;
    2142: T208 = 1'h0;
    2143: T208 = 1'h0;
    2144: T208 = 1'h0;
    2145: T208 = 1'h0;
    2146: T208 = 1'h0;
    2147: T208 = 1'h0;
    2148: T208 = 1'h0;
    2149: T208 = 1'h0;
    2150: T208 = 1'h0;
    2151: T208 = 1'h0;
    2152: T208 = 1'h0;
    2153: T208 = 1'h0;
    2154: T208 = 1'h0;
    2155: T208 = 1'h0;
    2156: T208 = 1'h0;
    2157: T208 = 1'h0;
    2158: T208 = 1'h0;
    2159: T208 = 1'h0;
    2160: T208 = 1'h0;
    2161: T208 = 1'h0;
    2162: T208 = 1'h0;
    2163: T208 = 1'h0;
    2164: T208 = 1'h0;
    2165: T208 = 1'h0;
    2166: T208 = 1'h0;
    2167: T208 = 1'h0;
    2168: T208 = 1'h0;
    2169: T208 = 1'h0;
    2170: T208 = 1'h0;
    2171: T208 = 1'h0;
    2172: T208 = 1'h0;
    2173: T208 = 1'h0;
    2174: T208 = 1'h0;
    2175: T208 = 1'h0;
    2176: T208 = 1'h0;
    2177: T208 = 1'h0;
    2178: T208 = 1'h0;
    2179: T208 = 1'h0;
    2180: T208 = 1'h0;
    2181: T208 = 1'h0;
    2182: T208 = 1'h0;
    2183: T208 = 1'h0;
    2184: T208 = 1'h0;
    2185: T208 = 1'h0;
    2186: T208 = 1'h0;
    2187: T208 = 1'h0;
    2188: T208 = 1'h0;
    2189: T208 = 1'h0;
    2190: T208 = 1'h0;
    2191: T208 = 1'h0;
    2192: T208 = 1'h0;
    2193: T208 = 1'h0;
    2194: T208 = 1'h0;
    2195: T208 = 1'h0;
    2196: T208 = 1'h0;
    2197: T208 = 1'h0;
    2198: T208 = 1'h0;
    2199: T208 = 1'h0;
    2200: T208 = 1'h0;
    2201: T208 = 1'h0;
    2202: T208 = 1'h0;
    2203: T208 = 1'h0;
    2204: T208 = 1'h0;
    2205: T208 = 1'h0;
    2206: T208 = 1'h0;
    2207: T208 = 1'h0;
    2208: T208 = 1'h0;
    2209: T208 = 1'h0;
    2210: T208 = 1'h0;
    2211: T208 = 1'h0;
    2212: T208 = 1'h0;
    2213: T208 = 1'h0;
    2214: T208 = 1'h0;
    2215: T208 = 1'h0;
    2216: T208 = 1'h0;
    2217: T208 = 1'h0;
    2218: T208 = 1'h0;
    2219: T208 = 1'h0;
    2220: T208 = 1'h0;
    2221: T208 = 1'h0;
    2222: T208 = 1'h0;
    2223: T208 = 1'h0;
    2224: T208 = 1'h0;
    2225: T208 = 1'h0;
    2226: T208 = 1'h0;
    2227: T208 = 1'h0;
    2228: T208 = 1'h0;
    2229: T208 = 1'h0;
    2230: T208 = 1'h0;
    2231: T208 = 1'h0;
    2232: T208 = 1'h0;
    2233: T208 = 1'h0;
    2234: T208 = 1'h0;
    2235: T208 = 1'h0;
    2236: T208 = 1'h0;
    2237: T208 = 1'h0;
    2238: T208 = 1'h0;
    2239: T208 = 1'h0;
    2240: T208 = 1'h0;
    2241: T208 = 1'h0;
    2242: T208 = 1'h0;
    2243: T208 = 1'h0;
    2244: T208 = 1'h0;
    2245: T208 = 1'h0;
    2246: T208 = 1'h0;
    2247: T208 = 1'h0;
    2248: T208 = 1'h0;
    2249: T208 = 1'h0;
    2250: T208 = 1'h0;
    2251: T208 = 1'h0;
    2252: T208 = 1'h0;
    2253: T208 = 1'h0;
    2254: T208 = 1'h0;
    2255: T208 = 1'h0;
    2256: T208 = 1'h0;
    2257: T208 = 1'h0;
    2258: T208 = 1'h0;
    2259: T208 = 1'h0;
    2260: T208 = 1'h0;
    2261: T208 = 1'h0;
    2262: T208 = 1'h0;
    2263: T208 = 1'h0;
    2264: T208 = 1'h0;
    2265: T208 = 1'h0;
    2266: T208 = 1'h0;
    2267: T208 = 1'h0;
    2268: T208 = 1'h0;
    2269: T208 = 1'h0;
    2270: T208 = 1'h0;
    2271: T208 = 1'h0;
    2272: T208 = 1'h0;
    2273: T208 = 1'h0;
    2274: T208 = 1'h0;
    2275: T208 = 1'h0;
    2276: T208 = 1'h0;
    2277: T208 = 1'h0;
    2278: T208 = 1'h0;
    2279: T208 = 1'h0;
    2280: T208 = 1'h0;
    2281: T208 = 1'h0;
    2282: T208 = 1'h0;
    2283: T208 = 1'h0;
    2284: T208 = 1'h0;
    2285: T208 = 1'h0;
    2286: T208 = 1'h0;
    2287: T208 = 1'h0;
    2288: T208 = 1'h0;
    2289: T208 = 1'h0;
    2290: T208 = 1'h0;
    2291: T208 = 1'h0;
    2292: T208 = 1'h0;
    2293: T208 = 1'h0;
    2294: T208 = 1'h0;
    2295: T208 = 1'h0;
    2296: T208 = 1'h0;
    2297: T208 = 1'h0;
    2298: T208 = 1'h0;
    2299: T208 = 1'h0;
    2300: T208 = 1'h0;
    2301: T208 = 1'h0;
    2302: T208 = 1'h0;
    2303: T208 = 1'h0;
    2304: T208 = 1'h0;
    2305: T208 = 1'h0;
    2306: T208 = 1'h0;
    2307: T208 = 1'h0;
    2308: T208 = 1'h0;
    2309: T208 = 1'h0;
    2310: T208 = 1'h0;
    2311: T208 = 1'h0;
    2312: T208 = 1'h0;
    2313: T208 = 1'h0;
    2314: T208 = 1'h0;
    2315: T208 = 1'h0;
    2316: T208 = 1'h0;
    2317: T208 = 1'h0;
    2318: T208 = 1'h0;
    2319: T208 = 1'h0;
    2320: T208 = 1'h0;
    2321: T208 = 1'h0;
    2322: T208 = 1'h0;
    2323: T208 = 1'h0;
    2324: T208 = 1'h0;
    2325: T208 = 1'h0;
    2326: T208 = 1'h0;
    2327: T208 = 1'h0;
    2328: T208 = 1'h0;
    2329: T208 = 1'h0;
    2330: T208 = 1'h0;
    2331: T208 = 1'h0;
    2332: T208 = 1'h0;
    2333: T208 = 1'h0;
    2334: T208 = 1'h0;
    2335: T208 = 1'h0;
    2336: T208 = 1'h0;
    2337: T208 = 1'h0;
    2338: T208 = 1'h0;
    2339: T208 = 1'h0;
    2340: T208 = 1'h0;
    2341: T208 = 1'h0;
    2342: T208 = 1'h0;
    2343: T208 = 1'h0;
    2344: T208 = 1'h0;
    2345: T208 = 1'h0;
    2346: T208 = 1'h0;
    2347: T208 = 1'h0;
    2348: T208 = 1'h0;
    2349: T208 = 1'h0;
    2350: T208 = 1'h0;
    2351: T208 = 1'h0;
    2352: T208 = 1'h0;
    2353: T208 = 1'h0;
    2354: T208 = 1'h0;
    2355: T208 = 1'h0;
    2356: T208 = 1'h0;
    2357: T208 = 1'h0;
    2358: T208 = 1'h0;
    2359: T208 = 1'h0;
    2360: T208 = 1'h0;
    2361: T208 = 1'h0;
    2362: T208 = 1'h0;
    2363: T208 = 1'h0;
    2364: T208 = 1'h0;
    2365: T208 = 1'h0;
    2366: T208 = 1'h0;
    2367: T208 = 1'h0;
    2368: T208 = 1'h0;
    2369: T208 = 1'h0;
    2370: T208 = 1'h0;
    2371: T208 = 1'h0;
    2372: T208 = 1'h0;
    2373: T208 = 1'h0;
    2374: T208 = 1'h0;
    2375: T208 = 1'h0;
    2376: T208 = 1'h0;
    2377: T208 = 1'h0;
    2378: T208 = 1'h0;
    2379: T208 = 1'h0;
    2380: T208 = 1'h0;
    2381: T208 = 1'h0;
    2382: T208 = 1'h0;
    2383: T208 = 1'h0;
    2384: T208 = 1'h0;
    2385: T208 = 1'h0;
    2386: T208 = 1'h0;
    2387: T208 = 1'h0;
    2388: T208 = 1'h0;
    2389: T208 = 1'h0;
    2390: T208 = 1'h0;
    2391: T208 = 1'h0;
    2392: T208 = 1'h0;
    2393: T208 = 1'h0;
    2394: T208 = 1'h0;
    2395: T208 = 1'h0;
    2396: T208 = 1'h0;
    2397: T208 = 1'h0;
    2398: T208 = 1'h0;
    2399: T208 = 1'h0;
    2400: T208 = 1'h0;
    2401: T208 = 1'h0;
    2402: T208 = 1'h0;
    2403: T208 = 1'h0;
    2404: T208 = 1'h0;
    2405: T208 = 1'h0;
    2406: T208 = 1'h0;
    2407: T208 = 1'h0;
    2408: T208 = 1'h0;
    2409: T208 = 1'h0;
    2410: T208 = 1'h0;
    2411: T208 = 1'h0;
    2412: T208 = 1'h0;
    2413: T208 = 1'h0;
    2414: T208 = 1'h0;
    2415: T208 = 1'h0;
    2416: T208 = 1'h0;
    2417: T208 = 1'h0;
    2418: T208 = 1'h0;
    2419: T208 = 1'h0;
    2420: T208 = 1'h0;
    2421: T208 = 1'h0;
    2422: T208 = 1'h0;
    2423: T208 = 1'h0;
    2424: T208 = 1'h0;
    2425: T208 = 1'h0;
    2426: T208 = 1'h0;
    2427: T208 = 1'h0;
    2428: T208 = 1'h0;
    2429: T208 = 1'h0;
    2430: T208 = 1'h0;
    2431: T208 = 1'h0;
    2432: T208 = 1'h0;
    2433: T208 = 1'h0;
    2434: T208 = 1'h0;
    2435: T208 = 1'h0;
    2436: T208 = 1'h0;
    2437: T208 = 1'h0;
    2438: T208 = 1'h0;
    2439: T208 = 1'h0;
    2440: T208 = 1'h0;
    2441: T208 = 1'h0;
    2442: T208 = 1'h0;
    2443: T208 = 1'h0;
    2444: T208 = 1'h0;
    2445: T208 = 1'h0;
    2446: T208 = 1'h0;
    2447: T208 = 1'h0;
    2448: T208 = 1'h0;
    2449: T208 = 1'h0;
    2450: T208 = 1'h0;
    2451: T208 = 1'h0;
    2452: T208 = 1'h0;
    2453: T208 = 1'h0;
    2454: T208 = 1'h0;
    2455: T208 = 1'h0;
    2456: T208 = 1'h0;
    2457: T208 = 1'h0;
    2458: T208 = 1'h0;
    2459: T208 = 1'h0;
    2460: T208 = 1'h0;
    2461: T208 = 1'h0;
    2462: T208 = 1'h0;
    2463: T208 = 1'h0;
    2464: T208 = 1'h0;
    2465: T208 = 1'h0;
    2466: T208 = 1'h0;
    2467: T208 = 1'h0;
    2468: T208 = 1'h0;
    2469: T208 = 1'h0;
    2470: T208 = 1'h0;
    2471: T208 = 1'h0;
    2472: T208 = 1'h0;
    2473: T208 = 1'h0;
    2474: T208 = 1'h0;
    2475: T208 = 1'h0;
    2476: T208 = 1'h0;
    2477: T208 = 1'h0;
    2478: T208 = 1'h0;
    2479: T208 = 1'h0;
    2480: T208 = 1'h0;
    2481: T208 = 1'h0;
    2482: T208 = 1'h0;
    2483: T208 = 1'h0;
    2484: T208 = 1'h0;
    2485: T208 = 1'h0;
    2486: T208 = 1'h0;
    2487: T208 = 1'h0;
    2488: T208 = 1'h0;
    2489: T208 = 1'h0;
    2490: T208 = 1'h0;
    2491: T208 = 1'h0;
    2492: T208 = 1'h0;
    2493: T208 = 1'h0;
    2494: T208 = 1'h0;
    2495: T208 = 1'h0;
    2496: T208 = 1'h0;
    2497: T208 = 1'h0;
    2498: T208 = 1'h0;
    2499: T208 = 1'h0;
    2500: T208 = 1'h0;
    2501: T208 = 1'h0;
    2502: T208 = 1'h0;
    2503: T208 = 1'h0;
    2504: T208 = 1'h0;
    2505: T208 = 1'h0;
    2506: T208 = 1'h0;
    2507: T208 = 1'h0;
    2508: T208 = 1'h0;
    2509: T208 = 1'h0;
    2510: T208 = 1'h0;
    2511: T208 = 1'h0;
    2512: T208 = 1'h0;
    2513: T208 = 1'h0;
    2514: T208 = 1'h0;
    2515: T208 = 1'h0;
    2516: T208 = 1'h0;
    2517: T208 = 1'h0;
    2518: T208 = 1'h0;
    2519: T208 = 1'h0;
    2520: T208 = 1'h0;
    2521: T208 = 1'h0;
    2522: T208 = 1'h0;
    2523: T208 = 1'h0;
    2524: T208 = 1'h0;
    2525: T208 = 1'h0;
    2526: T208 = 1'h0;
    2527: T208 = 1'h0;
    2528: T208 = 1'h0;
    2529: T208 = 1'h0;
    2530: T208 = 1'h0;
    2531: T208 = 1'h0;
    2532: T208 = 1'h0;
    2533: T208 = 1'h0;
    2534: T208 = 1'h0;
    2535: T208 = 1'h0;
    2536: T208 = 1'h0;
    2537: T208 = 1'h0;
    2538: T208 = 1'h0;
    2539: T208 = 1'h0;
    2540: T208 = 1'h0;
    2541: T208 = 1'h0;
    2542: T208 = 1'h0;
    2543: T208 = 1'h0;
    2544: T208 = 1'h0;
    2545: T208 = 1'h0;
    2546: T208 = 1'h0;
    2547: T208 = 1'h0;
    2548: T208 = 1'h0;
    2549: T208 = 1'h0;
    2550: T208 = 1'h0;
    2551: T208 = 1'h0;
    2552: T208 = 1'h0;
    2553: T208 = 1'h0;
    2554: T208 = 1'h0;
    2555: T208 = 1'h0;
    2556: T208 = 1'h0;
    2557: T208 = 1'h0;
    2558: T208 = 1'h0;
    2559: T208 = 1'h0;
    2560: T208 = 1'h0;
    2561: T208 = 1'h0;
    2562: T208 = 1'h0;
    2563: T208 = 1'h0;
    2564: T208 = 1'h0;
    2565: T208 = 1'h0;
    2566: T208 = 1'h0;
    2567: T208 = 1'h0;
    2568: T208 = 1'h0;
    2569: T208 = 1'h0;
    2570: T208 = 1'h0;
    2571: T208 = 1'h0;
    2572: T208 = 1'h0;
    2573: T208 = 1'h0;
    2574: T208 = 1'h0;
    2575: T208 = 1'h0;
    2576: T208 = 1'h0;
    2577: T208 = 1'h0;
    2578: T208 = 1'h0;
    2579: T208 = 1'h0;
    2580: T208 = 1'h0;
    2581: T208 = 1'h0;
    2582: T208 = 1'h0;
    2583: T208 = 1'h0;
    2584: T208 = 1'h0;
    2585: T208 = 1'h0;
    2586: T208 = 1'h0;
    2587: T208 = 1'h0;
    2588: T208 = 1'h0;
    2589: T208 = 1'h0;
    2590: T208 = 1'h0;
    2591: T208 = 1'h0;
    2592: T208 = 1'h0;
    2593: T208 = 1'h0;
    2594: T208 = 1'h0;
    2595: T208 = 1'h0;
    2596: T208 = 1'h0;
    2597: T208 = 1'h0;
    2598: T208 = 1'h0;
    2599: T208 = 1'h0;
    2600: T208 = 1'h0;
    2601: T208 = 1'h0;
    2602: T208 = 1'h0;
    2603: T208 = 1'h0;
    2604: T208 = 1'h0;
    2605: T208 = 1'h0;
    2606: T208 = 1'h0;
    2607: T208 = 1'h0;
    2608: T208 = 1'h0;
    2609: T208 = 1'h0;
    2610: T208 = 1'h0;
    2611: T208 = 1'h0;
    2612: T208 = 1'h0;
    2613: T208 = 1'h0;
    2614: T208 = 1'h0;
    2615: T208 = 1'h0;
    2616: T208 = 1'h0;
    2617: T208 = 1'h0;
    2618: T208 = 1'h0;
    2619: T208 = 1'h0;
    2620: T208 = 1'h0;
    2621: T208 = 1'h0;
    2622: T208 = 1'h0;
    2623: T208 = 1'h0;
    2624: T208 = 1'h0;
    2625: T208 = 1'h0;
    2626: T208 = 1'h0;
    2627: T208 = 1'h0;
    2628: T208 = 1'h0;
    2629: T208 = 1'h0;
    2630: T208 = 1'h0;
    2631: T208 = 1'h0;
    2632: T208 = 1'h0;
    2633: T208 = 1'h0;
    2634: T208 = 1'h0;
    2635: T208 = 1'h0;
    2636: T208 = 1'h0;
    2637: T208 = 1'h0;
    2638: T208 = 1'h0;
    2639: T208 = 1'h0;
    2640: T208 = 1'h0;
    2641: T208 = 1'h0;
    2642: T208 = 1'h0;
    2643: T208 = 1'h0;
    2644: T208 = 1'h0;
    2645: T208 = 1'h0;
    2646: T208 = 1'h0;
    2647: T208 = 1'h0;
    2648: T208 = 1'h0;
    2649: T208 = 1'h0;
    2650: T208 = 1'h0;
    2651: T208 = 1'h0;
    2652: T208 = 1'h0;
    2653: T208 = 1'h0;
    2654: T208 = 1'h0;
    2655: T208 = 1'h0;
    2656: T208 = 1'h0;
    2657: T208 = 1'h0;
    2658: T208 = 1'h0;
    2659: T208 = 1'h0;
    2660: T208 = 1'h0;
    2661: T208 = 1'h0;
    2662: T208 = 1'h0;
    2663: T208 = 1'h0;
    2664: T208 = 1'h0;
    2665: T208 = 1'h0;
    2666: T208 = 1'h0;
    2667: T208 = 1'h0;
    2668: T208 = 1'h0;
    2669: T208 = 1'h0;
    2670: T208 = 1'h0;
    2671: T208 = 1'h0;
    2672: T208 = 1'h0;
    2673: T208 = 1'h0;
    2674: T208 = 1'h0;
    2675: T208 = 1'h0;
    2676: T208 = 1'h0;
    2677: T208 = 1'h0;
    2678: T208 = 1'h0;
    2679: T208 = 1'h0;
    2680: T208 = 1'h0;
    2681: T208 = 1'h0;
    2682: T208 = 1'h0;
    2683: T208 = 1'h0;
    2684: T208 = 1'h0;
    2685: T208 = 1'h0;
    2686: T208 = 1'h0;
    2687: T208 = 1'h0;
    2688: T208 = 1'h0;
    2689: T208 = 1'h0;
    2690: T208 = 1'h0;
    2691: T208 = 1'h0;
    2692: T208 = 1'h0;
    2693: T208 = 1'h0;
    2694: T208 = 1'h0;
    2695: T208 = 1'h0;
    2696: T208 = 1'h0;
    2697: T208 = 1'h0;
    2698: T208 = 1'h0;
    2699: T208 = 1'h0;
    2700: T208 = 1'h0;
    2701: T208 = 1'h0;
    2702: T208 = 1'h0;
    2703: T208 = 1'h0;
    2704: T208 = 1'h0;
    2705: T208 = 1'h0;
    2706: T208 = 1'h0;
    2707: T208 = 1'h0;
    2708: T208 = 1'h0;
    2709: T208 = 1'h0;
    2710: T208 = 1'h0;
    2711: T208 = 1'h0;
    2712: T208 = 1'h0;
    2713: T208 = 1'h0;
    2714: T208 = 1'h0;
    2715: T208 = 1'h0;
    2716: T208 = 1'h0;
    2717: T208 = 1'h0;
    2718: T208 = 1'h0;
    2719: T208 = 1'h0;
    2720: T208 = 1'h0;
    2721: T208 = 1'h0;
    2722: T208 = 1'h0;
    2723: T208 = 1'h0;
    2724: T208 = 1'h0;
    2725: T208 = 1'h0;
    2726: T208 = 1'h0;
    2727: T208 = 1'h0;
    2728: T208 = 1'h0;
    2729: T208 = 1'h0;
    2730: T208 = 1'h0;
    2731: T208 = 1'h0;
    2732: T208 = 1'h0;
    2733: T208 = 1'h0;
    2734: T208 = 1'h0;
    2735: T208 = 1'h0;
    2736: T208 = 1'h0;
    2737: T208 = 1'h0;
    2738: T208 = 1'h0;
    2739: T208 = 1'h0;
    2740: T208 = 1'h0;
    2741: T208 = 1'h0;
    2742: T208 = 1'h0;
    2743: T208 = 1'h0;
    2744: T208 = 1'h0;
    2745: T208 = 1'h0;
    2746: T208 = 1'h0;
    2747: T208 = 1'h0;
    2748: T208 = 1'h0;
    2749: T208 = 1'h0;
    2750: T208 = 1'h0;
    2751: T208 = 1'h0;
    2752: T208 = 1'h0;
    2753: T208 = 1'h0;
    2754: T208 = 1'h0;
    2755: T208 = 1'h0;
    2756: T208 = 1'h0;
    2757: T208 = 1'h0;
    2758: T208 = 1'h0;
    2759: T208 = 1'h0;
    2760: T208 = 1'h0;
    2761: T208 = 1'h0;
    2762: T208 = 1'h0;
    2763: T208 = 1'h0;
    2764: T208 = 1'h0;
    2765: T208 = 1'h0;
    2766: T208 = 1'h0;
    2767: T208 = 1'h0;
    2768: T208 = 1'h0;
    2769: T208 = 1'h0;
    2770: T208 = 1'h0;
    2771: T208 = 1'h0;
    2772: T208 = 1'h0;
    2773: T208 = 1'h0;
    2774: T208 = 1'h0;
    2775: T208 = 1'h0;
    2776: T208 = 1'h0;
    2777: T208 = 1'h0;
    2778: T208 = 1'h0;
    2779: T208 = 1'h0;
    2780: T208 = 1'h0;
    2781: T208 = 1'h0;
    2782: T208 = 1'h0;
    2783: T208 = 1'h0;
    2784: T208 = 1'h0;
    2785: T208 = 1'h0;
    2786: T208 = 1'h0;
    2787: T208 = 1'h0;
    2788: T208 = 1'h0;
    2789: T208 = 1'h0;
    2790: T208 = 1'h0;
    2791: T208 = 1'h0;
    2792: T208 = 1'h0;
    2793: T208 = 1'h0;
    2794: T208 = 1'h0;
    2795: T208 = 1'h0;
    2796: T208 = 1'h0;
    2797: T208 = 1'h0;
    2798: T208 = 1'h0;
    2799: T208 = 1'h0;
    2800: T208 = 1'h0;
    2801: T208 = 1'h0;
    2802: T208 = 1'h0;
    2803: T208 = 1'h0;
    2804: T208 = 1'h0;
    2805: T208 = 1'h0;
    2806: T208 = 1'h0;
    2807: T208 = 1'h0;
    2808: T208 = 1'h0;
    2809: T208 = 1'h0;
    2810: T208 = 1'h0;
    2811: T208 = 1'h0;
    2812: T208 = 1'h0;
    2813: T208 = 1'h0;
    2814: T208 = 1'h0;
    2815: T208 = 1'h0;
    2816: T208 = 1'h0;
    2817: T208 = 1'h0;
    2818: T208 = 1'h0;
    2819: T208 = 1'h0;
    2820: T208 = 1'h0;
    2821: T208 = 1'h0;
    2822: T208 = 1'h0;
    2823: T208 = 1'h0;
    2824: T208 = 1'h0;
    2825: T208 = 1'h0;
    2826: T208 = 1'h0;
    2827: T208 = 1'h0;
    2828: T208 = 1'h0;
    2829: T208 = 1'h0;
    2830: T208 = 1'h0;
    2831: T208 = 1'h0;
    2832: T208 = 1'h0;
    2833: T208 = 1'h0;
    2834: T208 = 1'h0;
    2835: T208 = 1'h0;
    2836: T208 = 1'h0;
    2837: T208 = 1'h0;
    2838: T208 = 1'h0;
    2839: T208 = 1'h0;
    2840: T208 = 1'h0;
    2841: T208 = 1'h0;
    2842: T208 = 1'h0;
    2843: T208 = 1'h0;
    2844: T208 = 1'h0;
    2845: T208 = 1'h0;
    2846: T208 = 1'h0;
    2847: T208 = 1'h0;
    2848: T208 = 1'h0;
    2849: T208 = 1'h0;
    2850: T208 = 1'h0;
    2851: T208 = 1'h0;
    2852: T208 = 1'h0;
    2853: T208 = 1'h0;
    2854: T208 = 1'h0;
    2855: T208 = 1'h0;
    2856: T208 = 1'h0;
    2857: T208 = 1'h0;
    2858: T208 = 1'h0;
    2859: T208 = 1'h0;
    2860: T208 = 1'h0;
    2861: T208 = 1'h0;
    2862: T208 = 1'h0;
    2863: T208 = 1'h0;
    2864: T208 = 1'h0;
    2865: T208 = 1'h0;
    2866: T208 = 1'h0;
    2867: T208 = 1'h0;
    2868: T208 = 1'h0;
    2869: T208 = 1'h0;
    2870: T208 = 1'h0;
    2871: T208 = 1'h0;
    2872: T208 = 1'h0;
    2873: T208 = 1'h0;
    2874: T208 = 1'h0;
    2875: T208 = 1'h0;
    2876: T208 = 1'h0;
    2877: T208 = 1'h0;
    2878: T208 = 1'h0;
    2879: T208 = 1'h0;
    2880: T208 = 1'h0;
    2881: T208 = 1'h0;
    2882: T208 = 1'h0;
    2883: T208 = 1'h0;
    2884: T208 = 1'h0;
    2885: T208 = 1'h0;
    2886: T208 = 1'h0;
    2887: T208 = 1'h0;
    2888: T208 = 1'h0;
    2889: T208 = 1'h0;
    2890: T208 = 1'h0;
    2891: T208 = 1'h0;
    2892: T208 = 1'h0;
    2893: T208 = 1'h0;
    2894: T208 = 1'h0;
    2895: T208 = 1'h0;
    2896: T208 = 1'h0;
    2897: T208 = 1'h0;
    2898: T208 = 1'h0;
    2899: T208 = 1'h0;
    2900: T208 = 1'h0;
    2901: T208 = 1'h0;
    2902: T208 = 1'h0;
    2903: T208 = 1'h0;
    2904: T208 = 1'h0;
    2905: T208 = 1'h0;
    2906: T208 = 1'h0;
    2907: T208 = 1'h0;
    2908: T208 = 1'h0;
    2909: T208 = 1'h0;
    2910: T208 = 1'h0;
    2911: T208 = 1'h0;
    2912: T208 = 1'h0;
    2913: T208 = 1'h0;
    2914: T208 = 1'h0;
    2915: T208 = 1'h0;
    2916: T208 = 1'h0;
    2917: T208 = 1'h0;
    2918: T208 = 1'h0;
    2919: T208 = 1'h0;
    2920: T208 = 1'h0;
    2921: T208 = 1'h0;
    2922: T208 = 1'h0;
    2923: T208 = 1'h0;
    2924: T208 = 1'h0;
    2925: T208 = 1'h0;
    2926: T208 = 1'h0;
    2927: T208 = 1'h0;
    2928: T208 = 1'h0;
    2929: T208 = 1'h0;
    2930: T208 = 1'h0;
    2931: T208 = 1'h0;
    2932: T208 = 1'h0;
    2933: T208 = 1'h0;
    2934: T208 = 1'h0;
    2935: T208 = 1'h0;
    2936: T208 = 1'h0;
    2937: T208 = 1'h0;
    2938: T208 = 1'h0;
    2939: T208 = 1'h0;
    2940: T208 = 1'h0;
    2941: T208 = 1'h0;
    2942: T208 = 1'h0;
    2943: T208 = 1'h0;
    2944: T208 = 1'h0;
    2945: T208 = 1'h0;
    2946: T208 = 1'h0;
    2947: T208 = 1'h0;
    2948: T208 = 1'h0;
    2949: T208 = 1'h0;
    2950: T208 = 1'h0;
    2951: T208 = 1'h0;
    2952: T208 = 1'h0;
    2953: T208 = 1'h0;
    2954: T208 = 1'h0;
    2955: T208 = 1'h0;
    2956: T208 = 1'h0;
    2957: T208 = 1'h0;
    2958: T208 = 1'h0;
    2959: T208 = 1'h0;
    2960: T208 = 1'h0;
    2961: T208 = 1'h0;
    2962: T208 = 1'h0;
    2963: T208 = 1'h0;
    2964: T208 = 1'h0;
    2965: T208 = 1'h0;
    2966: T208 = 1'h0;
    2967: T208 = 1'h0;
    2968: T208 = 1'h0;
    2969: T208 = 1'h0;
    2970: T208 = 1'h0;
    2971: T208 = 1'h0;
    2972: T208 = 1'h0;
    2973: T208 = 1'h0;
    2974: T208 = 1'h0;
    2975: T208 = 1'h0;
    2976: T208 = 1'h0;
    2977: T208 = 1'h0;
    2978: T208 = 1'h0;
    2979: T208 = 1'h0;
    2980: T208 = 1'h0;
    2981: T208 = 1'h0;
    2982: T208 = 1'h0;
    2983: T208 = 1'h0;
    2984: T208 = 1'h0;
    2985: T208 = 1'h0;
    2986: T208 = 1'h0;
    2987: T208 = 1'h0;
    2988: T208 = 1'h0;
    2989: T208 = 1'h0;
    2990: T208 = 1'h0;
    2991: T208 = 1'h0;
    2992: T208 = 1'h0;
    2993: T208 = 1'h0;
    2994: T208 = 1'h0;
    2995: T208 = 1'h0;
    2996: T208 = 1'h0;
    2997: T208 = 1'h0;
    2998: T208 = 1'h0;
    2999: T208 = 1'h0;
    3000: T208 = 1'h0;
    3001: T208 = 1'h0;
    3002: T208 = 1'h0;
    3003: T208 = 1'h0;
    3004: T208 = 1'h0;
    3005: T208 = 1'h0;
    3006: T208 = 1'h0;
    3007: T208 = 1'h0;
    3008: T208 = 1'h0;
    3009: T208 = 1'h0;
    3010: T208 = 1'h0;
    3011: T208 = 1'h0;
    3012: T208 = 1'h0;
    3013: T208 = 1'h0;
    3014: T208 = 1'h0;
    3015: T208 = 1'h0;
    3016: T208 = 1'h0;
    3017: T208 = 1'h0;
    3018: T208 = 1'h0;
    3019: T208 = 1'h0;
    3020: T208 = 1'h0;
    3021: T208 = 1'h0;
    3022: T208 = 1'h0;
    3023: T208 = 1'h0;
    3024: T208 = 1'h0;
    3025: T208 = 1'h0;
    3026: T208 = 1'h0;
    3027: T208 = 1'h0;
    3028: T208 = 1'h0;
    3029: T208 = 1'h0;
    3030: T208 = 1'h0;
    3031: T208 = 1'h0;
    3032: T208 = 1'h0;
    3033: T208 = 1'h0;
    3034: T208 = 1'h0;
    3035: T208 = 1'h0;
    3036: T208 = 1'h0;
    3037: T208 = 1'h0;
    3038: T208 = 1'h0;
    3039: T208 = 1'h0;
    3040: T208 = 1'h0;
    3041: T208 = 1'h0;
    3042: T208 = 1'h0;
    3043: T208 = 1'h0;
    3044: T208 = 1'h0;
    3045: T208 = 1'h0;
    3046: T208 = 1'h0;
    3047: T208 = 1'h0;
    3048: T208 = 1'h0;
    3049: T208 = 1'h0;
    3050: T208 = 1'h0;
    3051: T208 = 1'h0;
    3052: T208 = 1'h0;
    3053: T208 = 1'h0;
    3054: T208 = 1'h0;
    3055: T208 = 1'h0;
    3056: T208 = 1'h0;
    3057: T208 = 1'h0;
    3058: T208 = 1'h0;
    3059: T208 = 1'h0;
    3060: T208 = 1'h0;
    3061: T208 = 1'h0;
    3062: T208 = 1'h0;
    3063: T208 = 1'h0;
    3064: T208 = 1'h0;
    3065: T208 = 1'h0;
    3066: T208 = 1'h0;
    3067: T208 = 1'h0;
    3068: T208 = 1'h0;
    3069: T208 = 1'h0;
    3070: T208 = 1'h0;
    3071: T208 = 1'h0;
    3072: T208 = 1'h1;
    3073: T208 = 1'h1;
    3074: T208 = 1'h1;
    3075: T208 = 1'h0;
    3076: T208 = 1'h0;
    3077: T208 = 1'h0;
    3078: T208 = 1'h0;
    3079: T208 = 1'h0;
    3080: T208 = 1'h0;
    3081: T208 = 1'h0;
    3082: T208 = 1'h0;
    3083: T208 = 1'h0;
    3084: T208 = 1'h0;
    3085: T208 = 1'h0;
    3086: T208 = 1'h0;
    3087: T208 = 1'h0;
    3088: T208 = 1'h0;
    3089: T208 = 1'h0;
    3090: T208 = 1'h0;
    3091: T208 = 1'h0;
    3092: T208 = 1'h0;
    3093: T208 = 1'h0;
    3094: T208 = 1'h0;
    3095: T208 = 1'h0;
    3096: T208 = 1'h0;
    3097: T208 = 1'h0;
    3098: T208 = 1'h0;
    3099: T208 = 1'h0;
    3100: T208 = 1'h0;
    3101: T208 = 1'h0;
    3102: T208 = 1'h0;
    3103: T208 = 1'h0;
    3104: T208 = 1'h0;
    3105: T208 = 1'h0;
    3106: T208 = 1'h0;
    3107: T208 = 1'h0;
    3108: T208 = 1'h0;
    3109: T208 = 1'h0;
    3110: T208 = 1'h0;
    3111: T208 = 1'h0;
    3112: T208 = 1'h0;
    3113: T208 = 1'h0;
    3114: T208 = 1'h0;
    3115: T208 = 1'h0;
    3116: T208 = 1'h0;
    3117: T208 = 1'h0;
    3118: T208 = 1'h0;
    3119: T208 = 1'h0;
    3120: T208 = 1'h0;
    3121: T208 = 1'h0;
    3122: T208 = 1'h0;
    3123: T208 = 1'h0;
    3124: T208 = 1'h0;
    3125: T208 = 1'h0;
    3126: T208 = 1'h0;
    3127: T208 = 1'h0;
    3128: T208 = 1'h0;
    3129: T208 = 1'h0;
    3130: T208 = 1'h0;
    3131: T208 = 1'h0;
    3132: T208 = 1'h0;
    3133: T208 = 1'h0;
    3134: T208 = 1'h0;
    3135: T208 = 1'h0;
    3136: T208 = 1'h0;
    3137: T208 = 1'h0;
    3138: T208 = 1'h0;
    3139: T208 = 1'h0;
    3140: T208 = 1'h0;
    3141: T208 = 1'h0;
    3142: T208 = 1'h0;
    3143: T208 = 1'h0;
    3144: T208 = 1'h0;
    3145: T208 = 1'h0;
    3146: T208 = 1'h0;
    3147: T208 = 1'h0;
    3148: T208 = 1'h0;
    3149: T208 = 1'h0;
    3150: T208 = 1'h0;
    3151: T208 = 1'h0;
    3152: T208 = 1'h0;
    3153: T208 = 1'h0;
    3154: T208 = 1'h0;
    3155: T208 = 1'h0;
    3156: T208 = 1'h0;
    3157: T208 = 1'h0;
    3158: T208 = 1'h0;
    3159: T208 = 1'h0;
    3160: T208 = 1'h0;
    3161: T208 = 1'h0;
    3162: T208 = 1'h0;
    3163: T208 = 1'h0;
    3164: T208 = 1'h0;
    3165: T208 = 1'h0;
    3166: T208 = 1'h0;
    3167: T208 = 1'h0;
    3168: T208 = 1'h0;
    3169: T208 = 1'h0;
    3170: T208 = 1'h0;
    3171: T208 = 1'h0;
    3172: T208 = 1'h0;
    3173: T208 = 1'h0;
    3174: T208 = 1'h0;
    3175: T208 = 1'h0;
    3176: T208 = 1'h0;
    3177: T208 = 1'h0;
    3178: T208 = 1'h0;
    3179: T208 = 1'h0;
    3180: T208 = 1'h0;
    3181: T208 = 1'h0;
    3182: T208 = 1'h0;
    3183: T208 = 1'h0;
    3184: T208 = 1'h0;
    3185: T208 = 1'h0;
    3186: T208 = 1'h0;
    3187: T208 = 1'h0;
    3188: T208 = 1'h0;
    3189: T208 = 1'h0;
    3190: T208 = 1'h0;
    3191: T208 = 1'h0;
    3192: T208 = 1'h0;
    3193: T208 = 1'h0;
    3194: T208 = 1'h0;
    3195: T208 = 1'h0;
    3196: T208 = 1'h0;
    3197: T208 = 1'h0;
    3198: T208 = 1'h0;
    3199: T208 = 1'h0;
    3200: T208 = 1'h0;
    3201: T208 = 1'h0;
    3202: T208 = 1'h0;
    3203: T208 = 1'h0;
    3204: T208 = 1'h0;
    3205: T208 = 1'h0;
    3206: T208 = 1'h0;
    3207: T208 = 1'h0;
    3208: T208 = 1'h0;
    3209: T208 = 1'h0;
    3210: T208 = 1'h0;
    3211: T208 = 1'h0;
    3212: T208 = 1'h0;
    3213: T208 = 1'h0;
    3214: T208 = 1'h0;
    3215: T208 = 1'h0;
    3216: T208 = 1'h0;
    3217: T208 = 1'h0;
    3218: T208 = 1'h0;
    3219: T208 = 1'h0;
    3220: T208 = 1'h0;
    3221: T208 = 1'h0;
    3222: T208 = 1'h0;
    3223: T208 = 1'h0;
    3224: T208 = 1'h0;
    3225: T208 = 1'h0;
    3226: T208 = 1'h0;
    3227: T208 = 1'h0;
    3228: T208 = 1'h0;
    3229: T208 = 1'h0;
    3230: T208 = 1'h0;
    3231: T208 = 1'h0;
    3232: T208 = 1'h0;
    3233: T208 = 1'h0;
    3234: T208 = 1'h0;
    3235: T208 = 1'h0;
    3236: T208 = 1'h0;
    3237: T208 = 1'h0;
    3238: T208 = 1'h0;
    3239: T208 = 1'h0;
    3240: T208 = 1'h0;
    3241: T208 = 1'h0;
    3242: T208 = 1'h0;
    3243: T208 = 1'h0;
    3244: T208 = 1'h0;
    3245: T208 = 1'h0;
    3246: T208 = 1'h0;
    3247: T208 = 1'h0;
    3248: T208 = 1'h0;
    3249: T208 = 1'h0;
    3250: T208 = 1'h0;
    3251: T208 = 1'h0;
    3252: T208 = 1'h0;
    3253: T208 = 1'h0;
    3254: T208 = 1'h0;
    3255: T208 = 1'h0;
    3256: T208 = 1'h0;
    3257: T208 = 1'h0;
    3258: T208 = 1'h0;
    3259: T208 = 1'h0;
    3260: T208 = 1'h0;
    3261: T208 = 1'h0;
    3262: T208 = 1'h0;
    3263: T208 = 1'h0;
    3264: T208 = 1'h1;
    3265: T208 = 1'h1;
    3266: T208 = 1'h1;
    3267: T208 = 1'h1;
    3268: T208 = 1'h1;
    3269: T208 = 1'h1;
    3270: T208 = 1'h1;
    3271: T208 = 1'h1;
    3272: T208 = 1'h1;
    3273: T208 = 1'h1;
    3274: T208 = 1'h1;
    3275: T208 = 1'h1;
    3276: T208 = 1'h1;
    3277: T208 = 1'h1;
    3278: T208 = 1'h1;
    3279: T208 = 1'h1;
    3280: T208 = 1'h0;
    3281: T208 = 1'h0;
    3282: T208 = 1'h0;
    3283: T208 = 1'h0;
    3284: T208 = 1'h0;
    3285: T208 = 1'h0;
    3286: T208 = 1'h0;
    3287: T208 = 1'h0;
    3288: T208 = 1'h0;
    3289: T208 = 1'h0;
    3290: T208 = 1'h0;
    3291: T208 = 1'h0;
    3292: T208 = 1'h0;
    3293: T208 = 1'h0;
    3294: T208 = 1'h0;
    3295: T208 = 1'h0;
    3296: T208 = 1'h0;
    3297: T208 = 1'h0;
    3298: T208 = 1'h0;
    3299: T208 = 1'h0;
    3300: T208 = 1'h0;
    3301: T208 = 1'h0;
    3302: T208 = 1'h0;
    3303: T208 = 1'h0;
    3304: T208 = 1'h0;
    3305: T208 = 1'h0;
    3306: T208 = 1'h0;
    3307: T208 = 1'h0;
    3308: T208 = 1'h0;
    3309: T208 = 1'h0;
    3310: T208 = 1'h0;
    3311: T208 = 1'h0;
    3312: T208 = 1'h0;
    3313: T208 = 1'h0;
    3314: T208 = 1'h0;
    3315: T208 = 1'h0;
    3316: T208 = 1'h0;
    3317: T208 = 1'h0;
    3318: T208 = 1'h0;
    3319: T208 = 1'h0;
    3320: T208 = 1'h0;
    3321: T208 = 1'h0;
    3322: T208 = 1'h0;
    3323: T208 = 1'h0;
    3324: T208 = 1'h0;
    3325: T208 = 1'h0;
    3326: T208 = 1'h0;
    3327: T208 = 1'h0;
    3328: T208 = 1'h0;
    3329: T208 = 1'h0;
    3330: T208 = 1'h0;
    3331: T208 = 1'h0;
    3332: T208 = 1'h0;
    3333: T208 = 1'h0;
    3334: T208 = 1'h0;
    3335: T208 = 1'h0;
    3336: T208 = 1'h0;
    3337: T208 = 1'h0;
    3338: T208 = 1'h0;
    3339: T208 = 1'h0;
    3340: T208 = 1'h0;
    3341: T208 = 1'h0;
    3342: T208 = 1'h0;
    3343: T208 = 1'h0;
    3344: T208 = 1'h0;
    3345: T208 = 1'h0;
    3346: T208 = 1'h0;
    3347: T208 = 1'h0;
    3348: T208 = 1'h0;
    3349: T208 = 1'h0;
    3350: T208 = 1'h0;
    3351: T208 = 1'h0;
    3352: T208 = 1'h0;
    3353: T208 = 1'h0;
    3354: T208 = 1'h0;
    3355: T208 = 1'h0;
    3356: T208 = 1'h0;
    3357: T208 = 1'h0;
    3358: T208 = 1'h0;
    3359: T208 = 1'h0;
    3360: T208 = 1'h0;
    3361: T208 = 1'h0;
    3362: T208 = 1'h0;
    3363: T208 = 1'h0;
    3364: T208 = 1'h0;
    3365: T208 = 1'h0;
    3366: T208 = 1'h0;
    3367: T208 = 1'h0;
    3368: T208 = 1'h0;
    3369: T208 = 1'h0;
    3370: T208 = 1'h0;
    3371: T208 = 1'h0;
    3372: T208 = 1'h0;
    3373: T208 = 1'h0;
    3374: T208 = 1'h0;
    3375: T208 = 1'h0;
    3376: T208 = 1'h0;
    3377: T208 = 1'h0;
    3378: T208 = 1'h0;
    3379: T208 = 1'h0;
    3380: T208 = 1'h0;
    3381: T208 = 1'h0;
    3382: T208 = 1'h0;
    3383: T208 = 1'h0;
    3384: T208 = 1'h0;
    3385: T208 = 1'h0;
    3386: T208 = 1'h0;
    3387: T208 = 1'h0;
    3388: T208 = 1'h0;
    3389: T208 = 1'h0;
    3390: T208 = 1'h0;
    3391: T208 = 1'h0;
    3392: T208 = 1'h0;
    3393: T208 = 1'h0;
    3394: T208 = 1'h0;
    3395: T208 = 1'h0;
    3396: T208 = 1'h0;
    3397: T208 = 1'h0;
    3398: T208 = 1'h0;
    3399: T208 = 1'h0;
    3400: T208 = 1'h0;
    3401: T208 = 1'h0;
    3402: T208 = 1'h0;
    3403: T208 = 1'h0;
    3404: T208 = 1'h0;
    3405: T208 = 1'h0;
    3406: T208 = 1'h0;
    3407: T208 = 1'h0;
    3408: T208 = 1'h0;
    3409: T208 = 1'h0;
    3410: T208 = 1'h0;
    3411: T208 = 1'h0;
    3412: T208 = 1'h0;
    3413: T208 = 1'h0;
    3414: T208 = 1'h0;
    3415: T208 = 1'h0;
    3416: T208 = 1'h0;
    3417: T208 = 1'h0;
    3418: T208 = 1'h0;
    3419: T208 = 1'h0;
    3420: T208 = 1'h0;
    3421: T208 = 1'h0;
    3422: T208 = 1'h0;
    3423: T208 = 1'h0;
    3424: T208 = 1'h0;
    3425: T208 = 1'h0;
    3426: T208 = 1'h0;
    3427: T208 = 1'h0;
    3428: T208 = 1'h0;
    3429: T208 = 1'h0;
    3430: T208 = 1'h0;
    3431: T208 = 1'h0;
    3432: T208 = 1'h0;
    3433: T208 = 1'h0;
    3434: T208 = 1'h0;
    3435: T208 = 1'h0;
    3436: T208 = 1'h0;
    3437: T208 = 1'h0;
    3438: T208 = 1'h0;
    3439: T208 = 1'h0;
    3440: T208 = 1'h0;
    3441: T208 = 1'h0;
    3442: T208 = 1'h0;
    3443: T208 = 1'h0;
    3444: T208 = 1'h0;
    3445: T208 = 1'h0;
    3446: T208 = 1'h0;
    3447: T208 = 1'h0;
    3448: T208 = 1'h0;
    3449: T208 = 1'h0;
    3450: T208 = 1'h0;
    3451: T208 = 1'h0;
    3452: T208 = 1'h0;
    3453: T208 = 1'h0;
    3454: T208 = 1'h0;
    3455: T208 = 1'h0;
    3456: T208 = 1'h0;
    3457: T208 = 1'h0;
    3458: T208 = 1'h0;
    3459: T208 = 1'h0;
    3460: T208 = 1'h0;
    3461: T208 = 1'h0;
    3462: T208 = 1'h0;
    3463: T208 = 1'h0;
    3464: T208 = 1'h0;
    3465: T208 = 1'h0;
    3466: T208 = 1'h0;
    3467: T208 = 1'h0;
    3468: T208 = 1'h0;
    3469: T208 = 1'h0;
    3470: T208 = 1'h0;
    3471: T208 = 1'h0;
    3472: T208 = 1'h0;
    3473: T208 = 1'h0;
    3474: T208 = 1'h0;
    3475: T208 = 1'h0;
    3476: T208 = 1'h0;
    3477: T208 = 1'h0;
    3478: T208 = 1'h0;
    3479: T208 = 1'h0;
    3480: T208 = 1'h0;
    3481: T208 = 1'h0;
    3482: T208 = 1'h0;
    3483: T208 = 1'h0;
    3484: T208 = 1'h0;
    3485: T208 = 1'h0;
    3486: T208 = 1'h0;
    3487: T208 = 1'h0;
    3488: T208 = 1'h0;
    3489: T208 = 1'h0;
    3490: T208 = 1'h0;
    3491: T208 = 1'h0;
    3492: T208 = 1'h0;
    3493: T208 = 1'h0;
    3494: T208 = 1'h0;
    3495: T208 = 1'h0;
    3496: T208 = 1'h0;
    3497: T208 = 1'h0;
    3498: T208 = 1'h0;
    3499: T208 = 1'h0;
    3500: T208 = 1'h0;
    3501: T208 = 1'h0;
    3502: T208 = 1'h0;
    3503: T208 = 1'h0;
    3504: T208 = 1'h0;
    3505: T208 = 1'h0;
    3506: T208 = 1'h0;
    3507: T208 = 1'h0;
    3508: T208 = 1'h0;
    3509: T208 = 1'h0;
    3510: T208 = 1'h0;
    3511: T208 = 1'h0;
    3512: T208 = 1'h0;
    3513: T208 = 1'h0;
    3514: T208 = 1'h0;
    3515: T208 = 1'h0;
    3516: T208 = 1'h0;
    3517: T208 = 1'h0;
    3518: T208 = 1'h0;
    3519: T208 = 1'h0;
    3520: T208 = 1'h0;
    3521: T208 = 1'h0;
    3522: T208 = 1'h0;
    3523: T208 = 1'h0;
    3524: T208 = 1'h0;
    3525: T208 = 1'h0;
    3526: T208 = 1'h0;
    3527: T208 = 1'h0;
    3528: T208 = 1'h0;
    3529: T208 = 1'h0;
    3530: T208 = 1'h0;
    3531: T208 = 1'h0;
    3532: T208 = 1'h0;
    3533: T208 = 1'h0;
    3534: T208 = 1'h0;
    3535: T208 = 1'h0;
    3536: T208 = 1'h0;
    3537: T208 = 1'h0;
    3538: T208 = 1'h0;
    3539: T208 = 1'h0;
    3540: T208 = 1'h0;
    3541: T208 = 1'h0;
    3542: T208 = 1'h0;
    3543: T208 = 1'h0;
    3544: T208 = 1'h0;
    3545: T208 = 1'h0;
    3546: T208 = 1'h0;
    3547: T208 = 1'h0;
    3548: T208 = 1'h0;
    3549: T208 = 1'h0;
    3550: T208 = 1'h0;
    3551: T208 = 1'h0;
    3552: T208 = 1'h0;
    3553: T208 = 1'h0;
    3554: T208 = 1'h0;
    3555: T208 = 1'h0;
    3556: T208 = 1'h0;
    3557: T208 = 1'h0;
    3558: T208 = 1'h0;
    3559: T208 = 1'h0;
    3560: T208 = 1'h0;
    3561: T208 = 1'h0;
    3562: T208 = 1'h0;
    3563: T208 = 1'h0;
    3564: T208 = 1'h0;
    3565: T208 = 1'h0;
    3566: T208 = 1'h0;
    3567: T208 = 1'h0;
    3568: T208 = 1'h0;
    3569: T208 = 1'h0;
    3570: T208 = 1'h0;
    3571: T208 = 1'h0;
    3572: T208 = 1'h0;
    3573: T208 = 1'h0;
    3574: T208 = 1'h0;
    3575: T208 = 1'h0;
    3576: T208 = 1'h0;
    3577: T208 = 1'h0;
    3578: T208 = 1'h0;
    3579: T208 = 1'h0;
    3580: T208 = 1'h0;
    3581: T208 = 1'h0;
    3582: T208 = 1'h0;
    3583: T208 = 1'h0;
    3584: T208 = 1'h0;
    3585: T208 = 1'h0;
    3586: T208 = 1'h0;
    3587: T208 = 1'h0;
    3588: T208 = 1'h0;
    3589: T208 = 1'h0;
    3590: T208 = 1'h0;
    3591: T208 = 1'h0;
    3592: T208 = 1'h0;
    3593: T208 = 1'h0;
    3594: T208 = 1'h0;
    3595: T208 = 1'h0;
    3596: T208 = 1'h0;
    3597: T208 = 1'h0;
    3598: T208 = 1'h0;
    3599: T208 = 1'h0;
    3600: T208 = 1'h0;
    3601: T208 = 1'h0;
    3602: T208 = 1'h0;
    3603: T208 = 1'h0;
    3604: T208 = 1'h0;
    3605: T208 = 1'h0;
    3606: T208 = 1'h0;
    3607: T208 = 1'h0;
    3608: T208 = 1'h0;
    3609: T208 = 1'h0;
    3610: T208 = 1'h0;
    3611: T208 = 1'h0;
    3612: T208 = 1'h0;
    3613: T208 = 1'h0;
    3614: T208 = 1'h0;
    3615: T208 = 1'h0;
    3616: T208 = 1'h0;
    3617: T208 = 1'h0;
    3618: T208 = 1'h0;
    3619: T208 = 1'h0;
    3620: T208 = 1'h0;
    3621: T208 = 1'h0;
    3622: T208 = 1'h0;
    3623: T208 = 1'h0;
    3624: T208 = 1'h0;
    3625: T208 = 1'h0;
    3626: T208 = 1'h0;
    3627: T208 = 1'h0;
    3628: T208 = 1'h0;
    3629: T208 = 1'h0;
    3630: T208 = 1'h0;
    3631: T208 = 1'h0;
    3632: T208 = 1'h0;
    3633: T208 = 1'h0;
    3634: T208 = 1'h0;
    3635: T208 = 1'h0;
    3636: T208 = 1'h0;
    3637: T208 = 1'h0;
    3638: T208 = 1'h0;
    3639: T208 = 1'h0;
    3640: T208 = 1'h0;
    3641: T208 = 1'h0;
    3642: T208 = 1'h0;
    3643: T208 = 1'h0;
    3644: T208 = 1'h0;
    3645: T208 = 1'h0;
    3646: T208 = 1'h0;
    3647: T208 = 1'h0;
    3648: T208 = 1'h0;
    3649: T208 = 1'h0;
    3650: T208 = 1'h0;
    3651: T208 = 1'h0;
    3652: T208 = 1'h0;
    3653: T208 = 1'h0;
    3654: T208 = 1'h0;
    3655: T208 = 1'h0;
    3656: T208 = 1'h0;
    3657: T208 = 1'h0;
    3658: T208 = 1'h0;
    3659: T208 = 1'h0;
    3660: T208 = 1'h0;
    3661: T208 = 1'h0;
    3662: T208 = 1'h0;
    3663: T208 = 1'h0;
    3664: T208 = 1'h0;
    3665: T208 = 1'h0;
    3666: T208 = 1'h0;
    3667: T208 = 1'h0;
    3668: T208 = 1'h0;
    3669: T208 = 1'h0;
    3670: T208 = 1'h0;
    3671: T208 = 1'h0;
    3672: T208 = 1'h0;
    3673: T208 = 1'h0;
    3674: T208 = 1'h0;
    3675: T208 = 1'h0;
    3676: T208 = 1'h0;
    3677: T208 = 1'h0;
    3678: T208 = 1'h0;
    3679: T208 = 1'h0;
    3680: T208 = 1'h0;
    3681: T208 = 1'h0;
    3682: T208 = 1'h0;
    3683: T208 = 1'h0;
    3684: T208 = 1'h0;
    3685: T208 = 1'h0;
    3686: T208 = 1'h0;
    3687: T208 = 1'h0;
    3688: T208 = 1'h0;
    3689: T208 = 1'h0;
    3690: T208 = 1'h0;
    3691: T208 = 1'h0;
    3692: T208 = 1'h0;
    3693: T208 = 1'h0;
    3694: T208 = 1'h0;
    3695: T208 = 1'h0;
    3696: T208 = 1'h0;
    3697: T208 = 1'h0;
    3698: T208 = 1'h0;
    3699: T208 = 1'h0;
    3700: T208 = 1'h0;
    3701: T208 = 1'h0;
    3702: T208 = 1'h0;
    3703: T208 = 1'h0;
    3704: T208 = 1'h0;
    3705: T208 = 1'h0;
    3706: T208 = 1'h0;
    3707: T208 = 1'h0;
    3708: T208 = 1'h0;
    3709: T208 = 1'h0;
    3710: T208 = 1'h0;
    3711: T208 = 1'h0;
    3712: T208 = 1'h0;
    3713: T208 = 1'h0;
    3714: T208 = 1'h0;
    3715: T208 = 1'h0;
    3716: T208 = 1'h0;
    3717: T208 = 1'h0;
    3718: T208 = 1'h0;
    3719: T208 = 1'h0;
    3720: T208 = 1'h0;
    3721: T208 = 1'h0;
    3722: T208 = 1'h0;
    3723: T208 = 1'h0;
    3724: T208 = 1'h0;
    3725: T208 = 1'h0;
    3726: T208 = 1'h0;
    3727: T208 = 1'h0;
    3728: T208 = 1'h0;
    3729: T208 = 1'h0;
    3730: T208 = 1'h0;
    3731: T208 = 1'h0;
    3732: T208 = 1'h0;
    3733: T208 = 1'h0;
    3734: T208 = 1'h0;
    3735: T208 = 1'h0;
    3736: T208 = 1'h0;
    3737: T208 = 1'h0;
    3738: T208 = 1'h0;
    3739: T208 = 1'h0;
    3740: T208 = 1'h0;
    3741: T208 = 1'h0;
    3742: T208 = 1'h0;
    3743: T208 = 1'h0;
    3744: T208 = 1'h0;
    3745: T208 = 1'h0;
    3746: T208 = 1'h0;
    3747: T208 = 1'h0;
    3748: T208 = 1'h0;
    3749: T208 = 1'h0;
    3750: T208 = 1'h0;
    3751: T208 = 1'h0;
    3752: T208 = 1'h0;
    3753: T208 = 1'h0;
    3754: T208 = 1'h0;
    3755: T208 = 1'h0;
    3756: T208 = 1'h0;
    3757: T208 = 1'h0;
    3758: T208 = 1'h0;
    3759: T208 = 1'h0;
    3760: T208 = 1'h0;
    3761: T208 = 1'h0;
    3762: T208 = 1'h0;
    3763: T208 = 1'h0;
    3764: T208 = 1'h0;
    3765: T208 = 1'h0;
    3766: T208 = 1'h0;
    3767: T208 = 1'h0;
    3768: T208 = 1'h0;
    3769: T208 = 1'h0;
    3770: T208 = 1'h0;
    3771: T208 = 1'h0;
    3772: T208 = 1'h0;
    3773: T208 = 1'h0;
    3774: T208 = 1'h0;
    3775: T208 = 1'h0;
    3776: T208 = 1'h0;
    3777: T208 = 1'h0;
    3778: T208 = 1'h0;
    3779: T208 = 1'h0;
    3780: T208 = 1'h0;
    3781: T208 = 1'h0;
    3782: T208 = 1'h0;
    3783: T208 = 1'h0;
    3784: T208 = 1'h0;
    3785: T208 = 1'h0;
    3786: T208 = 1'h0;
    3787: T208 = 1'h0;
    3788: T208 = 1'h0;
    3789: T208 = 1'h0;
    3790: T208 = 1'h0;
    3791: T208 = 1'h0;
    3792: T208 = 1'h0;
    3793: T208 = 1'h0;
    3794: T208 = 1'h0;
    3795: T208 = 1'h0;
    3796: T208 = 1'h0;
    3797: T208 = 1'h0;
    3798: T208 = 1'h0;
    3799: T208 = 1'h0;
    3800: T208 = 1'h0;
    3801: T208 = 1'h0;
    3802: T208 = 1'h0;
    3803: T208 = 1'h0;
    3804: T208 = 1'h0;
    3805: T208 = 1'h0;
    3806: T208 = 1'h0;
    3807: T208 = 1'h0;
    3808: T208 = 1'h0;
    3809: T208 = 1'h0;
    3810: T208 = 1'h0;
    3811: T208 = 1'h0;
    3812: T208 = 1'h0;
    3813: T208 = 1'h0;
    3814: T208 = 1'h0;
    3815: T208 = 1'h0;
    3816: T208 = 1'h0;
    3817: T208 = 1'h0;
    3818: T208 = 1'h0;
    3819: T208 = 1'h0;
    3820: T208 = 1'h0;
    3821: T208 = 1'h0;
    3822: T208 = 1'h0;
    3823: T208 = 1'h0;
    3824: T208 = 1'h0;
    3825: T208 = 1'h0;
    3826: T208 = 1'h0;
    3827: T208 = 1'h0;
    3828: T208 = 1'h0;
    3829: T208 = 1'h0;
    3830: T208 = 1'h0;
    3831: T208 = 1'h0;
    3832: T208 = 1'h0;
    3833: T208 = 1'h0;
    3834: T208 = 1'h0;
    3835: T208 = 1'h0;
    3836: T208 = 1'h0;
    3837: T208 = 1'h0;
    3838: T208 = 1'h0;
    3839: T208 = 1'h0;
    3840: T208 = 1'h0;
    3841: T208 = 1'h0;
    3842: T208 = 1'h0;
    3843: T208 = 1'h0;
    3844: T208 = 1'h0;
    3845: T208 = 1'h0;
    3846: T208 = 1'h0;
    3847: T208 = 1'h0;
    3848: T208 = 1'h0;
    3849: T208 = 1'h0;
    3850: T208 = 1'h0;
    3851: T208 = 1'h0;
    3852: T208 = 1'h0;
    3853: T208 = 1'h0;
    3854: T208 = 1'h0;
    3855: T208 = 1'h0;
    3856: T208 = 1'h0;
    3857: T208 = 1'h0;
    3858: T208 = 1'h0;
    3859: T208 = 1'h0;
    3860: T208 = 1'h0;
    3861: T208 = 1'h0;
    3862: T208 = 1'h0;
    3863: T208 = 1'h0;
    3864: T208 = 1'h0;
    3865: T208 = 1'h0;
    3866: T208 = 1'h0;
    3867: T208 = 1'h0;
    3868: T208 = 1'h0;
    3869: T208 = 1'h0;
    3870: T208 = 1'h0;
    3871: T208 = 1'h0;
    3872: T208 = 1'h0;
    3873: T208 = 1'h0;
    3874: T208 = 1'h0;
    3875: T208 = 1'h0;
    3876: T208 = 1'h0;
    3877: T208 = 1'h0;
    3878: T208 = 1'h0;
    3879: T208 = 1'h0;
    3880: T208 = 1'h0;
    3881: T208 = 1'h0;
    3882: T208 = 1'h0;
    3883: T208 = 1'h0;
    3884: T208 = 1'h0;
    3885: T208 = 1'h0;
    3886: T208 = 1'h0;
    3887: T208 = 1'h0;
    3888: T208 = 1'h0;
    3889: T208 = 1'h0;
    3890: T208 = 1'h0;
    3891: T208 = 1'h0;
    3892: T208 = 1'h0;
    3893: T208 = 1'h0;
    3894: T208 = 1'h0;
    3895: T208 = 1'h0;
    3896: T208 = 1'h0;
    3897: T208 = 1'h0;
    3898: T208 = 1'h0;
    3899: T208 = 1'h0;
    3900: T208 = 1'h0;
    3901: T208 = 1'h0;
    3902: T208 = 1'h0;
    3903: T208 = 1'h0;
    3904: T208 = 1'h0;
    3905: T208 = 1'h0;
    3906: T208 = 1'h0;
    3907: T208 = 1'h0;
    3908: T208 = 1'h0;
    3909: T208 = 1'h0;
    3910: T208 = 1'h0;
    3911: T208 = 1'h0;
    3912: T208 = 1'h0;
    3913: T208 = 1'h0;
    3914: T208 = 1'h0;
    3915: T208 = 1'h0;
    3916: T208 = 1'h0;
    3917: T208 = 1'h0;
    3918: T208 = 1'h0;
    3919: T208 = 1'h0;
    3920: T208 = 1'h0;
    3921: T208 = 1'h0;
    3922: T208 = 1'h0;
    3923: T208 = 1'h0;
    3924: T208 = 1'h0;
    3925: T208 = 1'h0;
    3926: T208 = 1'h0;
    3927: T208 = 1'h0;
    3928: T208 = 1'h0;
    3929: T208 = 1'h0;
    3930: T208 = 1'h0;
    3931: T208 = 1'h0;
    3932: T208 = 1'h0;
    3933: T208 = 1'h0;
    3934: T208 = 1'h0;
    3935: T208 = 1'h0;
    3936: T208 = 1'h0;
    3937: T208 = 1'h0;
    3938: T208 = 1'h0;
    3939: T208 = 1'h0;
    3940: T208 = 1'h0;
    3941: T208 = 1'h0;
    3942: T208 = 1'h0;
    3943: T208 = 1'h0;
    3944: T208 = 1'h0;
    3945: T208 = 1'h0;
    3946: T208 = 1'h0;
    3947: T208 = 1'h0;
    3948: T208 = 1'h0;
    3949: T208 = 1'h0;
    3950: T208 = 1'h0;
    3951: T208 = 1'h0;
    3952: T208 = 1'h0;
    3953: T208 = 1'h0;
    3954: T208 = 1'h0;
    3955: T208 = 1'h0;
    3956: T208 = 1'h0;
    3957: T208 = 1'h0;
    3958: T208 = 1'h0;
    3959: T208 = 1'h0;
    3960: T208 = 1'h0;
    3961: T208 = 1'h0;
    3962: T208 = 1'h0;
    3963: T208 = 1'h0;
    3964: T208 = 1'h0;
    3965: T208 = 1'h0;
    3966: T208 = 1'h0;
    3967: T208 = 1'h0;
    3968: T208 = 1'h0;
    3969: T208 = 1'h0;
    3970: T208 = 1'h0;
    3971: T208 = 1'h0;
    3972: T208 = 1'h0;
    3973: T208 = 1'h0;
    3974: T208 = 1'h0;
    3975: T208 = 1'h0;
    3976: T208 = 1'h0;
    3977: T208 = 1'h0;
    3978: T208 = 1'h0;
    3979: T208 = 1'h0;
    3980: T208 = 1'h0;
    3981: T208 = 1'h0;
    3982: T208 = 1'h0;
    3983: T208 = 1'h0;
    3984: T208 = 1'h0;
    3985: T208 = 1'h0;
    3986: T208 = 1'h0;
    3987: T208 = 1'h0;
    3988: T208 = 1'h0;
    3989: T208 = 1'h0;
    3990: T208 = 1'h0;
    3991: T208 = 1'h0;
    3992: T208 = 1'h0;
    3993: T208 = 1'h0;
    3994: T208 = 1'h0;
    3995: T208 = 1'h0;
    3996: T208 = 1'h0;
    3997: T208 = 1'h0;
    3998: T208 = 1'h0;
    3999: T208 = 1'h0;
    4000: T208 = 1'h0;
    4001: T208 = 1'h0;
    4002: T208 = 1'h0;
    4003: T208 = 1'h0;
    4004: T208 = 1'h0;
    4005: T208 = 1'h0;
    4006: T208 = 1'h0;
    4007: T208 = 1'h0;
    4008: T208 = 1'h0;
    4009: T208 = 1'h0;
    4010: T208 = 1'h0;
    4011: T208 = 1'h0;
    4012: T208 = 1'h0;
    4013: T208 = 1'h0;
    4014: T208 = 1'h0;
    4015: T208 = 1'h0;
    4016: T208 = 1'h0;
    4017: T208 = 1'h0;
    4018: T208 = 1'h0;
    4019: T208 = 1'h0;
    4020: T208 = 1'h0;
    4021: T208 = 1'h0;
    4022: T208 = 1'h0;
    4023: T208 = 1'h0;
    4024: T208 = 1'h0;
    4025: T208 = 1'h0;
    4026: T208 = 1'h0;
    4027: T208 = 1'h0;
    4028: T208 = 1'h0;
    4029: T208 = 1'h0;
    4030: T208 = 1'h0;
    4031: T208 = 1'h0;
    4032: T208 = 1'h0;
    4033: T208 = 1'h0;
    4034: T208 = 1'h0;
    4035: T208 = 1'h0;
    4036: T208 = 1'h0;
    4037: T208 = 1'h0;
    4038: T208 = 1'h0;
    4039: T208 = 1'h0;
    4040: T208 = 1'h0;
    4041: T208 = 1'h0;
    4042: T208 = 1'h0;
    4043: T208 = 1'h0;
    4044: T208 = 1'h0;
    4045: T208 = 1'h0;
    4046: T208 = 1'h0;
    4047: T208 = 1'h0;
    4048: T208 = 1'h0;
    4049: T208 = 1'h0;
    4050: T208 = 1'h0;
    4051: T208 = 1'h0;
    4052: T208 = 1'h0;
    4053: T208 = 1'h0;
    4054: T208 = 1'h0;
    4055: T208 = 1'h0;
    4056: T208 = 1'h0;
    4057: T208 = 1'h0;
    4058: T208 = 1'h0;
    4059: T208 = 1'h0;
    4060: T208 = 1'h0;
    4061: T208 = 1'h0;
    4062: T208 = 1'h0;
    4063: T208 = 1'h0;
    4064: T208 = 1'h0;
    4065: T208 = 1'h0;
    4066: T208 = 1'h0;
    4067: T208 = 1'h0;
    4068: T208 = 1'h0;
    4069: T208 = 1'h0;
    4070: T208 = 1'h0;
    4071: T208 = 1'h0;
    4072: T208 = 1'h0;
    4073: T208 = 1'h0;
    4074: T208 = 1'h0;
    4075: T208 = 1'h0;
    4076: T208 = 1'h0;
    4077: T208 = 1'h0;
    4078: T208 = 1'h0;
    4079: T208 = 1'h0;
    4080: T208 = 1'h0;
    4081: T208 = 1'h0;
    4082: T208 = 1'h0;
    4083: T208 = 1'h0;
    4084: T208 = 1'h0;
    4085: T208 = 1'h0;
    4086: T208 = 1'h0;
    4087: T208 = 1'h0;
    4088: T208 = 1'h0;
    4089: T208 = 1'h0;
    4090: T208 = 1'h0;
    4091: T208 = 1'h0;
    4092: T208 = 1'h0;
    4093: T208 = 1'h0;
    4094: T208 = 1'h0;
    4095: T208 = 1'h0;
`ifndef SYNTHESIS
    default: T208 = {1{$random}};
`else
    default: T208 = 1'bx;
`endif
  endcase
  assign T210 = T211 ^ 1'h1;
  assign T211 = T214 | T212;
  assign T212 = T213 == 32'h33;
  assign T213 = io_dpath_inst & 32'hfc007077;
  assign T214 = T217 | T215;
  assign T215 = T216 == 32'h4063;
  assign T216 = io_dpath_inst & 32'h407f;
  assign T217 = T220 | T218;
  assign T218 = T219 == 32'h1063;
  assign T219 = io_dpath_inst & 32'h306f;
  assign T220 = T223 | T221;
  assign T221 = T222 == 32'h23;
  assign T222 = io_dpath_inst & 32'h603f;
  assign T223 = T226 | T224;
  assign T224 = T225 == 32'he0000053;
  assign T225 = io_dpath_inst & 32'hedf0707f;
  assign T226 = T229 | T227;
  assign T227 = T228 == 32'he0000053;
  assign T228 = io_dpath_inst & 32'hfdf0607f;
  assign T229 = T232 | T230;
  assign T230 = T231 == 32'hc0000053;
  assign T231 = io_dpath_inst & 32'hedc0007f;
  assign T232 = T235 | T233;
  assign T233 = T234 == 32'h42000053;
  assign T234 = io_dpath_inst & 32'h7ff0007f;
  assign T235 = T238 | T236;
  assign T236 = T237 == 32'h40100053;
  assign T237 = io_dpath_inst & 32'h7ff0007f;
  assign T238 = T241 | T239;
  assign T239 = T240 == 32'h20000053;
  assign T240 = io_dpath_inst & 32'h7c00507f;
  assign T241 = T244 | T242;
  assign T242 = T243 == 32'h20000053;
  assign T243 = io_dpath_inst & 32'h7c00607f;
  assign T244 = T247 | T245;
  assign T245 = T246 == 32'h20000053;
  assign T246 = io_dpath_inst & 32'hf400607f;
  assign T247 = T248 | T69;
  assign T248 = T249 | T72;
  assign T249 = T252 | T250;
  assign T250 = T251 == 32'h2004033;
  assign T251 = io_dpath_inst & 32'hfe004077;
  assign T252 = T255 | T253;
  assign T253 = T254 == 32'h5033;
  assign T254 = io_dpath_inst & 32'hbe007077;
  assign T255 = T258 | T256;
  assign T256 = T257 == 32'h501b;
  assign T257 = io_dpath_inst & 32'hbe00705f;
  assign T258 = T261 | T259;
  assign T259 = T260 == 32'h5013;
  assign T260 = io_dpath_inst & 32'hbc00707f;
  assign T261 = T264 | T262;
  assign T262 = T263 == 32'h2073;
  assign T263 = io_dpath_inst & 32'h207f;
  assign T264 = T265 | T75;
  assign T265 = T268 | T266;
  assign T266 = T267 == 32'h2013;
  assign T267 = io_dpath_inst & 32'h207f;
  assign T268 = T269 | T78;
  assign T269 = T272 | T270;
  assign T270 = T271 == 32'h101b;
  assign T271 = io_dpath_inst & 32'hfe00305f;
  assign T272 = T275 | T273;
  assign T273 = T274 == 32'h1013;
  assign T274 = io_dpath_inst & 32'hfc00305f;
  assign T275 = T278 | T276;
  assign T276 = T277 == 32'h73;
  assign T277 = io_dpath_inst & 32'h7fffffff;
  assign T278 = T281 | T279;
  assign T279 = T280 == 32'h6f;
  assign T280 = io_dpath_inst & 32'h7f;
  assign T281 = T284 | T282;
  assign T282 = T283 == 32'h63;
  assign T283 = io_dpath_inst & 32'h707b;
  assign T284 = T287 | T285;
  assign T285 = T286 == 32'h53;
  assign T286 = io_dpath_inst & 32'hec00007f;
  assign T287 = T290 | T288;
  assign T288 = T289 == 32'h53;
  assign T289 = io_dpath_inst & 32'hf400007f;
  assign T290 = T293 | T291;
  assign T291 = T292 == 32'h43;
  assign T292 = io_dpath_inst & 32'h4000073;
  assign T293 = T296 | T294;
  assign T294 = T295 == 32'h33;
  assign T295 = io_dpath_inst & 32'hbe007077;
  assign T296 = T299 | T297;
  assign T297 = T298 == 32'h33;
  assign T298 = io_dpath_inst & 32'hfc00007f;
  assign T299 = T302 | T300;
  assign T300 = T301 == 32'h17;
  assign T301 = io_dpath_inst & 32'h5f;
  assign T302 = T305 | T303;
  assign T303 = T304 == 32'h13;
  assign T304 = io_dpath_inst & 32'h7077;
  assign T305 = T308 | T306;
  assign T306 = T307 == 32'hf;
  assign T307 = io_dpath_inst & 32'h607f;
  assign T308 = T84 | T309;
  assign T309 = T310 == 32'h3;
  assign T310 = io_dpath_inst & 32'h106f;
  assign T311 = T312 | io_imem_resp_bits_xcpt_if;
  assign T312 = id_interrupt | io_imem_resp_bits_xcpt_ma;
  assign T313 = T314 & io_imem_resp_valid;
  assign T314 = id_interrupt & T315;
  assign T315 = take_pc_mem_wb ^ 1'h1;
  assign T316 = T318 & T317;
  assign T317 = mem_reg_replay_next ^ 1'h1;
  assign T318 = T319 & ex_reg_xcpt_interrupt;
  assign T319 = take_pc_mem_wb ^ 1'h1;
  assign killm_common = T323 | T320;
  assign T320 = mem_reg_valid ^ 1'h1;
  assign T321 = ctrl_killx ? 1'h0 : ex_reg_valid;
  assign T322 = ctrl_killd ? 1'h0 : 1'h1;
  assign T323 = T324 | mem_reg_xcpt;
  assign T324 = dcache_kill_mem | take_pc_wb;
  assign dcache_kill_mem = mem_reg_wen & io_dmem_replay_next_valid;
  assign T325 = ctrl_killx ? 1'h0 : ex_reg_wen;
  assign T326 = ctrl_killd ? 1'h0 : T327;
  assign T327 = T330 | T328;
  assign T328 = T329 == 32'h80000010;
  assign T329 = io_dpath_inst & 32'h90000030;
  assign T330 = T333 | T331;
  assign T331 = T332 == 32'h2030;
  assign T332 = io_dpath_inst & 32'h2030;
  assign T333 = T336 | T334;
  assign T334 = T335 == 32'h1030;
  assign T335 = io_dpath_inst & 32'h1030;
  assign T336 = T339 | T337;
  assign T337 = T338 == 32'h28;
  assign T338 = io_dpath_inst & 32'h28;
  assign T339 = T342 | T340;
  assign T340 = T341 == 32'h24;
  assign T341 = io_dpath_inst & 32'h2024;
  assign T342 = T345 | T343;
  assign T343 = T344 == 32'h10;
  assign T344 = io_dpath_inst & 32'h50;
  assign T345 = T346 == 32'h0;
  assign T346 = io_dpath_inst & 32'h64;
  assign replay_wb_common = T347 | io_dpath_csr_replay;
  assign T347 = io_dmem_resp_bits_nack | wb_reg_replay;
  assign T348 = replay_mem & T349;
  assign T349 = take_pc_wb ^ 1'h1;
  assign replay_mem = T350 | fpu_kill_mem;
  assign T350 = dcache_kill_mem | mem_reg_replay;
  assign T351 = T352 | io_fpu_sboard_set;
  assign T352 = wb_dcache_miss & wb_reg_fp_wen;
  assign T353 = ctrl_killm ? 1'h0 : mem_reg_fp_wen;
  assign T354 = ctrl_killx ? 1'h0 : ex_reg_fp_wen;
  assign T355 = ctrl_killd ? 1'h0 : T356;
  assign T356 = T152 & io_fpu_dec_wen;
  assign wb_dcache_miss = wb_reg_mem_val & T357;
  assign T357 = io_dmem_resp_valid ^ 1'h1;
  assign T358 = ctrl_killm ? 1'h0 : mem_reg_mem_val;
  assign T359 = T123 & T360;
  assign T360 = ~ T361;
  assign T361 = io_dpath_fp_sboard_clr ? T362 : 32'h0;
  assign T362 = 1'h1 << io_dpath_fp_sboard_clra;
  assign T363 = T126 | io_dpath_fp_sboard_clr;
  assign T364 = T359 & T365;
  assign T365 = ~ T366;
  assign T366 = io_fpu_sboard_clr ? T367 : 32'h0;
  assign T367 = 1'h1 << io_fpu_sboard_clra;
  assign T368 = T363 | io_fpu_sboard_clr;
  assign T369 = T378 | T370;
  assign T370 = io_fpu_dec_ren3 & T371;
  assign T371 = T377 & T372;
  assign T372 = T373 - 1'h1;
  assign T373 = 1'h1 << T374;
  assign T374 = T375 + 5'h1;
  assign T375 = T376 - T376;
  assign T376 = io_dpath_inst[5'h1f:5'h1b];
  assign T377 = R118 >> T376;
  assign T378 = T387 | T379;
  assign T379 = io_fpu_dec_ren2 & T380;
  assign T380 = T386 & T381;
  assign T381 = T382 - 1'h1;
  assign T382 = 1'h1 << T383;
  assign T383 = T384 + 5'h1;
  assign T384 = T385 - T385;
  assign T385 = io_dpath_inst[5'h18:5'h14];
  assign T386 = R118 >> T385;
  assign T387 = T395 | T388;
  assign T388 = io_fpu_dec_ren1 & T389;
  assign T389 = T394 & T390;
  assign T390 = T391 - 1'h1;
  assign T391 = 1'h1 << T392;
  assign T392 = T393 + 5'h1;
  assign T393 = T29 - T29;
  assign T394 = R118 >> T29;
  assign T395 = T30 & T396;
  assign T396 = io_fpu_fcsr_rdy ^ 1'h1;
  assign T397 = T470 | id_sboard_hazard;
  assign id_sboard_hazard = T428 | T398;
  assign T398 = id_wen_not0 & T399;
  assign T399 = T404 & T400;
  assign T400 = T401 - 1'h1;
  assign T401 = 1'h1 << T402;
  assign T402 = T403 + 5'h1;
  assign T403 = T116 - T116;
  assign T404 = T405 >> T116;
  assign T405 = R409 & T406;
  assign T406 = ~ T407;
  assign T407 = io_dpath_ll_wen ? T408 : 32'h0;
  assign T408 = 1'h1 << io_dpath_ll_waddr;
  assign T410 = reset ? 32'h0 : T411;
  assign T411 = T426 ? T413 : T412;
  assign T412 = io_dpath_ll_wen ? T405 : R409;
  assign T413 = T405 | T414;
  assign T414 = T416 ? T415 : 32'h0;
  assign T415 = 1'h1 << io_dpath_wb_waddr;
  assign T416 = wb_set_sboard & io_dpath_wb_wen;
  assign wb_set_sboard = T417 | wb_reg_rocc_val;
  assign T417 = wb_reg_div_mul_val | wb_dcache_miss;
  assign T418 = ctrl_killm ? 1'h0 : mem_reg_div_mul_val;
  assign T419 = ex_reg_div_mul_val & io_dpath_div_mul_rdy;
  assign T420 = ctrl_killd ? 1'h0 : T421;
  assign T421 = T424 | T422;
  assign T422 = T423 == 32'h2004020;
  assign T423 = io_dpath_inst & 32'h2004064;
  assign T424 = T425 == 32'h2000030;
  assign T425 = io_dpath_inst & 32'h2004074;
  assign T426 = io_dpath_ll_wen | T416;
  assign id_wen_not0 = T327 & T427;
  assign T427 = T116 != 5'h0;
  assign T428 = T445 | T429;
  assign T429 = id_renx2_not0 & T430;
  assign T430 = T435 & T431;
  assign T431 = T432 - 1'h1;
  assign T432 = 1'h1 << T433;
  assign T433 = T434 + 5'h1;
  assign T434 = T385 - T385;
  assign T435 = T405 >> T385;
  assign id_renx2_not0 = T437 & T436;
  assign T436 = T385 != 5'h0;
  assign T437 = T440 | T438;
  assign T438 = T439 == 32'h2008;
  assign T439 = io_dpath_inst & 32'h2048;
  assign T440 = T443 | T441;
  assign T441 = T442 == 32'h20;
  assign T442 = io_dpath_inst & 32'h34;
  assign T443 = T444 == 32'h20;
  assign T444 = io_dpath_inst & 32'h64;
  assign T445 = id_renx1_not0 & T446;
  assign T446 = T451 & T447;
  assign T447 = T448 - 1'h1;
  assign T448 = 1'h1 << T449;
  assign T449 = T450 + 5'h1;
  assign T450 = T29 - T29;
  assign T451 = T405 >> T29;
  assign id_renx1_not0 = T453 & T452;
  assign T452 = T29 != 5'h0;
  assign T453 = T456 | T454;
  assign T454 = T455 == 32'h90000010;
  assign T455 = io_dpath_inst & 32'h90000034;
  assign T456 = T459 | T457;
  assign T457 = T458 == 32'h2020;
  assign T458 = io_dpath_inst & 32'h6024;
  assign T459 = T462 | T460;
  assign T460 = T461 == 32'h2000;
  assign T461 = io_dpath_inst & 32'h2050;
  assign T462 = T465 | T463;
  assign T463 = T464 == 32'h1020;
  assign T464 = io_dpath_inst & 32'h5024;
  assign T465 = T468 | T466;
  assign T466 = T467 == 32'h20;
  assign T467 = io_dpath_inst & 32'h38;
  assign T468 = T469 == 32'h0;
  assign T469 = io_dpath_inst & 32'h44;
  assign T470 = T495 | id_wb_hazard;
  assign id_wb_hazard = T485 | T471;
  assign T471 = fp_data_hazard_wb & T472;
  assign T472 = wb_dcache_miss | wb_reg_fp_val;
  assign T473 = ctrl_killm ? 1'h0 : mem_reg_fp_val;
  assign fp_data_hazard_wb = wb_reg_fp_wen & T474;
  assign T474 = T477 | T475;
  assign T475 = io_fpu_dec_wen & T476;
  assign T476 = T116 == io_dpath_wb_waddr;
  assign T477 = T480 | T478;
  assign T478 = io_fpu_dec_ren3 & T479;
  assign T479 = T376 == io_dpath_wb_waddr;
  assign T480 = T483 | T481;
  assign T481 = io_fpu_dec_ren2 & T482;
  assign T482 = T385 == io_dpath_wb_waddr;
  assign T483 = io_fpu_dec_ren1 & T484;
  assign T484 = T29 == io_dpath_wb_waddr;
  assign T485 = data_hazard_wb & wb_set_sboard;
  assign data_hazard_wb = wb_reg_wen & T486;
  assign T486 = T489 | T487;
  assign T487 = id_wen_not0 & T488;
  assign T488 = T116 == io_dpath_wb_waddr;
  assign T489 = T492 | T490;
  assign T490 = id_renx2_not0 & T491;
  assign T491 = T385 == io_dpath_wb_waddr;
  assign T492 = id_renx1_not0 & T493;
  assign T493 = T29 == io_dpath_wb_waddr;
  assign T494 = ctrl_killm ? 1'h0 : mem_reg_wen;
  assign T495 = id_ex_hazard | id_mem_hazard;
  assign id_mem_hazard = T508 | T496;
  assign T496 = fp_data_hazard_mem & mem_reg_fp_val;
  assign fp_data_hazard_mem = mem_reg_fp_wen & T497;
  assign T497 = T500 | T498;
  assign T498 = io_fpu_dec_wen & T499;
  assign T499 = T116 == io_dpath_mem_waddr;
  assign T500 = T503 | T501;
  assign T501 = io_fpu_dec_ren3 & T502;
  assign T502 = T376 == io_dpath_mem_waddr;
  assign T503 = T506 | T504;
  assign T504 = io_fpu_dec_ren2 & T505;
  assign T505 = T385 == io_dpath_mem_waddr;
  assign T506 = io_fpu_dec_ren1 & T507;
  assign T507 = T29 == io_dpath_mem_waddr;
  assign T508 = data_hazard_mem & T509;
  assign T509 = T510 | mem_reg_rocc_val;
  assign T510 = T511 | mem_reg_fp_val;
  assign T511 = T512 | mem_reg_div_mul_val;
  assign T512 = T561 | T513;
  assign T513 = mem_reg_mem_val & mem_reg_slow_bypass;
  assign T514 = T560 ? ex_slow_bypass : mem_reg_slow_bypass;
  assign ex_slow_bypass = T533 | T515;
  assign T515 = T528 | T516;
  assign T516 = 3'h5 == ex_reg_mem_type;
  assign T517 = T527 ? T518 : ex_reg_mem_type;
  assign T518 = T519;
  assign T519 = {T525, T520};
  assign T520 = {T523, T521};
  assign T521 = T522 == 32'h1000;
  assign T522 = io_dpath_inst & 32'h1000;
  assign T523 = T524 == 32'h2000;
  assign T524 = io_dpath_inst & 32'h2000;
  assign T525 = T526 == 32'h4000;
  assign T526 = io_dpath_inst & 32'h4000;
  assign T527 = ctrl_killd ^ 1'h1;
  assign T528 = T530 | T529;
  assign T529 = 3'h1 == ex_reg_mem_type;
  assign T530 = T532 | T531;
  assign T531 = 3'h4 == ex_reg_mem_type;
  assign T532 = 3'h0 == ex_reg_mem_type;
  assign T533 = ex_reg_mem_cmd == 5'h7;
  assign T534 = T527 ? T535 : ex_reg_mem_cmd;
  assign T535 = {1'h0, T536};
  assign T536 = {T558, T537};
  assign T537 = {T552, T538};
  assign T538 = {T547, T539};
  assign T539 = T542 | T540;
  assign T540 = T541 == 32'h20000020;
  assign T541 = io_dpath_inst & 32'h20000020;
  assign T542 = T545 | T543;
  assign T543 = T544 == 32'h18000020;
  assign T544 = io_dpath_inst & 32'h18000020;
  assign T545 = T546 == 32'h20;
  assign T546 = io_dpath_inst & 32'h28;
  assign T547 = T550 | T548;
  assign T548 = T549 == 32'h40000008;
  assign T549 = io_dpath_inst & 32'h40000008;
  assign T550 = T551 == 32'h10000008;
  assign T551 = io_dpath_inst & 32'h10000008;
  assign T552 = T555 | T553;
  assign T553 = T554 == 32'h80000008;
  assign T554 = io_dpath_inst & 32'h80000008;
  assign T555 = T556 | T550;
  assign T556 = T557 == 32'h8000008;
  assign T557 = io_dpath_inst & 32'h8000008;
  assign T558 = T559 == 32'h8;
  assign T559 = io_dpath_inst & 32'h18000008;
  assign T560 = ctrl_killx ^ 1'h1;
  assign T561 = mem_reg_csr != 2'h0;
  assign T562 = ctrl_killx ? 2'h0 : ex_reg_csr;
  assign T563 = ctrl_killd ? 2'h0 : T22;
  assign data_hazard_mem = mem_reg_wen & T564;
  assign T564 = T567 | T565;
  assign T565 = id_wen_not0 & T566;
  assign T566 = T116 == io_dpath_mem_waddr;
  assign T567 = T570 | T568;
  assign T568 = id_renx2_not0 & T569;
  assign T569 = T385 == io_dpath_mem_waddr;
  assign T570 = id_renx1_not0 & T571;
  assign T571 = T29 == io_dpath_mem_waddr;
  assign id_ex_hazard = T585 | T572;
  assign T572 = fp_data_hazard_ex & T573;
  assign T573 = ex_reg_mem_val | ex_reg_fp_val;
  assign fp_data_hazard_ex = ex_reg_fp_wen & T574;
  assign T574 = T577 | T575;
  assign T575 = io_fpu_dec_wen & T576;
  assign T576 = T116 == io_dpath_ex_waddr;
  assign T577 = T580 | T578;
  assign T578 = io_fpu_dec_ren3 & T579;
  assign T579 = T376 == io_dpath_ex_waddr;
  assign T580 = T583 | T581;
  assign T581 = io_fpu_dec_ren2 & T582;
  assign T582 = T385 == io_dpath_ex_waddr;
  assign T583 = io_fpu_dec_ren1 & T584;
  assign T584 = T29 == io_dpath_ex_waddr;
  assign T585 = data_hazard_ex & T586;
  assign T586 = T587 | ex_reg_rocc_val;
  assign T587 = T588 | ex_reg_fp_val;
  assign T588 = T589 | ex_reg_div_mul_val;
  assign T589 = T590 | ex_reg_mem_val;
  assign T590 = T591 | ex_reg_jalr;
  assign T591 = ex_reg_csr != 2'h0;
  assign data_hazard_ex = ex_reg_wen & T592;
  assign T592 = T595 | T593;
  assign T593 = id_wen_not0 & T594;
  assign T594 = T116 == io_dpath_ex_waddr;
  assign T595 = T598 | T596;
  assign T596 = id_renx2_not0 & T597;
  assign T597 = T385 == io_dpath_ex_waddr;
  assign T598 = id_renx1_not0 & T599;
  assign T599 = T29 == io_dpath_ex_waddr;
  assign T600 = T601 | take_pc_mem_wb;
  assign T601 = io_imem_resp_valid ^ 1'h1;
  assign T602 = wb_dcache_miss & ex_reg_load_use;
  assign T603 = ctrl_killd ? 1'h0 : id_load_use;
  assign id_load_use = T604;
  assign T604 = mem_reg_mem_val & T605;
  assign T605 = data_hazard_mem | fp_data_hazard_mem;
  assign replay_ex_structural = T608 | T606;
  assign T606 = ex_reg_div_mul_val & T607;
  assign T607 = io_dpath_div_mul_rdy ^ 1'h1;
  assign T608 = ex_reg_mem_val & T609;
  assign T609 = io_dmem_req_ready ^ 1'h1;
  assign T610 = take_pc_mem_wb ^ 1'h1;
  assign T611 = ctrl_killx ? 1'h0 : ex_reg_sret;
  assign T612 = ctrl_killd ? 1'h0 : T182;
  assign T613 = replay_wb | wb_reg_xcpt;
  assign io_rocc_s = io_dpath_status_s;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign wb_rocc_val = wb_reg_rocc_val & T614;
  assign T614 = replay_wb_common ^ 1'h1;
  assign io_fpu_killm = killm_common;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_valid = T615;
  assign T615 = T616 & T152;
  assign T616 = ctrl_killd ^ 1'h1;
  assign io_dmem_req_bits_cmd = ex_reg_mem_cmd;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_typ = ex_reg_mem_type;
  assign io_dmem_req_bits_kill = T617;
  assign T617 = killm_common | mem_xcpt;
  assign io_dmem_req_valid = ex_reg_mem_val;
  assign io_imem_invalidate = wb_reg_flush_inst;
  assign T618 = ctrl_killm ? 1'h0 : mem_reg_flush_inst;
  assign T619 = ctrl_killx ? 1'h0 : ex_reg_flush_inst;
  assign T620 = ctrl_killd ? 1'h0 : T101;
  assign io_imem_btb_update_bits_incorrectTarget = take_pc_mem;
  assign io_imem_btb_update_bits_isReturn = T621;
  assign T621 = mem_reg_jalr & io_dpath_mem_rs1_ra;
  assign io_imem_btb_update_bits_isCall = T622;
  assign T622 = mem_reg_wen & T623;
  assign T623 = io_dpath_mem_waddr[1'h0:1'h0];
  assign io_imem_btb_update_bits_isJump = T624;
  assign T624 = mem_reg_jal | mem_reg_jalr;
  assign io_imem_btb_update_bits_taken = T625;
  assign T625 = mem_reg_jal | T626;
  assign T626 = mem_reg_branch & io_dpath_mem_br_taken;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign T627 = T630 ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T628 = T629 ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T629 = T527 & io_imem_btb_resp_valid;
  assign T630 = T560 & ex_reg_btb_hit;
  assign T631 = ctrl_killd ? 1'h0 : io_imem_btb_resp_valid;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = mem_reg_btb_resp_bht_index;
  assign T632 = T630 ? ex_reg_btb_resp_bht_index : mem_reg_btb_resp_bht_index;
  assign T633 = T629 ? io_imem_btb_resp_bits_bht_index : ex_reg_btb_resp_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign T634 = T630 ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign T635 = T629 ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign T636 = T630 ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign T637 = T629 ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign T638 = T630 ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign T639 = T629 ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign T640 = T560 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign io_imem_btb_update_valid = T641;
  assign T641 = T642 | mem_reg_jalr;
  assign T642 = mem_reg_branch | mem_reg_jal;
  assign io_imem_resp_ready = T643;
  assign T643 = T644 | ctrl_draind;
  assign T644 = ctrl_stalld ^ 1'h1;
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_dpath_badvaddr_wen = wb_reg_xcpt;
  assign io_dpath_cause = wb_reg_cause;
  assign T645 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign mem_cause = T166 ? mem_reg_cause : T646;
  assign T646 = {60'h0, T647};
  assign T647 = T165 ? 4'h8 : T648;
  assign T648 = T163 ? 4'h9 : T649;
  assign T649 = T161 ? 4'ha : 4'hb;
  assign T650 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign ex_cause = T169 ? ex_reg_cause : 64'h2;
  assign T651 = id_xcpt ? id_cause : ex_reg_cause;
  assign id_cause = id_interrupt ? id_interrupt_cause : T652;
  assign T652 = {60'h0, T653};
  assign T653 = io_imem_resp_bits_xcpt_ma ? 4'h0 : T654;
  assign T654 = io_imem_resp_bits_xcpt_if ? 4'h1 : T655;
  assign T655 = T206 ? 4'h2 : T656;
  assign T656 = id_csr_privileged ? 4'h3 : T657;
  assign T657 = T180 ? 4'h3 : T658;
  assign T658 = T174 ? 4'h4 : T659;
  assign T659 = T171 ? 4'h6 : 4'hc;
  assign id_interrupt_cause = T61 ? 64'h8000000000000000 : T660;
  assign T660 = T58 ? 64'h8000000000000001 : T661;
  assign T661 = T54 ? 64'h8000000000000002 : T662;
  assign T662 = T50 ? 64'h8000000000000003 : T663;
  assign T663 = T46 ? 64'h8000000000000004 : T664;
  assign T664 = T42 ? 64'h8000000000000005 : T665;
  assign T665 = T38 ? 64'h8000000000000006 : 64'h8000000000000007;
  assign io_dpath_exception = wb_reg_xcpt;
  assign io_dpath_retire = T666;
  assign T666 = wb_reg_valid & T667;
  assign T667 = replay_wb ^ 1'h1;
  assign T668 = ctrl_killm ? 1'h0 : mem_reg_valid;
  assign io_dpath_ll_ready = T669;
  assign T669 = wb_reg_wen ^ 1'h1;
  assign io_dpath_bypass_src_0 = T670;
  assign T670 = T679 ? 2'h0 : T671;
  assign T671 = T677 ? 2'h1 : T672;
  assign T672 = T673 ? 2'h2 : 2'h3;
  assign T673 = T675 & T674;
  assign T674 = io_dpath_mem_waddr == T29;
  assign T675 = mem_reg_wen & T676;
  assign T676 = mem_reg_mem_val ^ 1'h1;
  assign T677 = ex_reg_wen & T678;
  assign T678 = io_dpath_ex_waddr == T29;
  assign T679 = 5'h0 == T29;
  assign io_dpath_bypass_src_1 = T680;
  assign T680 = T687 ? 2'h0 : T681;
  assign T681 = T685 ? 2'h1 : T682;
  assign T682 = T683 ? 2'h2 : 2'h3;
  assign T683 = T675 & T684;
  assign T684 = io_dpath_mem_waddr == T385;
  assign T685 = ex_reg_wen & T686;
  assign T686 = io_dpath_ex_waddr == T385;
  assign T687 = 5'h0 == T385;
  assign io_dpath_bypass_0 = T688;
  assign T688 = T691 | T689;
  assign T689 = mem_reg_wen & T690;
  assign T690 = io_dpath_mem_waddr == T29;
  assign T691 = T692 | T673;
  assign T692 = T679 | T677;
  assign io_dpath_bypass_1 = T693;
  assign T693 = T696 | T694;
  assign T694 = mem_reg_wen & T695;
  assign T695 = io_dpath_mem_waddr == T385;
  assign T696 = T697 | T683;
  assign T697 = T687 | T685;
  assign io_dpath_mem_rocc_val = mem_reg_rocc_val;
  assign io_dpath_ex_rocc_val = ex_reg_rocc_val;
  assign io_dpath_ex_rs2_val = T698;
  assign T698 = T699 | ex_reg_rocc_val;
  assign T699 = ex_reg_mem_val & T700;
  assign T700 = T704 | T701;
  assign T701 = T703 | T702;
  assign T702 = ex_reg_mem_cmd == 5'h4;
  assign T703 = ex_reg_mem_cmd[2'h3:2'h3];
  assign T704 = T706 | T705;
  assign T705 = ex_reg_mem_cmd == 5'h7;
  assign T706 = ex_reg_mem_cmd == 5'h1;
  assign io_dpath_ex_mem_type = ex_reg_mem_type;
  assign io_dpath_wb_wen = T707;
  assign T707 = wb_reg_wen & T708;
  assign T708 = replay_wb ^ 1'h1;
  assign io_dpath_mem_wen = mem_reg_wen;
  assign io_dpath_mem_branch = mem_reg_branch;
  assign io_dpath_mem_jalr = mem_reg_jalr;
  assign io_dpath_ex_valid = ex_reg_valid;
  assign io_dpath_ex_wen = ex_reg_wen;
  assign io_dpath_mem_fp_val = mem_reg_fp_val;
  assign io_dpath_ex_fp_val = ex_reg_fp_val;
  assign io_dpath_wb_load = T709;
  assign T709 = wb_reg_mem_val & wb_reg_wen;
  assign io_dpath_mem_load = T710;
  assign T710 = mem_reg_mem_val & mem_reg_wen;
  assign io_dpath_sret = wb_reg_sret;
  assign io_dpath_csr = T711;
  assign T711 = {1'h0, wb_reg_csr};
  assign T712 = ctrl_killm ? 2'h0 : mem_reg_csr;
  assign io_dpath_div_mul_kill = T713;
  assign T713 = mem_reg_div_mul_val & killm_common;
  assign io_dpath_div_mul_val = ex_reg_div_mul_val;
  assign io_dpath_fn_alu = T714;
  assign T714 = T715;
  assign T715 = {T751, T716};
  assign T716 = {T740, T717};
  assign T717 = {T726, T718};
  assign T718 = T721 | T719;
  assign T719 = T720 == 32'h7000;
  assign T720 = io_dpath_inst & 32'h7044;
  assign T721 = T724 | T722;
  assign T722 = T723 == 32'h1040;
  assign T723 = io_dpath_inst & 32'h1058;
  assign T724 = T725 == 32'h1010;
  assign T725 = io_dpath_inst & 32'h3054;
  assign T726 = T729 | T727;
  assign T727 = T728 == 32'h40001010;
  assign T728 = io_dpath_inst & 32'h40001054;
  assign T729 = T732 | T730;
  assign T730 = T731 == 32'h40000030;
  assign T731 = io_dpath_inst & 32'h40003034;
  assign T732 = T735 | T733;
  assign T733 = T734 == 32'h6010;
  assign T734 = io_dpath_inst & 32'h6054;
  assign T735 = T738 | T736;
  assign T736 = T737 == 32'h3010;
  assign T737 = io_dpath_inst & 32'h3054;
  assign T738 = T739 == 32'h2040;
  assign T739 = io_dpath_inst & 32'h2058;
  assign T740 = T743 | T741;
  assign T741 = T742 == 32'h4040;
  assign T742 = io_dpath_inst & 32'h4058;
  assign T743 = T746 | T744;
  assign T744 = T745 == 32'h4010;
  assign T745 = io_dpath_inst & 32'h5054;
  assign T746 = T749 | T747;
  assign T747 = T748 == 32'h4010;
  assign T748 = io_dpath_inst & 32'h40004054;
  assign T749 = T750 == 32'h2010;
  assign T750 = io_dpath_inst & 32'h2054;
  assign T751 = T754 | T752;
  assign T752 = T753 == 32'h40001010;
  assign T753 = io_dpath_inst & 32'h40003054;
  assign T754 = T755 | T730;
  assign T755 = T758 | T756;
  assign T756 = T757 == 32'h2010;
  assign T757 = io_dpath_inst & 32'h6054;
  assign T758 = T759 == 32'h40;
  assign T759 = io_dpath_inst & 32'h54;
  assign io_dpath_fn_dw = T760;
  assign T760 = T761;
  assign T761 = T764 | T762;
  assign T762 = T763 == 32'h0;
  assign T763 = io_dpath_inst & 32'h8;
  assign T764 = T765 == 32'h0;
  assign T765 = io_dpath_inst & 32'h10;
  assign io_dpath_sel_imm = T766;
  assign T766 = T767;
  assign T767 = {T777, T768};
  assign T768 = {T774, T769};
  assign T769 = T772 | T770;
  assign T770 = T771 == 32'h40;
  assign T771 = io_dpath_inst & 32'h44;
  assign T772 = T773 == 32'h8;
  assign T773 = io_dpath_inst & 32'h18;
  assign T774 = T772 | T775;
  assign T775 = T776 == 32'h14;
  assign T776 = io_dpath_inst & 32'h14;
  assign T777 = T780 | T778;
  assign T778 = T779 == 32'h10;
  assign T779 = io_dpath_inst & 32'h14;
  assign T780 = T783 | T781;
  assign T781 = T782 == 32'h4;
  assign T782 = io_dpath_inst & 32'h201c;
  assign T783 = T784 == 32'h0;
  assign T784 = io_dpath_inst & 32'h30;
  assign io_dpath_sel_alu1 = T785;
  assign T785 = T786;
  assign T786 = {T799, T787};
  assign T787 = T790 | T788;
  assign T788 = T789 == 32'h0;
  assign T789 = io_dpath_inst & 32'h18;
  assign T790 = T793 | T791;
  assign T791 = T792 == 32'h0;
  assign T792 = io_dpath_inst & 32'h24;
  assign T793 = T794 | T468;
  assign T794 = T797 | T795;
  assign T795 = T796 == 32'h0;
  assign T796 = io_dpath_inst & 32'h50;
  assign T797 = T798 == 32'h0;
  assign T798 = io_dpath_inst & 32'h4004;
  assign T799 = T802 | T800;
  assign T800 = T801 == 32'h48;
  assign T801 = io_dpath_inst & 32'h48;
  assign T802 = T803 == 32'h14;
  assign T803 = io_dpath_inst & 32'h34;
  assign io_dpath_sel_alu2 = T804;
  assign T804 = {1'h0, T805};
  assign T805 = T806;
  assign T806 = {T819, T807};
  assign T807 = T810 | T808;
  assign T808 = T809 == 32'h4050;
  assign T809 = io_dpath_inst & 32'h4050;
  assign T810 = T811 | T800;
  assign T811 = T814 | T812;
  assign T812 = T813 == 32'h4;
  assign T813 = io_dpath_inst & 32'hc;
  assign T814 = T817 | T815;
  assign T815 = T816 == 32'h0;
  assign T816 = io_dpath_inst & 32'h20;
  assign T817 = T818 == 32'h0;
  assign T818 = io_dpath_inst & 32'h58;
  assign T819 = T822 | T820;
  assign T820 = T821 == 32'h4000;
  assign T821 = io_dpath_inst & 32'h4008;
  assign T822 = T823 | T788;
  assign T823 = T824 | T468;
  assign T824 = T825 == 32'h0;
  assign T825 = io_dpath_inst & 32'h48;
  assign io_dpath_ren_0 = T453;
  assign io_dpath_ren_1 = T437;
  assign io_dpath_killd = T826;
  assign T826 = take_pc_mem_wb | T827;
  assign T827 = ctrl_stalld & T828;
  assign T828 = ctrl_draind ^ 1'h1;
  assign io_dpath_sel_pc = T829;
  assign T829 = {1'h0, T830};
  assign T830 = wb_reg_xcpt ? 2'h3 : T831;
  assign T831 = wb_reg_sret ? 2'h3 : T832;
  assign T832 = replay_wb ? 2'h2 : 2'h1;

  always @(posedge clk) begin
    wb_reg_xcpt <= T1;
    if(ctrl_killm) begin
      wb_reg_sret <= 1'h0;
    end else begin
      wb_reg_sret <= T5;
    end
    mem_reg_replay <= T7;
    if(ctrl_killx) begin
      mem_reg_replay_next <= 1'h0;
    end else begin
      mem_reg_replay_next <= ex_reg_replay_next;
    end
    if(ctrl_killd) begin
      ex_reg_replay_next <= 1'h0;
    end else begin
      ex_reg_replay_next <= T10;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T89;
    end
    if(ctrl_killd) begin
      ex_reg_mem_val <= 1'h0;
    end else begin
      ex_reg_mem_val <= T92;
    end
    if(reset) begin
      R118 <= 32'h0;
    end else if(T368) begin
      R118 <= T364;
    end else if(T363) begin
      R118 <= T359;
    end else if(T126) begin
      R118 <= T123;
    end
    if(ctrl_killm) begin
      wb_reg_rocc_val <= 1'h0;
    end else begin
      wb_reg_rocc_val <= mem_reg_rocc_val;
    end
    if(ctrl_killx) begin
      mem_reg_rocc_val <= 1'h0;
    end else begin
      mem_reg_rocc_val <= ex_reg_rocc_val;
    end
    if(ctrl_killd) begin
      ex_reg_rocc_val <= 1'h0;
    end else begin
      ex_reg_rocc_val <= T133;
    end
    if(ctrl_killx) begin
      mem_reg_jal <= 1'h0;
    end else begin
      mem_reg_jal <= ex_reg_jal;
    end
    if(ctrl_killd) begin
      ex_reg_jal <= 1'h0;
    end else begin
      ex_reg_jal <= T138;
    end
    if(ctrl_killx) begin
      mem_reg_jalr <= 1'h0;
    end else begin
      mem_reg_jalr <= ex_reg_jalr;
    end
    if(ctrl_killd) begin
      ex_reg_jalr <= 1'h0;
    end else begin
      ex_reg_jalr <= T143;
    end
    if(ctrl_killx) begin
      mem_reg_branch <= 1'h0;
    end else begin
      mem_reg_branch <= ex_reg_branch;
    end
    if(ctrl_killd) begin
      ex_reg_branch <= 1'h0;
    end else begin
      ex_reg_branch <= T147;
    end
    if(ctrl_killx) begin
      mem_reg_fp_val <= 1'h0;
    end else begin
      mem_reg_fp_val <= ex_reg_fp_val;
    end
    if(ctrl_killd) begin
      ex_reg_fp_val <= 1'h0;
    end else begin
      ex_reg_fp_val <= T152;
    end
    if(ctrl_killx) begin
      mem_reg_mem_val <= 1'h0;
    end else begin
      mem_reg_mem_val <= ex_reg_mem_val;
    end
    if(ctrl_killx) begin
      mem_reg_xcpt <= 1'h0;
    end else begin
      mem_reg_xcpt <= ex_xcpt;
    end
    if(ctrl_killd) begin
      ex_reg_xcpt <= 1'h0;
    end else begin
      ex_reg_xcpt <= id_xcpt;
    end
    ex_reg_xcpt_interrupt <= T313;
    mem_reg_xcpt_interrupt <= T316;
    if(ctrl_killx) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= ex_reg_valid;
    end
    if(ctrl_killd) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= 1'h1;
    end
    if(ctrl_killx) begin
      mem_reg_wen <= 1'h0;
    end else begin
      mem_reg_wen <= ex_reg_wen;
    end
    if(ctrl_killd) begin
      ex_reg_wen <= 1'h0;
    end else begin
      ex_reg_wen <= T327;
    end
    wb_reg_replay <= T348;
    if(ctrl_killm) begin
      wb_reg_fp_wen <= 1'h0;
    end else begin
      wb_reg_fp_wen <= mem_reg_fp_wen;
    end
    if(ctrl_killx) begin
      mem_reg_fp_wen <= 1'h0;
    end else begin
      mem_reg_fp_wen <= ex_reg_fp_wen;
    end
    if(ctrl_killd) begin
      ex_reg_fp_wen <= 1'h0;
    end else begin
      ex_reg_fp_wen <= T356;
    end
    if(ctrl_killm) begin
      wb_reg_mem_val <= 1'h0;
    end else begin
      wb_reg_mem_val <= mem_reg_mem_val;
    end
    if(reset) begin
      R409 <= 32'h0;
    end else if(T426) begin
      R409 <= T413;
    end else if(io_dpath_ll_wen) begin
      R409 <= T405;
    end
    if(ctrl_killm) begin
      wb_reg_div_mul_val <= 1'h0;
    end else begin
      wb_reg_div_mul_val <= mem_reg_div_mul_val;
    end
    mem_reg_div_mul_val <= T419;
    if(ctrl_killd) begin
      ex_reg_div_mul_val <= 1'h0;
    end else begin
      ex_reg_div_mul_val <= T421;
    end
    if(ctrl_killm) begin
      wb_reg_fp_val <= 1'h0;
    end else begin
      wb_reg_fp_val <= mem_reg_fp_val;
    end
    if(ctrl_killm) begin
      wb_reg_wen <= 1'h0;
    end else begin
      wb_reg_wen <= mem_reg_wen;
    end
    if(T560) begin
      mem_reg_slow_bypass <= ex_slow_bypass;
    end
    if(T527) begin
      ex_reg_mem_type <= T518;
    end
    if(T527) begin
      ex_reg_mem_cmd <= T535;
    end
    if(ctrl_killx) begin
      mem_reg_csr <= 2'h0;
    end else begin
      mem_reg_csr <= ex_reg_csr;
    end
    if(ctrl_killd) begin
      ex_reg_csr <= 2'h0;
    end else begin
      ex_reg_csr <= T22;
    end
    if(ctrl_killd) begin
      ex_reg_load_use <= 1'h0;
    end else begin
      ex_reg_load_use <= id_load_use;
    end
    if(ctrl_killx) begin
      mem_reg_sret <= 1'h0;
    end else begin
      mem_reg_sret <= ex_reg_sret;
    end
    if(ctrl_killd) begin
      ex_reg_sret <= 1'h0;
    end else begin
      ex_reg_sret <= T182;
    end
    if(ctrl_killm) begin
      wb_reg_flush_inst <= 1'h0;
    end else begin
      wb_reg_flush_inst <= mem_reg_flush_inst;
    end
    if(ctrl_killx) begin
      mem_reg_flush_inst <= 1'h0;
    end else begin
      mem_reg_flush_inst <= ex_reg_flush_inst;
    end
    if(ctrl_killd) begin
      ex_reg_flush_inst <= 1'h0;
    end else begin
      ex_reg_flush_inst <= T101;
    end
    if(T630) begin
      mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
    end
    if(T629) begin
      ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
    end
    if(ctrl_killd) begin
      ex_reg_btb_hit <= 1'h0;
    end else begin
      ex_reg_btb_hit <= io_imem_btb_resp_valid;
    end
    if(T630) begin
      mem_reg_btb_resp_bht_index <= ex_reg_btb_resp_bht_index;
    end
    if(T629) begin
      ex_reg_btb_resp_bht_index <= io_imem_btb_resp_bits_bht_index;
    end
    if(T630) begin
      mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
    end
    if(T629) begin
      ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
    end
    if(T630) begin
      mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
    end
    if(T629) begin
      ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
    end
    if(T630) begin
      mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
    end
    if(T629) begin
      ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
    end
    if(T560) begin
      mem_reg_btb_hit <= ex_reg_btb_hit;
    end
    if(mem_xcpt) begin
      wb_reg_cause <= mem_cause;
    end
    if(ex_xcpt) begin
      mem_reg_cause <= ex_cause;
    end
    if(id_xcpt) begin
      ex_reg_cause <= id_cause;
    end
    if(ctrl_killm) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= mem_reg_valid;
    end
    if(ctrl_killm) begin
      wb_reg_csr <= 2'h0;
    end else begin
      wb_reg_csr <= mem_reg_csr;
    end
  end
endmodule

module ALU(
    input  io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output[63:0] io_out,
    output[63:0] io_adder_out
);

  wire[63:0] sum;
  wire[63:0] T0;
  wire[63:0] T1;
  wire T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[31:0] T5;
  wire[63:0] out64;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T11;
  wire cmp;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire[63:0] T26;
  wire T27;
  wire[63:0] T28;
  wire T29;
  wire[63:0] T30;
  wire T31;
  wire[63:0] shout_l;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[62:0] T34;
  wire[63:0] T35;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[61:0] T38;
  wire[63:0] T39;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[59:0] T42;
  wire[63:0] T43;
  wire[63:0] T44;
  wire[63:0] T45;
  wire[55:0] T46;
  wire[63:0] T47;
  wire[63:0] T48;
  wire[63:0] T49;
  wire[47:0] T50;
  wire[63:0] T51;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[31:0] T54;
  wire[63:0] T55;
  wire[64:0] T56;
  wire[5:0] shamt;
  wire[5:0] T57;
  wire[4:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[64:0] T62;
  wire[64:0] T63;
  wire[63:0] shin;
  wire[63:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire[62:0] T67;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[61:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[59:0] T75;
  wire[63:0] T76;
  wire[63:0] T77;
  wire[63:0] T78;
  wire[55:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[47:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[31:0] T87;
  wire[63:0] shin_r;
  wire[31:0] T88;
  wire[31:0] shin_hi;
  wire[31:0] shin_hi_32;
  wire[31:0] T89;
  wire[31:0] T90;
  wire T91;
  wire T92;
  wire[31:0] T93;
  wire T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire[31:0] T97;
  wire[63:0] T98;
  wire[63:0] T99;
  wire[47:0] T100;
  wire[63:0] T101;
  wire[63:0] T102;
  wire[55:0] T103;
  wire[63:0] T104;
  wire[63:0] T105;
  wire[59:0] T106;
  wire[63:0] T107;
  wire[63:0] T108;
  wire[61:0] T109;
  wire[63:0] T110;
  wire[63:0] T111;
  wire[62:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire[63:0] T119;
  wire[63:0] T120;
  wire[31:0] T121;
  wire[63:0] T122;
  wire[63:0] T123;
  wire[47:0] T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire[55:0] T127;
  wire[63:0] T128;
  wire[63:0] T129;
  wire[59:0] T130;
  wire[63:0] T131;
  wire[63:0] T132;
  wire[61:0] T133;
  wire[63:0] T134;
  wire[63:0] T135;
  wire[62:0] T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire[31:0] out_hi;
  wire[31:0] T144;
  wire[31:0] T145;
  wire T146;
  wire[31:0] T147;
  wire T148;


  assign io_adder_out = sum;
  assign sum = io_in1 + T0;
  assign T0 = T2 ? T1 : io_in2;
  assign T1 = 64'h0 - io_in2;
  assign T2 = io_fn[2'h3:2'h3];
  assign io_out = T3;
  assign T3 = T4;
  assign T4 = {out_hi, T5};
  assign T5 = out64[5'h1f:1'h0];
  assign out64 = T141 ? sum : T6;
  assign T6 = T138 ? T55 : T7;
  assign T7 = T137 ? shout_l : T8;
  assign T8 = T31 ? T30 : T9;
  assign T9 = T29 ? T28 : T10;
  assign T10 = T27 ? T26 : T11;
  assign T11 = {63'h0, cmp};
  assign cmp = T25 ^ T12;
  assign T12 = T23 ? T22 : T13;
  assign T13 = T19 ? T18 : T14;
  assign T14 = T17 ? T16 : T15;
  assign T15 = io_in1[6'h3f:6'h3f];
  assign T16 = io_in2[6'h3f:6'h3f];
  assign T17 = io_fn[1'h1:1'h1];
  assign T18 = sum[6'h3f:6'h3f];
  assign T19 = T21 == T20;
  assign T20 = io_in2[6'h3f:6'h3f];
  assign T21 = io_in1[6'h3f:6'h3f];
  assign T22 = sum == 64'h0;
  assign T23 = T24 ^ 1'h1;
  assign T24 = io_fn[2'h2:2'h2];
  assign T25 = io_fn[1'h0:1'h0];
  assign T26 = io_in1 ^ io_in2;
  assign T27 = io_fn == 4'h4;
  assign T28 = io_in1 | io_in2;
  assign T29 = io_fn == 4'h6;
  assign T30 = io_in1 & io_in2;
  assign T31 = io_fn == 4'h7;
  assign shout_l = T134 | T32;
  assign T32 = T33 & 64'haaaaaaaaaaaaaaaa;
  assign T33 = T34 << 1'h1;
  assign T34 = T35[6'h3e:1'h0];
  assign T35 = T131 | T36;
  assign T36 = T37 & 64'hcccccccccccccccc;
  assign T37 = T38 << 2'h2;
  assign T38 = T39[6'h3d:1'h0];
  assign T39 = T128 | T40;
  assign T40 = T41 & 64'hf0f0f0f0f0f0f0f0;
  assign T41 = T42 << 3'h4;
  assign T42 = T43[6'h3b:1'h0];
  assign T43 = T125 | T44;
  assign T44 = T45 & 64'hff00ff00ff00ff00;
  assign T45 = T46 << 4'h8;
  assign T46 = T47[6'h37:1'h0];
  assign T47 = T122 | T48;
  assign T48 = T49 & 64'hffff0000ffff0000;
  assign T49 = T50 << 5'h10;
  assign T50 = T51[6'h2f:1'h0];
  assign T51 = T119 | T52;
  assign T52 = T53 & 64'hffffffff00000000;
  assign T53 = T54 << 6'h20;
  assign T54 = T55[5'h1f:1'h0];
  assign T55 = T56[6'h3f:1'h0];
  assign T56 = $signed(T62) >>> shamt;
  assign shamt = T57;
  assign T57 = {T59, T58};
  assign T58 = io_in2[3'h4:1'h0];
  assign T59 = T61 & T60;
  assign T60 = io_dw == 1'h1;
  assign T61 = io_in2[3'h5:3'h5];
  assign T62 = T63;
  assign T63 = {T116, shin};
  assign shin = T113 ? shin_r : T64;
  assign T64 = T110 | T65;
  assign T65 = T66 & 64'haaaaaaaaaaaaaaaa;
  assign T66 = T67 << 1'h1;
  assign T67 = T68[6'h3e:1'h0];
  assign T68 = T107 | T69;
  assign T69 = T70 & 64'hcccccccccccccccc;
  assign T70 = T71 << 2'h2;
  assign T71 = T72[6'h3d:1'h0];
  assign T72 = T104 | T73;
  assign T73 = T74 & 64'hf0f0f0f0f0f0f0f0;
  assign T74 = T75 << 3'h4;
  assign T75 = T76[6'h3b:1'h0];
  assign T76 = T101 | T77;
  assign T77 = T78 & 64'hff00ff00ff00ff00;
  assign T78 = T79 << 4'h8;
  assign T79 = T80[6'h37:1'h0];
  assign T80 = T98 | T81;
  assign T81 = T82 & 64'hffff0000ffff0000;
  assign T82 = T83 << 5'h10;
  assign T83 = T84[6'h2f:1'h0];
  assign T84 = T95 | T85;
  assign T85 = T86 & 64'hffffffff00000000;
  assign T86 = T87 << 6'h20;
  assign T87 = shin_r[5'h1f:1'h0];
  assign shin_r = {shin_hi, T88};
  assign T88 = io_in1[5'h1f:1'h0];
  assign shin_hi = T94 ? T93 : shin_hi_32;
  assign shin_hi_32 = T92 ? T89 : 32'h0;
  assign T89 = 32'h0 - T90;
  assign T90 = {31'h0, T91};
  assign T91 = io_in1[5'h1f:5'h1f];
  assign T92 = io_fn[2'h3:2'h3];
  assign T93 = io_in1[6'h3f:6'h20];
  assign T94 = io_dw == 1'h1;
  assign T95 = T96 & 64'hffffffff;
  assign T96 = {32'h0, T97};
  assign T97 = shin_r >> 6'h20;
  assign T98 = T99 & 64'hffff0000ffff;
  assign T99 = {16'h0, T100};
  assign T100 = T84 >> 5'h10;
  assign T101 = T102 & 64'hff00ff00ff00ff;
  assign T102 = {8'h0, T103};
  assign T103 = T80 >> 4'h8;
  assign T104 = T105 & 64'hf0f0f0f0f0f0f0f;
  assign T105 = {4'h0, T106};
  assign T106 = T76 >> 3'h4;
  assign T107 = T108 & 64'h3333333333333333;
  assign T108 = {2'h0, T109};
  assign T109 = T72 >> 2'h2;
  assign T110 = T111 & 64'h5555555555555555;
  assign T111 = {1'h0, T112};
  assign T112 = T68 >> 1'h1;
  assign T113 = T115 | T114;
  assign T114 = io_fn == 4'hb;
  assign T115 = io_fn == 4'h5;
  assign T116 = T118 & T117;
  assign T117 = shin[6'h3f:6'h3f];
  assign T118 = io_fn[2'h3:2'h3];
  assign T119 = T120 & 64'hffffffff;
  assign T120 = {32'h0, T121};
  assign T121 = T55 >> 6'h20;
  assign T122 = T123 & 64'hffff0000ffff;
  assign T123 = {16'h0, T124};
  assign T124 = T51 >> 5'h10;
  assign T125 = T126 & 64'hff00ff00ff00ff;
  assign T126 = {8'h0, T127};
  assign T127 = T47 >> 4'h8;
  assign T128 = T129 & 64'hf0f0f0f0f0f0f0f;
  assign T129 = {4'h0, T130};
  assign T130 = T43 >> 3'h4;
  assign T131 = T132 & 64'h3333333333333333;
  assign T132 = {2'h0, T133};
  assign T133 = T39 >> 2'h2;
  assign T134 = T135 & 64'h5555555555555555;
  assign T135 = {1'h0, T136};
  assign T136 = T35 >> 1'h1;
  assign T137 = io_fn == 4'h1;
  assign T138 = T140 | T139;
  assign T139 = io_fn == 4'hb;
  assign T140 = io_fn == 4'h5;
  assign T141 = T143 | T142;
  assign T142 = io_fn == 4'ha;
  assign T143 = io_fn == 4'h0;
  assign out_hi = T148 ? T147 : T144;
  assign T144 = 32'h0 - T145;
  assign T145 = {31'h0, T146};
  assign T146 = out64[5'h1f:5'h1f];
  assign T147 = out64[6'h3f:6'h20];
  assign T148 = io_dw == 1'h1;
endmodule

module MulDiv(input clk, input reset,
    output io_req_ready,
    input  io_req_valid,
    input [3:0] io_req_bits_fn,
    input  io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input  io_kill,
    input  io_resp_ready,
    output io_resp_valid,
    output[63:0] io_resp_bits_data,
    output[4:0] io_resp_bits_tag
);

  reg [4:0] req_tag;
  wire[4:0] T0;
  wire T1;
  wire[63:0] T2;
  wire[63:0] T3;
  reg [129:0] remainder;
  wire[129:0] T4;
  wire[129:0] T5;
  wire[129:0] T6;
  wire[129:0] T7;
  wire[129:0] T8;
  wire[129:0] T9;
  wire[129:0] T10;
  wire[63:0] negated_remainder;
  wire[63:0] T11;
  wire T12;
  wire T13;
  reg  isMul;
  wire T14;
  wire T15;
  wire T16;
  wire[3:0] T17;
  wire T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  reg [2:0] state;
  wire[2:0] T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire[2:0] T26;
  wire[2:0] T27;
  wire[2:0] T28;
  wire[2:0] T29;
  wire T30;
  wire[2:0] T31;
  reg  neg_out;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  isHi;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire[3:0] T41;
  wire T42;
  wire[3:0] T43;
  wire T44;
  wire T45;
  wire T46;
  wire[64:0] subtractor;
  reg [64:0] divisor;
  wire[64:0] T47;
  wire[64:0] T48;
  wire T49;
  wire T50;
  wire T51;
  wire[64:0] T52;
  wire[63:0] rhs_in;
  wire[31:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[31:0] T56;
  wire rhs_sign;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire[3:0] T63;
  wire[31:0] T64;
  wire T65;
  wire[64:0] T66;
  wire T67;
  reg [6:0] count;
  wire[6:0] T68;
  wire[6:0] T69;
  wire[6:0] T70;
  wire[6:0] T71;
  wire T72;
  wire T73;
  wire[6:0] T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire lhs_sign;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[3:0] T87;
  wire T88;
  wire T89;
  wire T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire[2:0] T94;
  wire[2:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[2:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire[129:0] T104;
  wire[129:0] T105;
  wire[63:0] T106;
  wire[129:0] T107;
  wire[129:0] T108;
  wire[64:0] T109;
  wire[63:0] T110;
  wire[128:0] T111;
  wire[63:0] T112;
  wire[128:0] T113;
  wire[128:0] T114;
  wire[62:0] T115;
  wire[63:0] T116;
  wire[128:0] T117;
  wire[63:0] T118;
  wire[64:0] T119;
  wire[65:0] T120;
  wire[65:0] T121;
  wire[64:0] T122;
  wire[64:0] T123;
  wire T124;
  wire[65:0] T125;
  wire[1:0] T126;
  wire[1:0] T127;
  wire T128;
  wire[64:0] T129;
  wire[64:0] T130;
  wire[64:0] T131;
  wire[129:0] T132;
  wire[128:0] T133;
  wire[64:0] T134;
  wire T135;
  wire[63:0] T136;
  wire[63:0] T137;
  wire[63:0] T138;
  wire[63:0] T139;
  wire[129:0] T140;
  wire[63:0] lhs_in;
  wire[31:0] T141;
  wire[31:0] T142;
  wire[31:0] T143;
  wire[31:0] T144;
  wire[31:0] T145;
  wire T146;
  wire[63:0] T147;
  wire[31:0] T148;
  wire[31:0] T149;
  wire[31:0] T150;
  wire T151;
  wire T152;
  reg  req_dw;
  wire T153;
  wire T154;
  wire T155;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    req_tag = {1{$random}};
    remainder = {5{$random}};
    isMul = {1{$random}};
    state = {1{$random}};
    neg_out = {1{$random}};
    isHi = {1{$random}};
    divisor = {3{$random}};
    count = {1{$random}};
    req_dw = {1{$random}};
  end
`endif

  assign io_resp_bits_tag = req_tag;
  assign T0 = T1 ? io_req_bits_tag : req_tag;
  assign T1 = io_req_ready & io_req_valid;
  assign io_resp_bits_data = T2;
  assign T2 = T152 ? T147 : T3;
  assign T3 = remainder[6'h3f:1'h0];
  assign T4 = T1 ? T140 : T5;
  assign T5 = T75 ? T132 : T6;
  assign T6 = T72 ? T107 : T7;
  assign T7 = T90 ? T105 : T8;
  assign T8 = T30 ? T104 : T9;
  assign T9 = T12 ? T10 : remainder;
  assign T10 = {66'h0, negated_remainder};
  assign negated_remainder = 64'h0 - T11;
  assign T11 = remainder[6'h3f:1'h0];
  assign T12 = T21 & T13;
  assign T13 = T20 | isMul;
  assign T14 = T1 ? T15 : isMul;
  assign T15 = T18 | T16;
  assign T16 = T17 == 4'h8;
  assign T17 = io_req_bits_fn & 4'h8;
  assign T18 = T19 == 4'h0;
  assign T19 = io_req_bits_fn & 4'h4;
  assign T20 = remainder[6'h3f:6'h3f];
  assign T21 = state == 3'h1;
  assign T22 = reset ? 3'h0 : T23;
  assign T23 = T1 ? T100 : T24;
  assign T24 = T98 ? 3'h0 : T25;
  assign T25 = T96 ? T94 : T26;
  assign T26 = T92 ? T91 : T27;
  assign T27 = T90 ? T31 : T28;
  assign T28 = T30 ? 3'h5 : T29;
  assign T29 = T21 ? 3'h2 : state;
  assign T30 = state == 3'h4;
  assign T31 = neg_out ? 3'h4 : 3'h5;
  assign T32 = T1 ? T78 : T33;
  assign T33 = T34 ? 1'h0 : neg_out;
  assign T34 = T75 & T35;
  assign T35 = T44 & T36;
  assign T36 = isHi ^ 1'h1;
  assign T37 = T1 ? T38 : isHi;
  assign T38 = T39 | T16;
  assign T39 = T42 | T40;
  assign T40 = T41 == 4'h2;
  assign T41 = io_req_bits_fn & 4'h2;
  assign T42 = T43 == 4'h1;
  assign T43 = io_req_bits_fn & 4'h5;
  assign T44 = T67 & T45;
  assign T45 = T46 ^ 1'h1;
  assign T46 = subtractor[7'h40:7'h40];
  assign subtractor = T66 - divisor;
  assign T47 = T1 ? T52 : T48;
  assign T48 = T49 ? subtractor : divisor;
  assign T49 = T21 & T50;
  assign T50 = T51 | isMul;
  assign T51 = divisor[6'h3f:6'h3f];
  assign T52 = {rhs_sign, rhs_in};
  assign rhs_in = {T54, T53};
  assign T53 = io_req_bits_in2[5'h1f:1'h0];
  assign T54 = T65 ? T64 : T55;
  assign T55 = 32'h0 - T56;
  assign T56 = {31'h0, rhs_sign};
  assign rhs_sign = T61 & T57;
  assign T57 = T60 ? T59 : T58;
  assign T58 = io_req_bits_in2[5'h1f:5'h1f];
  assign T59 = io_req_bits_in2[6'h3f:6'h3f];
  assign T60 = io_req_bits_dw == 1'h1;
  assign T61 = T62 | T18;
  assign T62 = T63 == 4'h0;
  assign T63 = io_req_bits_fn & 4'h9;
  assign T64 = io_req_bits_in2[6'h3f:6'h20];
  assign T65 = io_req_bits_dw == 1'h1;
  assign T66 = remainder[8'h80:7'h40];
  assign T67 = count == 7'h0;
  assign T68 = T1 ? 7'h0 : T69;
  assign T69 = T75 ? T74 : T70;
  assign T70 = T72 ? T71 : count;
  assign T71 = count + 7'h1;
  assign T72 = T73 & isMul;
  assign T73 = state == 3'h2;
  assign T74 = count + 7'h1;
  assign T75 = T77 & T76;
  assign T76 = isMul ^ 1'h1;
  assign T77 = state == 3'h2;
  assign T78 = T89 & T79;
  assign T79 = T38 ? lhs_sign : T80;
  assign T80 = lhs_sign != rhs_sign;
  assign lhs_sign = T85 & T81;
  assign T81 = T84 ? T83 : T82;
  assign T82 = io_req_bits_in1[5'h1f:5'h1f];
  assign T83 = io_req_bits_in1[6'h3f:6'h3f];
  assign T84 = io_req_bits_dw == 1'h1;
  assign T85 = T88 | T86;
  assign T86 = T87 == 4'h0;
  assign T87 = io_req_bits_fn & 4'h3;
  assign T88 = T62 | T18;
  assign T89 = T15 ^ 1'h1;
  assign T90 = state == 3'h3;
  assign T91 = isHi ? 3'h3 : 3'h5;
  assign T92 = T72 & T93;
  assign T93 = count == 7'h3f;
  assign T94 = isHi ? 3'h3 : T95;
  assign T95 = neg_out ? 3'h4 : 3'h5;
  assign T96 = T75 & T97;
  assign T97 = count == 7'h40;
  assign T98 = T99 | io_kill;
  assign T99 = io_resp_ready & io_resp_valid;
  assign T100 = T101 ? 3'h1 : 3'h2;
  assign T101 = lhs_sign | T102;
  assign T102 = rhs_sign & T103;
  assign T103 = T15 ^ 1'h1;
  assign T104 = {66'h0, negated_remainder};
  assign T105 = {66'h0, T106};
  assign T106 = remainder[8'h80:7'h41];
  assign T107 = T108;
  assign T108 = {T131, T109};
  assign T109 = {1'h0, T110};
  assign T110 = T111[6'h3f:1'h0];
  assign T111 = {T130, T112};
  assign T112 = T113[6'h3f:1'h0];
  assign T113 = T114;
  assign T114 = {T120, T115};
  assign T115 = T116[6'h3f:1'h1];
  assign T116 = T117[6'h3f:1'h0];
  assign T117 = {T119, T118};
  assign T118 = remainder[6'h3f:1'h0];
  assign T119 = remainder[8'h81:7'h41];
  assign T120 = T125 + T121;
  assign T121 = {T124, T122};
  assign T122 = T123;
  assign T123 = T117[8'h80:7'h40];
  assign T124 = T122[7'h40:7'h40];
  assign T125 = $signed(T129) * $signed(T126);
  assign T126 = T127;
  assign T127 = {1'h0, T128};
  assign T128 = T116[1'h0:1'h0];
  assign T129 = divisor;
  assign T130 = T113[8'h80:7'h40];
  assign T131 = T111 >> 7'h40;
  assign T132 = {1'h0, T133};
  assign T133 = {T137, T134};
  assign T134 = {T136, T135};
  assign T135 = T46 ^ 1'h1;
  assign T136 = remainder[6'h3f:1'h0];
  assign T137 = T46 ? T139 : T138;
  assign T138 = subtractor[6'h3f:1'h0];
  assign T139 = remainder[7'h7f:7'h40];
  assign T140 = {66'h0, lhs_in};
  assign lhs_in = {T142, T141};
  assign T141 = io_req_bits_in1[5'h1f:1'h0];
  assign T142 = T146 ? T145 : T143;
  assign T143 = 32'h0 - T144;
  assign T144 = {31'h0, lhs_sign};
  assign T145 = io_req_bits_in1[6'h3f:6'h20];
  assign T146 = io_req_bits_dw == 1'h1;
  assign T147 = {T149, T148};
  assign T148 = remainder[5'h1f:1'h0];
  assign T149 = 32'h0 - T150;
  assign T150 = {31'h0, T151};
  assign T151 = remainder[5'h1f:5'h1f];
  assign T152 = req_dw == 1'h0;
  assign T153 = T1 ? io_req_bits_dw : req_dw;
  assign io_resp_valid = T154;
  assign T154 = state == 3'h5;
  assign io_req_ready = T155;
  assign T155 = state == 3'h0;

  always @(posedge clk) begin
    if(T1) begin
      req_tag <= io_req_bits_tag;
    end
    if(T1) begin
      remainder <= T140;
    end else if(T75) begin
      remainder <= T132;
    end else if(T72) begin
      remainder <= T107;
    end else if(T90) begin
      remainder <= T105;
    end else if(T30) begin
      remainder <= T104;
    end else if(T12) begin
      remainder <= T10;
    end
    if(T1) begin
      isMul <= T15;
    end
    if(reset) begin
      state <= 3'h0;
    end else if(T1) begin
      state <= T100;
    end else if(T98) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= T94;
    end else if(T92) begin
      state <= T91;
    end else if(T90) begin
      state <= T31;
    end else if(T30) begin
      state <= 3'h5;
    end else if(T21) begin
      state <= 3'h2;
    end
    if(T1) begin
      neg_out <= T78;
    end else if(T34) begin
      neg_out <= 1'h0;
    end
    if(T1) begin
      isHi <= T38;
    end
    if(T1) begin
      divisor <= T52;
    end else if(T49) begin
      divisor <= subtractor;
    end
    if(T1) begin
      count <= 7'h0;
    end else if(T75) begin
      count <= T74;
    end else if(T72) begin
      count <= T71;
    end
    if(T1) begin
      req_dw <= io_req_bits_dw;
    end
  end
endmodule

module CSRFile(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [11:0] io_rw_addr,
    input [1:0] io_rw_cmd,
    output[63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    output[7:0] io_status_ip,
    output[7:0] io_status_im,
    output[6:0] io_status_zero,
    output io_status_er,
    output io_status_vm,
    output io_status_s64,
    output io_status_u64,
    output io_status_ef,
    output io_status_pei,
    output io_status_ei,
    output io_status_ps,
    output io_status_s,
    output[31:0] io_ptbr,
    output[43:0] io_evec,
    input  io_exception,
    input  io_retire,
    input  io_uarch_counters_15,
    input  io_uarch_counters_14,
    input  io_uarch_counters_13,
    input  io_uarch_counters_12,
    input  io_uarch_counters_11,
    input  io_uarch_counters_10,
    input  io_uarch_counters_9,
    input  io_uarch_counters_8,
    input  io_uarch_counters_7,
    input  io_uarch_counters_6,
    input  io_uarch_counters_5,
    input  io_uarch_counters_4,
    input  io_uarch_counters_3,
    input  io_uarch_counters_2,
    input  io_uarch_counters_1,
    input  io_uarch_counters_0,
    input [63:0] io_cause,
    input  io_badvaddr_wen,
    input [43:0] io_pc,
    input  io_sret,
    output io_fatc,
    output io_replay,
    output[63:0] io_time,
    output[2:0] io_fcsr_rm,
    input  io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    //output[6:0] io_rocc_cmd_bits_inst_funct
    //output[4:0] io_rocc_cmd_bits_inst_rs2
    //output[4:0] io_rocc_cmd_bits_inst_rs1
    //output io_rocc_cmd_bits_inst_xd
    //output io_rocc_cmd_bits_inst_xs1
    //output io_rocc_cmd_bits_inst_xs2
    //output[4:0] io_rocc_cmd_bits_inst_rd
    //output[6:0] io_rocc_cmd_bits_inst_opcode
    //output[63:0] io_rocc_cmd_bits_rs1
    //output[63:0] io_rocc_cmd_bits_rs2
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  reg [2:0] reg_frm;
  wire[2:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] wdata;
  reg [63:0] host_pcr_bits_data;
  wire[63:0] T4;
  wire[63:0] T5;
  wire T6;
  wire host_pcr_req_fire;
  wire T7;
  wire T8;
  reg  host_pcr_req_valid;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  reg [41:0] T13;
  wire[11:0] addr;
  wire[11:0] T15;
  wire[10:0] T16;
  wire[10:0] T17;
  reg [4:0] host_pcr_bits_addr;
  wire[4:0] T18;
  wire wen;
  wire T19;
  reg  host_pcr_bits_rw;
  wire T20;
  wire[63:0] T21;
  wire[58:0] T22;
  wire T23;
  wire T24;
  wire[63:0] T25;
  reg [5:0] R26;
  wire[5:0] T27;
  wire[5:0] T28;
  wire[5:0] T29;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[5:0] T32;
  wire[63:0] T33;
  wire T34;
  wire T35;
  reg [57:0] R36;
  wire[57:0] T37;
  wire[57:0] T38;
  wire[57:0] T39;
  wire[57:0] T40;
  wire T41;
  wire[57:0] T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[43:0] T47;
  wire[43:0] T48;
  reg [43:0] reg_epc;
  wire[43:0] T49;
  wire[43:0] T50;
  wire[43:0] T51;
  wire[43:0] T52;
  wire[43:0] T53;
  wire T54;
  wire T55;
  wire[43:0] T56;
  wire[42:0] T57;
  reg [42:0] reg_evec;
  wire[42:0] T58;
  wire[42:0] T59;
  wire[42:0] T60;
  wire T61;
  wire T62;
  wire T63;
  reg [31:0] reg_ptbr;
  wire[31:0] T64;
  wire[31:0] T65;
  wire[31:0] T66;
  wire[18:0] T67;
  wire T68;
  wire T69;
  reg  reg_status_s;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  reg  reg_status_ps;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  reg  reg_status_ei;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  reg  reg_status_pei;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg  reg_status_ef;
  wire T90;
  wire T91;
  wire T92;
  reg  reg_status_u64;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  reg  reg_status_s64;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg  reg_status_vm;
  wire T101;
  wire T102;
  wire T103;
  reg  reg_status_er;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  reg [6:0] reg_status_zero;
  wire[6:0] T108;
  wire[6:0] T109;
  wire[6:0] T110;
  wire[6:0] T111;
  reg [7:0] reg_status_im;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[3:0] T116;
  wire[1:0] T117;
  reg  r_irq_ipi;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire[1:0] T124;
  wire T125;
  reg [63:0] reg_fromhost;
  wire[63:0] T126;
  wire[63:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  reg  r_irq_timer;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  reg [31:0] reg_compare;
  wire[31:0] T138;
  wire[31:0] T139;
  wire[31:0] T140;
  wire T141;
  wire T142;
  wire[31:0] T143;
  wire[63:0] T144;
  wire[63:0] T145;
  wire[63:0] T146;
  reg [5:0] R147;
  wire[5:0] T148;
  wire[5:0] T149;
  wire[5:0] T150;
  wire[6:0] T151;
  wire[6:0] T152;
  wire T153;
  reg [57:0] R154;
  wire[57:0] T155;
  wire[57:0] T156;
  wire[57:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[63:0] T161;
  wire[63:0] T162;
  wire[63:0] T163;
  reg [5:0] R164;
  wire[5:0] T165;
  wire[5:0] T166;
  wire[5:0] T167;
  wire[6:0] T168;
  wire[6:0] T169;
  wire T170;
  reg [57:0] R171;
  wire[57:0] T172;
  wire[57:0] T173;
  wire[57:0] T174;
  wire T175;
  wire T176;
  wire T177;
  wire[63:0] T178;
  wire[63:0] T179;
  wire[63:0] T180;
  reg [5:0] R181;
  wire[5:0] T182;
  wire[5:0] T183;
  wire[5:0] T184;
  wire[6:0] T185;
  wire[6:0] T186;
  wire T187;
  reg [57:0] R188;
  wire[57:0] T189;
  wire[57:0] T190;
  wire[57:0] T191;
  wire T192;
  wire T193;
  wire T194;
  wire[63:0] T195;
  wire[63:0] T196;
  wire[63:0] T197;
  reg [5:0] R198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[6:0] T202;
  wire[6:0] T203;
  wire T204;
  reg [57:0] R205;
  wire[57:0] T206;
  wire[57:0] T207;
  wire[57:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire[63:0] T212;
  wire[63:0] T213;
  wire[63:0] T214;
  reg [5:0] R215;
  wire[5:0] T216;
  wire[5:0] T217;
  wire[5:0] T218;
  wire[6:0] T219;
  wire[6:0] T220;
  wire T221;
  reg [57:0] R222;
  wire[57:0] T223;
  wire[57:0] T224;
  wire[57:0] T225;
  wire T226;
  wire T227;
  wire T228;
  wire[63:0] T229;
  wire[63:0] T230;
  wire[63:0] T231;
  reg [5:0] R232;
  wire[5:0] T233;
  wire[5:0] T234;
  wire[5:0] T235;
  wire[6:0] T236;
  wire[6:0] T237;
  wire T238;
  reg [57:0] R239;
  wire[57:0] T240;
  wire[57:0] T241;
  wire[57:0] T242;
  wire T243;
  wire T244;
  wire T245;
  wire[63:0] T246;
  wire[63:0] T247;
  wire[63:0] T248;
  reg [5:0] R249;
  wire[5:0] T250;
  wire[5:0] T251;
  wire[5:0] T252;
  wire[6:0] T253;
  wire[6:0] T254;
  wire T255;
  reg [57:0] R256;
  wire[57:0] T257;
  wire[57:0] T258;
  wire[57:0] T259;
  wire T260;
  wire T261;
  wire T262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire[63:0] T265;
  reg [5:0] R266;
  wire[5:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[6:0] T270;
  wire[6:0] T271;
  wire T272;
  reg [57:0] R273;
  wire[57:0] T274;
  wire[57:0] T275;
  wire[57:0] T276;
  wire T277;
  wire T278;
  wire T279;
  wire[63:0] T280;
  wire[63:0] T281;
  wire[63:0] T282;
  reg [5:0] R283;
  wire[5:0] T284;
  wire[5:0] T285;
  wire[5:0] T286;
  wire[6:0] T287;
  wire[6:0] T288;
  wire T289;
  reg [57:0] R290;
  wire[57:0] T291;
  wire[57:0] T292;
  wire[57:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[63:0] T297;
  wire[63:0] T298;
  wire[63:0] T299;
  reg [5:0] R300;
  wire[5:0] T301;
  wire[5:0] T302;
  wire[5:0] T303;
  wire[6:0] T304;
  wire[6:0] T305;
  wire T306;
  reg [57:0] R307;
  wire[57:0] T308;
  wire[57:0] T309;
  wire[57:0] T310;
  wire T311;
  wire T312;
  wire T313;
  wire[63:0] T314;
  wire[63:0] T315;
  wire[63:0] T316;
  reg [5:0] R317;
  wire[5:0] T318;
  wire[5:0] T319;
  wire[5:0] T320;
  wire[6:0] T321;
  wire[6:0] T322;
  wire T323;
  reg [57:0] R324;
  wire[57:0] T325;
  wire[57:0] T326;
  wire[57:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[63:0] T331;
  wire[63:0] T332;
  wire[63:0] T333;
  reg [5:0] R334;
  wire[5:0] T335;
  wire[5:0] T336;
  wire[5:0] T337;
  wire[6:0] T338;
  wire[6:0] T339;
  wire T340;
  reg [57:0] R341;
  wire[57:0] T342;
  wire[57:0] T343;
  wire[57:0] T344;
  wire T345;
  wire T346;
  wire T347;
  wire[63:0] T348;
  wire[63:0] T349;
  wire[63:0] T350;
  reg [5:0] R351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[6:0] T355;
  wire[6:0] T356;
  wire T357;
  reg [57:0] R358;
  wire[57:0] T359;
  wire[57:0] T360;
  wire[57:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire[63:0] T365;
  wire[63:0] T366;
  wire[63:0] T367;
  reg [5:0] R368;
  wire[5:0] T369;
  wire[5:0] T370;
  wire[5:0] T371;
  wire[6:0] T372;
  wire[6:0] T373;
  wire T374;
  reg [57:0] R375;
  wire[57:0] T376;
  wire[57:0] T377;
  wire[57:0] T378;
  wire T379;
  wire T380;
  wire T381;
  wire[63:0] T382;
  wire[63:0] T383;
  wire[63:0] T384;
  reg [5:0] R385;
  wire[5:0] T386;
  wire[5:0] T387;
  wire[5:0] T388;
  wire[6:0] T389;
  wire[6:0] T390;
  wire T391;
  reg [57:0] R392;
  wire[57:0] T393;
  wire[57:0] T394;
  wire[57:0] T395;
  wire T396;
  wire T397;
  wire T398;
  wire[63:0] T399;
  wire[63:0] T400;
  wire[63:0] T401;
  reg [5:0] R402;
  wire[5:0] T403;
  wire[5:0] T404;
  wire[5:0] T405;
  wire[6:0] T406;
  wire[6:0] T407;
  wire T408;
  reg [57:0] R409;
  wire[57:0] T410;
  wire[57:0] T411;
  wire[57:0] T412;
  wire T413;
  wire T414;
  wire T415;
  wire[63:0] T416;
  wire[63:0] T417;
  wire[63:0] T418;
  wire[63:0] T419;
  reg [63:0] reg_tohost;
  wire[63:0] T420;
  wire[63:0] T421;
  wire[63:0] T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire[63:0] T431;
  wire[63:0] T432;
  wire T433;
  reg  reg_stats;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire[63:0] T439;
  wire[63:0] T440;
  wire[1:0] T441;
  wire[63:0] T442;
  wire[63:0] T443;
  wire[1:0] T444;
  wire T445;
  wire[63:0] T446;
  wire[63:0] T447;
  wire[1:0] T448;
  wire[63:0] T449;
  wire[63:0] T450;
  wire[1:0] T451;
  wire T452;
  wire[63:0] T453;
  wire[63:0] T454;
  wire T455;
  wire T456;
  wire[63:0] T457;
  wire[63:0] T458;
  wire[31:0] T459;
  wire[31:0] T460;
  wire[31:0] T461;
  wire[5:0] T462;
  wire[2:0] T463;
  wire[1:0] T464;
  wire[2:0] T465;
  wire[1:0] T466;
  wire[25:0] T467;
  wire[2:0] T468;
  wire[1:0] T469;
  wire[22:0] T470;
  wire[14:0] T471;
  wire[63:0] T472;
  wire[63:0] T473;
  reg [63:0] reg_cause;
  wire[63:0] T474;
  wire T475;
  wire[63:0] T476;
  wire[63:0] T477;
  wire[42:0] T478;
  wire[63:0] T479;
  wire[63:0] T480;
  wire[31:0] T481;
  wire[63:0] T482;
  wire[63:0] T483;
  wire[63:0] T484;
  wire[63:0] T485;
  wire[63:0] T486;
  wire[31:0] T487;
  wire[31:0] read_ptbr;
  wire[18:0] T488;
  wire[63:0] T489;
  wire[63:0] T490;
  wire[42:0] T491;
  reg [42:0] reg_badvaddr;
  wire[42:0] T492;
  wire[43:0] T493;
  wire[43:0] T494;
  wire[43:0] T495;
  wire[43:0] T496;
  wire[42:0] T497;
  wire T498;
  wire T499;
  wire[20:0] T500;
  wire T501;
  wire T502;
  wire[42:0] T503;
  wire T504;
  wire[63:0] T505;
  wire[63:0] T506;
  wire[43:0] T507;
  wire[63:0] T508;
  wire[63:0] T509;
  reg [63:0] reg_sup1;
  wire[63:0] T510;
  wire T511;
  wire T512;
  wire[63:0] T513;
  wire[63:0] T514;
  reg [63:0] reg_sup0;
  wire[63:0] T515;
  wire T516;
  wire T517;
  wire[63:0] T518;
  wire[63:0] T519;
  wire[63:0] T520;
  reg [5:0] R521;
  wire[5:0] T522;
  wire[5:0] T523;
  wire[5:0] T524;
  wire[6:0] T525;
  wire[6:0] T526;
  wire T527;
  reg [57:0] R528;
  wire[57:0] T529;
  wire[57:0] T530;
  wire[57:0] T531;
  wire T532;
  wire T533;
  wire T534;
  wire[63:0] T535;
  wire[63:0] T536;
  wire T537;
  wire[63:0] T538;
  wire[63:0] T539;
  wire T540;
  wire[63:0] T541;
  wire[7:0] T542;
  wire[7:0] T543;
  wire[7:0] T544;
  reg [4:0] reg_fflags;
  wire[4:0] T545;
  wire[63:0] T546;
  wire[63:0] T547;
  wire[63:0] T548;
  wire[4:0] T549;
  wire[4:0] T550;
  wire T551;
  wire T552;
  wire[7:0] T553;
  wire[4:0] T554;
  wire[4:0] T555;
  wire[2:0] T556;
  wire[4:0] T557;
  wire T558;
  wire T559;
  reg  host_pcr_rep_valid;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    reg_frm = {1{$random}};
    host_pcr_bits_data = {2{$random}};
    host_pcr_req_valid = {1{$random}};
    host_pcr_bits_addr = {1{$random}};
    host_pcr_bits_rw = {1{$random}};
    R26 = {1{$random}};
    R36 = {2{$random}};
    reg_epc = {2{$random}};
    reg_evec = {2{$random}};
    reg_ptbr = {1{$random}};
    reg_status_s = {1{$random}};
    reg_status_ps = {1{$random}};
    reg_status_ei = {1{$random}};
    reg_status_pei = {1{$random}};
    reg_status_ef = {1{$random}};
    reg_status_u64 = {1{$random}};
    reg_status_s64 = {1{$random}};
    reg_status_vm = {1{$random}};
    reg_status_er = {1{$random}};
    reg_status_zero = {1{$random}};
    reg_status_im = {1{$random}};
    r_irq_ipi = {1{$random}};
    reg_fromhost = {2{$random}};
    r_irq_timer = {1{$random}};
    reg_compare = {1{$random}};
    R147 = {1{$random}};
    R154 = {2{$random}};
    R164 = {1{$random}};
    R171 = {2{$random}};
    R181 = {1{$random}};
    R188 = {2{$random}};
    R198 = {1{$random}};
    R205 = {2{$random}};
    R215 = {1{$random}};
    R222 = {2{$random}};
    R232 = {1{$random}};
    R239 = {2{$random}};
    R249 = {1{$random}};
    R256 = {2{$random}};
    R266 = {1{$random}};
    R273 = {2{$random}};
    R283 = {1{$random}};
    R290 = {2{$random}};
    R300 = {1{$random}};
    R307 = {2{$random}};
    R317 = {1{$random}};
    R324 = {2{$random}};
    R334 = {1{$random}};
    R341 = {2{$random}};
    R351 = {1{$random}};
    R358 = {2{$random}};
    R368 = {1{$random}};
    R375 = {2{$random}};
    R385 = {1{$random}};
    R392 = {2{$random}};
    R402 = {1{$random}};
    R409 = {2{$random}};
    reg_tohost = {2{$random}};
    reg_stats = {1{$random}};
    reg_cause = {2{$random}};
    reg_badvaddr = {2{$random}};
    reg_sup1 = {2{$random}};
    reg_sup0 = {2{$random}};
    R521 = {1{$random}};
    R528 = {2{$random}};
    reg_fflags = {1{$random}};
    host_pcr_rep_valid = {1{$random}};
  end
`endif

  assign io_fcsr_rm = reg_frm;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = T23 ? T21 : T2;
  assign T2 = T11 ? wdata : T3;
  assign T3 = {61'h0, reg_frm};
  assign wdata = T8 ? io_rw_wdata : host_pcr_bits_data;
  assign T4 = host_pcr_req_fire ? io_rw_rdata : T5;
  assign T5 = T6 ? io_host_pcr_req_bits_data : host_pcr_bits_data;
  assign T6 = io_host_pcr_req_ready & io_host_pcr_req_valid;
  assign host_pcr_req_fire = host_pcr_req_valid & T7;
  assign T7 = T8 ^ 1'h1;
  assign T8 = io_rw_cmd != 2'h0;
  assign T9 = host_pcr_req_fire ? 1'h0 : T10;
  assign T10 = T6 ? 1'h1 : host_pcr_req_valid;
  assign T11 = wen & T12;
  assign T12 = T13[1'h1:1'h1];
  always @(*) case (addr)
    1: T13 = 42'h1;
    2: T13 = 42'h2;
    3: T13 = 42'h4;
    192: T13 = 42'h8;
    1280: T13 = 42'h10;
    1281: T13 = 42'h20;
    1282: T13 = 42'h40;
    1283: T13 = 42'h80;
    1284: T13 = 42'h100;
    1285: T13 = 42'h200;
    1286: T13 = 42'h400;
    1287: T13 = 42'h800;
    1288: T13 = 42'h1000;
    1289: T13 = 42'h2000;
    1290: T13 = 42'h4000;
    1291: T13 = 42'h8000;
    1292: T13 = 42'h10000;
    1293: T13 = 42'h20000;
    1294: T13 = 42'h40000;
    1295: T13 = 42'h80000;
    1309: T13 = 42'h100000;
    1310: T13 = 42'h200000;
    1311: T13 = 42'h400000;
    3072: T13 = 42'h800000;
    3073: T13 = 42'h1000000;
    3074: T13 = 42'h2000000;
    3264: T13 = 42'h4000000;
    3265: T13 = 42'h8000000;
    3266: T13 = 42'h10000000;
    3267: T13 = 42'h20000000;
    3268: T13 = 42'h40000000;
    3269: T13 = 42'h80000000;
    3270: T13 = 42'h100000000;
    3271: T13 = 42'h200000000;
    3272: T13 = 42'h400000000;
    3273: T13 = 42'h800000000;
    3274: T13 = 42'h1000000000;
    3275: T13 = 42'h2000000000;
    3276: T13 = 42'h4000000000;
    3277: T13 = 42'h8000000000;
    3278: T13 = 42'h10000000000;
    3279: T13 = 42'h20000000000;
`ifndef SYNTHESIS
    default: T13 = {2{$random}};
`else
    default: T13 = 42'bx;
`endif
  endcase
  assign addr = T8 ? io_rw_addr : T15;
  assign T15 = {1'h0, T16};
  assign T16 = T17 | 11'h500;
  assign T17 = {6'h0, host_pcr_bits_addr};
  assign T18 = T6 ? io_host_pcr_req_bits_addr : host_pcr_bits_addr;
  assign wen = T8 | T19;
  assign T19 = host_pcr_req_fire & host_pcr_bits_rw;
  assign T20 = T6 ? io_host_pcr_req_bits_rw : host_pcr_bits_rw;
  assign T21 = {5'h0, T22};
  assign T22 = wdata >> 3'h5;
  assign T23 = wen & T24;
  assign T24 = T13[2'h2:2'h2];
  assign io_time = T25;
  assign T25 = {R36, R26};
  assign T27 = reset ? 6'h0 : T28;
  assign T28 = T34 ? T32 : T29;
  assign T29 = T30[3'h5:1'h0];
  assign T30 = T31 + 7'h1;
  assign T31 = {1'h0, R26};
  assign T32 = T33[3'h5:1'h0];
  assign T33 = wdata;
  assign T34 = wen & T35;
  assign T35 = T13[4'ha:4'ha];
  assign T37 = reset ? 58'h0 : T38;
  assign T38 = T34 ? T42 : T39;
  assign T39 = T41 ? T40 : R36;
  assign T40 = R36 + 58'h1;
  assign T41 = T30[3'h6:3'h6];
  assign T42 = T33[6'h3f:3'h6];
  assign io_replay = T43;
  assign T43 = io_host_ipi_req_valid & T44;
  assign T44 = io_host_ipi_req_ready ^ 1'h1;
  assign io_fatc = T45;
  assign T45 = wen & T46;
  assign T46 = T13[5'h11:5'h11];
  assign io_evec = T47;
  assign T47 = T48;
  assign T48 = io_exception ? T56 : reg_epc;
  assign T49 = T54 ? T52 : T50;
  assign T50 = io_exception ? T51 : reg_epc;
  assign T51 = io_pc;
  assign T52 = T53;
  assign T53 = wdata[6'h2b:1'h0];
  assign T54 = wen & T55;
  assign T55 = T13[3'h6:3'h6];
  assign T56 = {T63, T57};
  assign T57 = reg_evec;
  assign T58 = T61 ? T59 : reg_evec;
  assign T59 = T60;
  assign T60 = wdata[6'h2a:1'h0];
  assign T61 = wen & T62;
  assign T62 = T13[4'hc:4'hc];
  assign T63 = T57[6'h2a:6'h2a];
  assign io_ptbr = reg_ptbr;
  assign T64 = T68 ? T65 : reg_ptbr;
  assign T65 = T66;
  assign T66 = {T67, 13'h0};
  assign T67 = wdata[5'h1f:4'hd];
  assign T68 = wen & T69;
  assign T69 = T13[4'h8:4'h8];
  assign io_status_s = reg_status_s;
  assign T70 = reset ? 1'h1 : T71;
  assign T71 = T78 ? T80 : T72;
  assign T72 = io_sret ? reg_status_ps : T73;
  assign T73 = io_exception ? 1'h1 : reg_status_s;
  assign T74 = reset ? 1'h0 : T75;
  assign T75 = T78 ? T77 : T76;
  assign T76 = io_exception ? reg_status_s : reg_status_ps;
  assign T77 = wdata[1'h1:1'h1];
  assign T78 = wen & T79;
  assign T79 = T13[4'he:4'he];
  assign T80 = wdata[1'h0:1'h0];
  assign io_status_ps = reg_status_ps;
  assign io_status_ei = reg_status_ei;
  assign T81 = reset ? 1'h0 : T82;
  assign T82 = T78 ? T89 : T83;
  assign T83 = io_sret ? reg_status_pei : T84;
  assign T84 = io_exception ? 1'h0 : reg_status_ei;
  assign T85 = reset ? 1'h0 : T86;
  assign T86 = T78 ? T88 : T87;
  assign T87 = io_exception ? reg_status_ei : reg_status_pei;
  assign T88 = wdata[2'h3:2'h3];
  assign T89 = wdata[2'h2:2'h2];
  assign io_status_pei = reg_status_pei;
  assign io_status_ef = reg_status_ef;
  assign T90 = reset ? 1'h0 : T91;
  assign T91 = T78 ? T92 : reg_status_ef;
  assign T92 = wdata[3'h4:3'h4];
  assign io_status_u64 = reg_status_u64;
  assign T93 = reset ? 1'h1 : T94;
  assign T94 = T78 ? 1'h1 : T95;
  assign T95 = T78 ? T96 : reg_status_u64;
  assign T96 = wdata[3'h5:3'h5];
  assign io_status_s64 = reg_status_s64;
  assign T97 = reset ? 1'h1 : T98;
  assign T98 = T78 ? 1'h1 : T99;
  assign T99 = T78 ? T100 : reg_status_s64;
  assign T100 = wdata[3'h6:3'h6];
  assign io_status_vm = reg_status_vm;
  assign T101 = reset ? 1'h0 : T102;
  assign T102 = T78 ? T103 : reg_status_vm;
  assign T103 = wdata[3'h7:3'h7];
  assign io_status_er = reg_status_er;
  assign T104 = reset ? 1'h0 : T105;
  assign T105 = T78 ? 1'h0 : T106;
  assign T106 = T78 ? T107 : reg_status_er;
  assign T107 = wdata[4'h8:4'h8];
  assign io_status_zero = reg_status_zero;
  assign T108 = reset ? 7'h0 : T109;
  assign T109 = T78 ? 7'h0 : T110;
  assign T110 = T78 ? T111 : reg_status_zero;
  assign T111 = wdata[4'hf:4'h9];
  assign io_status_im = reg_status_im;
  assign T112 = reset ? 8'h0 : T113;
  assign T113 = T78 ? T114 : reg_status_im;
  assign T114 = wdata[5'h17:5'h10];
  assign io_status_ip = T115;
  assign T115 = {T116, 4'h0};
  assign T116 = {T124, T117};
  assign T117 = {r_irq_ipi, 1'h0};
  assign T118 = reset ? 1'h1 : T119;
  assign T119 = io_host_ipi_rep_valid ? 1'h1 : T120;
  assign T120 = T122 ? T121 : r_irq_ipi;
  assign T121 = wdata[1'h0:1'h0];
  assign T122 = wen & T123;
  assign T123 = T13[5'h13:5'h13];
  assign T124 = {r_irq_timer, T125};
  assign T125 = reg_fromhost != 64'h0;
  assign T126 = reset ? 64'h0 : T127;
  assign T127 = T128 ? wdata : reg_fromhost;
  assign T128 = T132 & T129;
  assign T129 = T131 | T130;
  assign T130 = host_pcr_req_fire ^ 1'h1;
  assign T131 = reg_fromhost == 64'h0;
  assign T132 = wen & T133;
  assign T133 = T13[5'h16:5'h16];
  assign T134 = reset ? 1'h0 : T135;
  assign T135 = T141 ? 1'h0 : T136;
  assign T136 = T137 ? 1'h1 : r_irq_timer;
  assign T137 = T143 == reg_compare;
  assign T138 = T141 ? T139 : reg_compare;
  assign T139 = T140;
  assign T140 = wdata[5'h1f:1'h0];
  assign T141 = wen & T142;
  assign T142 = T13[4'hb:4'hb];
  assign T143 = T25[5'h1f:1'h0];
  assign io_rw_rdata = T144;
  assign T144 = T161 | T145;
  assign T145 = T160 ? T146 : 64'h0;
  assign T146 = {R154, R147};
  assign T148 = reset ? 6'h0 : T149;
  assign T149 = T153 ? T150 : R147;
  assign T150 = T151[3'h5:1'h0];
  assign T151 = T152 + 7'h1;
  assign T152 = {1'h0, R147};
  assign T153 = io_uarch_counters_15 != 1'h0;
  assign T155 = reset ? 58'h0 : T156;
  assign T156 = T158 ? T157 : R154;
  assign T157 = R154 + 58'h1;
  assign T158 = T153 & T159;
  assign T159 = T151[3'h6:3'h6];
  assign T160 = T13[6'h29:6'h29];
  assign T161 = T178 | T162;
  assign T162 = T177 ? T163 : 64'h0;
  assign T163 = {R171, R164};
  assign T165 = reset ? 6'h0 : T166;
  assign T166 = T170 ? T167 : R164;
  assign T167 = T168[3'h5:1'h0];
  assign T168 = T169 + 7'h1;
  assign T169 = {1'h0, R164};
  assign T170 = io_uarch_counters_14 != 1'h0;
  assign T172 = reset ? 58'h0 : T173;
  assign T173 = T175 ? T174 : R171;
  assign T174 = R171 + 58'h1;
  assign T175 = T170 & T176;
  assign T176 = T168[3'h6:3'h6];
  assign T177 = T13[6'h28:6'h28];
  assign T178 = T195 | T179;
  assign T179 = T194 ? T180 : 64'h0;
  assign T180 = {R188, R181};
  assign T182 = reset ? 6'h0 : T183;
  assign T183 = T187 ? T184 : R181;
  assign T184 = T185[3'h5:1'h0];
  assign T185 = T186 + 7'h1;
  assign T186 = {1'h0, R181};
  assign T187 = io_uarch_counters_13 != 1'h0;
  assign T189 = reset ? 58'h0 : T190;
  assign T190 = T192 ? T191 : R188;
  assign T191 = R188 + 58'h1;
  assign T192 = T187 & T193;
  assign T193 = T185[3'h6:3'h6];
  assign T194 = T13[6'h27:6'h27];
  assign T195 = T212 | T196;
  assign T196 = T211 ? T197 : 64'h0;
  assign T197 = {R205, R198};
  assign T199 = reset ? 6'h0 : T200;
  assign T200 = T204 ? T201 : R198;
  assign T201 = T202[3'h5:1'h0];
  assign T202 = T203 + 7'h1;
  assign T203 = {1'h0, R198};
  assign T204 = io_uarch_counters_12 != 1'h0;
  assign T206 = reset ? 58'h0 : T207;
  assign T207 = T209 ? T208 : R205;
  assign T208 = R205 + 58'h1;
  assign T209 = T204 & T210;
  assign T210 = T202[3'h6:3'h6];
  assign T211 = T13[6'h26:6'h26];
  assign T212 = T229 | T213;
  assign T213 = T228 ? T214 : 64'h0;
  assign T214 = {R222, R215};
  assign T216 = reset ? 6'h0 : T217;
  assign T217 = T221 ? T218 : R215;
  assign T218 = T219[3'h5:1'h0];
  assign T219 = T220 + 7'h1;
  assign T220 = {1'h0, R215};
  assign T221 = io_uarch_counters_11 != 1'h0;
  assign T223 = reset ? 58'h0 : T224;
  assign T224 = T226 ? T225 : R222;
  assign T225 = R222 + 58'h1;
  assign T226 = T221 & T227;
  assign T227 = T219[3'h6:3'h6];
  assign T228 = T13[6'h25:6'h25];
  assign T229 = T246 | T230;
  assign T230 = T245 ? T231 : 64'h0;
  assign T231 = {R239, R232};
  assign T233 = reset ? 6'h0 : T234;
  assign T234 = T238 ? T235 : R232;
  assign T235 = T236[3'h5:1'h0];
  assign T236 = T237 + 7'h1;
  assign T237 = {1'h0, R232};
  assign T238 = io_uarch_counters_10 != 1'h0;
  assign T240 = reset ? 58'h0 : T241;
  assign T241 = T243 ? T242 : R239;
  assign T242 = R239 + 58'h1;
  assign T243 = T238 & T244;
  assign T244 = T236[3'h6:3'h6];
  assign T245 = T13[6'h24:6'h24];
  assign T246 = T263 | T247;
  assign T247 = T262 ? T248 : 64'h0;
  assign T248 = {R256, R249};
  assign T250 = reset ? 6'h0 : T251;
  assign T251 = T255 ? T252 : R249;
  assign T252 = T253[3'h5:1'h0];
  assign T253 = T254 + 7'h1;
  assign T254 = {1'h0, R249};
  assign T255 = io_uarch_counters_9 != 1'h0;
  assign T257 = reset ? 58'h0 : T258;
  assign T258 = T260 ? T259 : R256;
  assign T259 = R256 + 58'h1;
  assign T260 = T255 & T261;
  assign T261 = T253[3'h6:3'h6];
  assign T262 = T13[6'h23:6'h23];
  assign T263 = T280 | T264;
  assign T264 = T279 ? T265 : 64'h0;
  assign T265 = {R273, R266};
  assign T267 = reset ? 6'h0 : T268;
  assign T268 = T272 ? T269 : R266;
  assign T269 = T270[3'h5:1'h0];
  assign T270 = T271 + 7'h1;
  assign T271 = {1'h0, R266};
  assign T272 = io_uarch_counters_8 != 1'h0;
  assign T274 = reset ? 58'h0 : T275;
  assign T275 = T277 ? T276 : R273;
  assign T276 = R273 + 58'h1;
  assign T277 = T272 & T278;
  assign T278 = T270[3'h6:3'h6];
  assign T279 = T13[6'h22:6'h22];
  assign T280 = T297 | T281;
  assign T281 = T296 ? T282 : 64'h0;
  assign T282 = {R290, R283};
  assign T284 = reset ? 6'h0 : T285;
  assign T285 = T289 ? T286 : R283;
  assign T286 = T287[3'h5:1'h0];
  assign T287 = T288 + 7'h1;
  assign T288 = {1'h0, R283};
  assign T289 = io_uarch_counters_7 != 1'h0;
  assign T291 = reset ? 58'h0 : T292;
  assign T292 = T294 ? T293 : R290;
  assign T293 = R290 + 58'h1;
  assign T294 = T289 & T295;
  assign T295 = T287[3'h6:3'h6];
  assign T296 = T13[6'h21:6'h21];
  assign T297 = T314 | T298;
  assign T298 = T313 ? T299 : 64'h0;
  assign T299 = {R307, R300};
  assign T301 = reset ? 6'h0 : T302;
  assign T302 = T306 ? T303 : R300;
  assign T303 = T304[3'h5:1'h0];
  assign T304 = T305 + 7'h1;
  assign T305 = {1'h0, R300};
  assign T306 = io_uarch_counters_6 != 1'h0;
  assign T308 = reset ? 58'h0 : T309;
  assign T309 = T311 ? T310 : R307;
  assign T310 = R307 + 58'h1;
  assign T311 = T306 & T312;
  assign T312 = T304[3'h6:3'h6];
  assign T313 = T13[6'h20:6'h20];
  assign T314 = T331 | T315;
  assign T315 = T330 ? T316 : 64'h0;
  assign T316 = {R324, R317};
  assign T318 = reset ? 6'h0 : T319;
  assign T319 = T323 ? T320 : R317;
  assign T320 = T321[3'h5:1'h0];
  assign T321 = T322 + 7'h1;
  assign T322 = {1'h0, R317};
  assign T323 = io_uarch_counters_5 != 1'h0;
  assign T325 = reset ? 58'h0 : T326;
  assign T326 = T328 ? T327 : R324;
  assign T327 = R324 + 58'h1;
  assign T328 = T323 & T329;
  assign T329 = T321[3'h6:3'h6];
  assign T330 = T13[5'h1f:5'h1f];
  assign T331 = T348 | T332;
  assign T332 = T347 ? T333 : 64'h0;
  assign T333 = {R341, R334};
  assign T335 = reset ? 6'h0 : T336;
  assign T336 = T340 ? T337 : R334;
  assign T337 = T338[3'h5:1'h0];
  assign T338 = T339 + 7'h1;
  assign T339 = {1'h0, R334};
  assign T340 = io_uarch_counters_4 != 1'h0;
  assign T342 = reset ? 58'h0 : T343;
  assign T343 = T345 ? T344 : R341;
  assign T344 = R341 + 58'h1;
  assign T345 = T340 & T346;
  assign T346 = T338[3'h6:3'h6];
  assign T347 = T13[5'h1e:5'h1e];
  assign T348 = T365 | T349;
  assign T349 = T364 ? T350 : 64'h0;
  assign T350 = {R358, R351};
  assign T352 = reset ? 6'h0 : T353;
  assign T353 = T357 ? T354 : R351;
  assign T354 = T355[3'h5:1'h0];
  assign T355 = T356 + 7'h1;
  assign T356 = {1'h0, R351};
  assign T357 = io_uarch_counters_3 != 1'h0;
  assign T359 = reset ? 58'h0 : T360;
  assign T360 = T362 ? T361 : R358;
  assign T361 = R358 + 58'h1;
  assign T362 = T357 & T363;
  assign T363 = T355[3'h6:3'h6];
  assign T364 = T13[5'h1d:5'h1d];
  assign T365 = T382 | T366;
  assign T366 = T381 ? T367 : 64'h0;
  assign T367 = {R375, R368};
  assign T369 = reset ? 6'h0 : T370;
  assign T370 = T374 ? T371 : R368;
  assign T371 = T372[3'h5:1'h0];
  assign T372 = T373 + 7'h1;
  assign T373 = {1'h0, R368};
  assign T374 = io_uarch_counters_2 != 1'h0;
  assign T376 = reset ? 58'h0 : T377;
  assign T377 = T379 ? T378 : R375;
  assign T378 = R375 + 58'h1;
  assign T379 = T374 & T380;
  assign T380 = T372[3'h6:3'h6];
  assign T381 = T13[5'h1c:5'h1c];
  assign T382 = T399 | T383;
  assign T383 = T398 ? T384 : 64'h0;
  assign T384 = {R392, R385};
  assign T386 = reset ? 6'h0 : T387;
  assign T387 = T391 ? T388 : R385;
  assign T388 = T389[3'h5:1'h0];
  assign T389 = T390 + 7'h1;
  assign T390 = {1'h0, R385};
  assign T391 = io_uarch_counters_1 != 1'h0;
  assign T393 = reset ? 58'h0 : T394;
  assign T394 = T396 ? T395 : R392;
  assign T395 = R392 + 58'h1;
  assign T396 = T391 & T397;
  assign T397 = T389[3'h6:3'h6];
  assign T398 = T13[5'h1b:5'h1b];
  assign T399 = T416 | T400;
  assign T400 = T415 ? T401 : 64'h0;
  assign T401 = {R409, R402};
  assign T403 = reset ? 6'h0 : T404;
  assign T404 = T408 ? T405 : R402;
  assign T405 = T406[3'h5:1'h0];
  assign T406 = T407 + 7'h1;
  assign T407 = {1'h0, R402};
  assign T408 = io_uarch_counters_0 != 1'h0;
  assign T410 = reset ? 58'h0 : T411;
  assign T411 = T413 ? T412 : R409;
  assign T412 = R409 + 58'h1;
  assign T413 = T408 & T414;
  assign T414 = T406[3'h6:3'h6];
  assign T415 = T13[5'h1a:5'h1a];
  assign T416 = T418 | T417;
  assign T417 = T133 ? reg_fromhost : 64'h0;
  assign T418 = T431 | T419;
  assign T419 = T424 ? reg_tohost : 64'h0;
  assign T420 = reset ? 64'h0 : T421;
  assign T421 = T427 ? wdata : T422;
  assign T422 = T423 ? 64'h0 : reg_tohost;
  assign T423 = T425 & T424;
  assign T424 = T13[5'h15:5'h15];
  assign T425 = host_pcr_req_fire & T426;
  assign T426 = host_pcr_bits_rw ^ 1'h1;
  assign T427 = T430 & T428;
  assign T428 = T429 | host_pcr_req_fire;
  assign T429 = reg_tohost == 64'h0;
  assign T430 = wen & T424;
  assign T431 = T439 | T432;
  assign T432 = {63'h0, T433};
  assign T433 = T438 ? reg_stats : 1'h0;
  assign T434 = reset ? 1'h0 : T435;
  assign T435 = T437 ? T436 : reg_stats;
  assign T436 = wdata[1'h0:1'h0];
  assign T437 = wen & T438;
  assign T438 = T13[2'h3:2'h3];
  assign T439 = T442 | T440;
  assign T440 = {62'h0, T441};
  assign T441 = T123 ? 2'h2 : 2'h0;
  assign T442 = T446 | T443;
  assign T443 = {62'h0, T444};
  assign T444 = T445 ? 2'h2 : 2'h0;
  assign T445 = T13[5'h12:5'h12];
  assign T446 = T449 | T447;
  assign T447 = {62'h0, T448};
  assign T448 = T46 ? 2'h2 : 2'h0;
  assign T449 = T453 | T450;
  assign T450 = {62'h0, T451};
  assign T451 = T452 ? 2'h2 : 2'h0;
  assign T452 = T13[5'h10:5'h10];
  assign T453 = T457 | T454;
  assign T454 = {63'h0, T455};
  assign T455 = T456 ? io_host_id : 1'h0;
  assign T456 = T13[4'hf:4'hf];
  assign T457 = T472 | T458;
  assign T458 = {32'h0, T459};
  assign T459 = T79 ? T460 : 32'h0;
  assign T460 = T461;
  assign T461 = {T467, T462};
  assign T462 = {T465, T463};
  assign T463 = {io_status_ei, T464};
  assign T464 = {io_status_ps, io_status_s};
  assign T465 = {io_status_u64, T466};
  assign T466 = {io_status_ef, io_status_pei};
  assign T467 = {T470, T468};
  assign T468 = {io_status_er, T469};
  assign T469 = {io_status_vm, io_status_s64};
  assign T470 = {io_status_ip, T471};
  assign T471 = {io_status_im, io_status_zero};
  assign T472 = T476 | T473;
  assign T473 = T475 ? reg_cause : 64'h0;
  assign T474 = io_exception ? io_cause : reg_cause;
  assign T475 = T13[4'hd:4'hd];
  assign T476 = T479 | T477;
  assign T477 = {21'h0, T478};
  assign T478 = T62 ? reg_evec : 43'h0;
  assign T479 = T482 | T480;
  assign T480 = {32'h0, T481};
  assign T481 = T142 ? reg_compare : 32'h0;
  assign T482 = T484 | T483;
  assign T483 = T35 ? T25 : 64'h0;
  assign T484 = T485 | 64'h0;
  assign T485 = T489 | T486;
  assign T486 = {32'h0, T487};
  assign T487 = T69 ? read_ptbr : 32'h0;
  assign read_ptbr = T488 << 4'hd;
  assign T488 = reg_ptbr[5'h1f:4'hd];
  assign T489 = T505 | T490;
  assign T490 = {21'h0, T491};
  assign T491 = T504 ? reg_badvaddr : 43'h0;
  assign T492 = T493[6'h2a:1'h0];
  assign T493 = io_badvaddr_wen ? T495 : T494;
  assign T494 = {1'h0, reg_badvaddr};
  assign T495 = T496;
  assign T496 = {T498, T497};
  assign T497 = io_rw_wdata[6'h2a:1'h0];
  assign T498 = T502 ? T501 : T499;
  assign T499 = T500 != 21'h0;
  assign T500 = io_rw_wdata[6'h3f:6'h2b];
  assign T501 = T500 == 21'h1fffff;
  assign T502 = $signed(T503) < $signed(1'h0);
  assign T503 = T497;
  assign T504 = T13[3'h7:3'h7];
  assign T505 = T508 | T506;
  assign T506 = {20'h0, T507};
  assign T507 = T55 ? reg_epc : 44'h0;
  assign T508 = T513 | T509;
  assign T509 = T512 ? reg_sup1 : 64'h0;
  assign T510 = T511 ? wdata : reg_sup1;
  assign T511 = wen & T512;
  assign T512 = T13[3'h5:3'h5];
  assign T513 = T518 | T514;
  assign T514 = T517 ? reg_sup0 : 64'h0;
  assign T515 = T516 ? wdata : reg_sup0;
  assign T516 = wen & T517;
  assign T517 = T13[3'h4:3'h4];
  assign T518 = T535 | T519;
  assign T519 = T534 ? T520 : 64'h0;
  assign T520 = {R528, R521};
  assign T522 = reset ? 6'h0 : T523;
  assign T523 = T527 ? T524 : R521;
  assign T524 = T525[3'h5:1'h0];
  assign T525 = T526 + 7'h1;
  assign T526 = {1'h0, R521};
  assign T527 = io_retire != 1'h0;
  assign T529 = reset ? 58'h0 : T530;
  assign T530 = T532 ? T531 : R528;
  assign T531 = R528 + 58'h1;
  assign T532 = T527 & T533;
  assign T533 = T525[3'h6:3'h6];
  assign T534 = T13[5'h19:5'h19];
  assign T535 = T538 | T536;
  assign T536 = T537 ? T25 : 64'h0;
  assign T537 = T13[5'h18:5'h18];
  assign T538 = T541 | T539;
  assign T539 = T540 ? T25 : 64'h0;
  assign T540 = T13[5'h17:5'h17];
  assign T541 = {56'h0, T542};
  assign T542 = T553 | T543;
  assign T543 = T24 ? T544 : 8'h0;
  assign T544 = {reg_frm, reg_fflags};
  assign T545 = T546[3'h4:1'h0];
  assign T546 = T23 ? wdata : T547;
  assign T547 = T551 ? wdata : T548;
  assign T548 = {59'h0, T549};
  assign T549 = io_fcsr_flags_valid ? T550 : reg_fflags;
  assign T550 = reg_fflags | io_fcsr_flags_bits;
  assign T551 = wen & T552;
  assign T552 = T13[1'h0:1'h0];
  assign T553 = {3'h0, T554};
  assign T554 = T557 | T555;
  assign T555 = {2'h0, T556};
  assign T556 = T12 ? reg_frm : 3'h0;
  assign T557 = T552 ? reg_fflags : 5'h0;
  assign io_host_debug_stats_pcr = reg_stats;
  assign io_host_ipi_rep_ready = 1'h1;
  assign io_host_ipi_req_bits = T558;
  assign T558 = io_rw_wdata[1'h0:1'h0];
  assign io_host_ipi_req_valid = T559;
  assign T559 = T8 & T445;
  assign io_host_pcr_rep_bits = host_pcr_bits_data;
  assign io_host_pcr_rep_valid = host_pcr_rep_valid;
  assign T560 = T562 ? 1'h0 : T561;
  assign T561 = host_pcr_req_fire ? 1'h1 : host_pcr_rep_valid;
  assign T562 = io_host_pcr_rep_ready & io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = T563;
  assign T563 = T565 & T564;
  assign T564 = host_pcr_rep_valid ^ 1'h1;
  assign T565 = host_pcr_req_valid ^ 1'h1;

  always @(posedge clk) begin
    reg_frm <= T0;
    if(host_pcr_req_fire) begin
      host_pcr_bits_data <= io_rw_rdata;
    end else if(T6) begin
      host_pcr_bits_data <= io_host_pcr_req_bits_data;
    end
    if(host_pcr_req_fire) begin
      host_pcr_req_valid <= 1'h0;
    end else if(T6) begin
      host_pcr_req_valid <= 1'h1;
    end
    if(T6) begin
      host_pcr_bits_addr <= io_host_pcr_req_bits_addr;
    end
    if(T6) begin
      host_pcr_bits_rw <= io_host_pcr_req_bits_rw;
    end
    if(reset) begin
      R26 <= 6'h0;
    end else if(T34) begin
      R26 <= T32;
    end else begin
      R26 <= T29;
    end
    if(reset) begin
      R36 <= 58'h0;
    end else if(T34) begin
      R36 <= T42;
    end else if(T41) begin
      R36 <= T40;
    end
    if(T54) begin
      reg_epc <= T52;
    end else if(io_exception) begin
      reg_epc <= T51;
    end
    if(T61) begin
      reg_evec <= T59;
    end
    if(T68) begin
      reg_ptbr <= T65;
    end
    if(reset) begin
      reg_status_s <= 1'h1;
    end else if(T78) begin
      reg_status_s <= T80;
    end else if(io_sret) begin
      reg_status_s <= reg_status_ps;
    end else if(io_exception) begin
      reg_status_s <= 1'h1;
    end
    if(reset) begin
      reg_status_ps <= 1'h0;
    end else if(T78) begin
      reg_status_ps <= T77;
    end else if(io_exception) begin
      reg_status_ps <= reg_status_s;
    end
    if(reset) begin
      reg_status_ei <= 1'h0;
    end else if(T78) begin
      reg_status_ei <= T89;
    end else if(io_sret) begin
      reg_status_ei <= reg_status_pei;
    end else if(io_exception) begin
      reg_status_ei <= 1'h0;
    end
    if(reset) begin
      reg_status_pei <= 1'h0;
    end else if(T78) begin
      reg_status_pei <= T88;
    end else if(io_exception) begin
      reg_status_pei <= reg_status_ei;
    end
    if(reset) begin
      reg_status_ef <= 1'h0;
    end else if(T78) begin
      reg_status_ef <= T92;
    end
    if(reset) begin
      reg_status_u64 <= 1'h1;
    end else if(T78) begin
      reg_status_u64 <= 1'h1;
    end else if(T78) begin
      reg_status_u64 <= T96;
    end
    if(reset) begin
      reg_status_s64 <= 1'h1;
    end else if(T78) begin
      reg_status_s64 <= 1'h1;
    end else if(T78) begin
      reg_status_s64 <= T100;
    end
    if(reset) begin
      reg_status_vm <= 1'h0;
    end else if(T78) begin
      reg_status_vm <= T103;
    end
    if(reset) begin
      reg_status_er <= 1'h0;
    end else if(T78) begin
      reg_status_er <= 1'h0;
    end else if(T78) begin
      reg_status_er <= T107;
    end
    if(reset) begin
      reg_status_zero <= 7'h0;
    end else if(T78) begin
      reg_status_zero <= 7'h0;
    end else if(T78) begin
      reg_status_zero <= T111;
    end
    if(reset) begin
      reg_status_im <= 8'h0;
    end else if(T78) begin
      reg_status_im <= T114;
    end
    if(reset) begin
      r_irq_ipi <= 1'h1;
    end else if(io_host_ipi_rep_valid) begin
      r_irq_ipi <= 1'h1;
    end else if(T122) begin
      r_irq_ipi <= T121;
    end
    if(reset) begin
      reg_fromhost <= 64'h0;
    end else if(T128) begin
      reg_fromhost <= wdata;
    end
    if(reset) begin
      r_irq_timer <= 1'h0;
    end else if(T141) begin
      r_irq_timer <= 1'h0;
    end else if(T137) begin
      r_irq_timer <= 1'h1;
    end
    if(T141) begin
      reg_compare <= T139;
    end
    if(reset) begin
      R147 <= 6'h0;
    end else if(T153) begin
      R147 <= T150;
    end
    if(reset) begin
      R154 <= 58'h0;
    end else if(T158) begin
      R154 <= T157;
    end
    if(reset) begin
      R164 <= 6'h0;
    end else if(T170) begin
      R164 <= T167;
    end
    if(reset) begin
      R171 <= 58'h0;
    end else if(T175) begin
      R171 <= T174;
    end
    if(reset) begin
      R181 <= 6'h0;
    end else if(T187) begin
      R181 <= T184;
    end
    if(reset) begin
      R188 <= 58'h0;
    end else if(T192) begin
      R188 <= T191;
    end
    if(reset) begin
      R198 <= 6'h0;
    end else if(T204) begin
      R198 <= T201;
    end
    if(reset) begin
      R205 <= 58'h0;
    end else if(T209) begin
      R205 <= T208;
    end
    if(reset) begin
      R215 <= 6'h0;
    end else if(T221) begin
      R215 <= T218;
    end
    if(reset) begin
      R222 <= 58'h0;
    end else if(T226) begin
      R222 <= T225;
    end
    if(reset) begin
      R232 <= 6'h0;
    end else if(T238) begin
      R232 <= T235;
    end
    if(reset) begin
      R239 <= 58'h0;
    end else if(T243) begin
      R239 <= T242;
    end
    if(reset) begin
      R249 <= 6'h0;
    end else if(T255) begin
      R249 <= T252;
    end
    if(reset) begin
      R256 <= 58'h0;
    end else if(T260) begin
      R256 <= T259;
    end
    if(reset) begin
      R266 <= 6'h0;
    end else if(T272) begin
      R266 <= T269;
    end
    if(reset) begin
      R273 <= 58'h0;
    end else if(T277) begin
      R273 <= T276;
    end
    if(reset) begin
      R283 <= 6'h0;
    end else if(T289) begin
      R283 <= T286;
    end
    if(reset) begin
      R290 <= 58'h0;
    end else if(T294) begin
      R290 <= T293;
    end
    if(reset) begin
      R300 <= 6'h0;
    end else if(T306) begin
      R300 <= T303;
    end
    if(reset) begin
      R307 <= 58'h0;
    end else if(T311) begin
      R307 <= T310;
    end
    if(reset) begin
      R317 <= 6'h0;
    end else if(T323) begin
      R317 <= T320;
    end
    if(reset) begin
      R324 <= 58'h0;
    end else if(T328) begin
      R324 <= T327;
    end
    if(reset) begin
      R334 <= 6'h0;
    end else if(T340) begin
      R334 <= T337;
    end
    if(reset) begin
      R341 <= 58'h0;
    end else if(T345) begin
      R341 <= T344;
    end
    if(reset) begin
      R351 <= 6'h0;
    end else if(T357) begin
      R351 <= T354;
    end
    if(reset) begin
      R358 <= 58'h0;
    end else if(T362) begin
      R358 <= T361;
    end
    if(reset) begin
      R368 <= 6'h0;
    end else if(T374) begin
      R368 <= T371;
    end
    if(reset) begin
      R375 <= 58'h0;
    end else if(T379) begin
      R375 <= T378;
    end
    if(reset) begin
      R385 <= 6'h0;
    end else if(T391) begin
      R385 <= T388;
    end
    if(reset) begin
      R392 <= 58'h0;
    end else if(T396) begin
      R392 <= T395;
    end
    if(reset) begin
      R402 <= 6'h0;
    end else if(T408) begin
      R402 <= T405;
    end
    if(reset) begin
      R409 <= 58'h0;
    end else if(T413) begin
      R409 <= T412;
    end
    if(reset) begin
      reg_tohost <= 64'h0;
    end else if(T427) begin
      reg_tohost <= wdata;
    end else if(T423) begin
      reg_tohost <= 64'h0;
    end
    if(reset) begin
      reg_stats <= 1'h0;
    end else if(T437) begin
      reg_stats <= T436;
    end
    if(io_exception) begin
      reg_cause <= io_cause;
    end
    reg_badvaddr <= T492;
    if(T511) begin
      reg_sup1 <= wdata;
    end
    if(T516) begin
      reg_sup0 <= wdata;
    end
    if(reset) begin
      R521 <= 6'h0;
    end else if(T527) begin
      R521 <= T524;
    end
    if(reset) begin
      R528 <= 58'h0;
    end else if(T532) begin
      R528 <= T531;
    end
    reg_fflags <= T545;
    if(T562) begin
      host_pcr_rep_valid <= 1'h0;
    end else if(host_pcr_req_fire) begin
      host_pcr_rep_valid <= 1'h1;
    end
  end
endmodule

module Datapath(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    input [2:0] io_ctrl_sel_pc,
    input  io_ctrl_killd,
    input  io_ctrl_ren_1,
    input  io_ctrl_ren_0,
    input [2:0] io_ctrl_sel_alu2,
    input [1:0] io_ctrl_sel_alu1,
    input [2:0] io_ctrl_sel_imm,
    input  io_ctrl_fn_dw,
    input [3:0] io_ctrl_fn_alu,
    input  io_ctrl_div_mul_val,
    input  io_ctrl_div_mul_kill,
    //input  io_ctrl_div_val
    //input  io_ctrl_div_kill
    input [2:0] io_ctrl_csr,
    input  io_ctrl_sret,
    input  io_ctrl_mem_load,
    input  io_ctrl_wb_load,
    input  io_ctrl_ex_fp_val,
    input  io_ctrl_mem_fp_val,
    input  io_ctrl_ex_wen,
    input  io_ctrl_ex_valid,
    input  io_ctrl_mem_jalr,
    input  io_ctrl_mem_branch,
    input  io_ctrl_mem_wen,
    input  io_ctrl_wb_wen,
    input [2:0] io_ctrl_ex_mem_type,
    input  io_ctrl_ex_rs2_val,
    input  io_ctrl_ex_rocc_val,
    input  io_ctrl_mem_rocc_val,
    input  io_ctrl_bypass_1,
    input  io_ctrl_bypass_0,
    input [1:0] io_ctrl_bypass_src_1,
    input [1:0] io_ctrl_bypass_src_0,
    input  io_ctrl_ll_ready,
    input  io_ctrl_retire,
    input  io_ctrl_exception,
    input [63:0] io_ctrl_cause,
    input  io_ctrl_badvaddr_wen,
    output[31:0] io_ctrl_inst,
    //output io_ctrl_jalr_eq
    output io_ctrl_mem_br_taken,
    output io_ctrl_mem_misprediction,
    output io_ctrl_div_mul_rdy,
    output io_ctrl_ll_wen,
    output[4:0] io_ctrl_ll_waddr,
    output[4:0] io_ctrl_ex_waddr,
    output io_ctrl_mem_rs1_ra,
    output[4:0] io_ctrl_mem_waddr,
    output[4:0] io_ctrl_wb_waddr,
    output[7:0] io_ctrl_status_ip,
    output[7:0] io_ctrl_status_im,
    output[6:0] io_ctrl_status_zero,
    output io_ctrl_status_er,
    output io_ctrl_status_vm,
    output io_ctrl_status_s64,
    output io_ctrl_status_u64,
    output io_ctrl_status_ef,
    output io_ctrl_status_pei,
    output io_ctrl_status_ei,
    output io_ctrl_status_ps,
    output io_ctrl_status_s,
    output io_ctrl_fp_sboard_clr,
    output[4:0] io_ctrl_fp_sboard_clra,
    output io_ctrl_csr_replay,
    input  io_dmem_req_ready,
    //output io_dmem_req_valid
    //output io_dmem_req_bits_kill
    //output[2:0] io_dmem_req_bits_typ
    //output io_dmem_req_bits_phys
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    //output[4:0] io_dmem_req_bits_cmd
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    //output io_imem_req_valid
    output[43:0] io_imem_req_bits_pc,
    //output io_imem_resp_ready
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    //output io_imem_btb_update_valid
    //output io_imem_btb_update_bits_prediction_valid
    //output io_imem_btb_update_bits_prediction_bits_taken
    //output[42:0] io_imem_btb_update_bits_prediction_bits_target
    //output[2:0] io_imem_btb_update_bits_prediction_bits_entry
    //output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index
    //output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    //output io_imem_btb_update_bits_taken
    //output io_imem_btb_update_bits_isJump
    //output io_imem_btb_update_bits_isCall
    //output io_imem_btb_update_bits_isReturn
    //output io_imem_btb_update_bits_incorrectTarget
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    //output io_imem_invalidate
    output[31:0] io_fpu_inst,
    output[63:0] io_fpu_fromint_data,
    output[2:0] io_fpu_fcsr_rm,
    input  io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output[2:0] io_fpu_dmem_resp_type,
    output[4:0] io_fpu_dmem_resp_tag,
    output[63:0] io_fpu_dmem_resp_data,
    input  io_rocc_cmd_ready,
    //output io_rocc_cmd_valid
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    //output io_rocc_s
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    //output io_rocc_exception
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] wb_reg_inst;
  wire[31:0] T2;
  reg [31:0] mem_reg_inst;
  wire[31:0] T3;
  reg [31:0] ex_reg_inst;
  wire[31:0] T4;
  wire T5;
  wire T6;
  reg  ex_reg_kill;
  wire T7;
  reg  mem_reg_kill;
  wire[31:0] T8;
  wire[63:0] T9;
  reg [63:0] R10;
  reg [63:0] R11;
  wire[63:0] ex_rs_1;
  wire[63:0] T12;
  reg [1:0] ex_reg_rs_lsb_1;
  wire[1:0] T13;
  wire[1:0] T14;
  wire[1:0] T15;
  wire[63:0] id_rs_1;
  wire[63:0] T16;
  wire[63:0] T17;
  reg [63:0] T18 [30:0];
  wire[63:0] T19;
  wire[63:0] wb_wdata;
  wire[63:0] T20;
  wire[63:0] T21;
  wire[63:0] T22;
  reg [63:0] wb_reg_wdata;
  wire[63:0] T23;
  wire[63:0] T24;
  wire[63:0] mem_int_wdata;
  reg [63:0] mem_reg_wdata;
  wire[63:0] T25;
  wire[63:0] alu_io_out;
  wire[63:0] T26;
  wire[44:0] mem_br_target;
  wire[44:0] T27;
  wire[44:0] T28;
  reg [43:0] mem_reg_pc;
  wire[43:0] T29;
  reg [43:0] ex_reg_pc;
  wire[43:0] T30;
  wire[44:0] T31;
  wire[21:0] T32;
  wire[21:0] T33;
  wire[21:0] T34;
  wire[21:0] T35;
  wire[11:0] T36;
  wire[4:0] T37;
  wire[3:0] T38;
  wire[6:0] T39;
  wire[5:0] T40;
  wire T41;
  wire T42;
  wire[9:0] T43;
  wire[8:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[21:0] T52;
  wire[14:0] T53;
  wire[14:0] T54;
  wire[11:0] T55;
  wire[4:0] T56;
  wire[3:0] T57;
  wire[6:0] T58;
  wire[5:0] T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[6:0] T66;
  wire T67;
  wire T68;
  wire[22:0] T69;
  wire T70;
  wire[18:0] T71;
  wire T72;
  wire T73;
  wire[63:0] pcr_io_rw_rdata;
  wire T74;
  wire[63:0] ll_wdata;
  wire[63:0] div_io_resp_bits_data;
  wire T75;
  wire dmem_resp_xpu;
  wire T76;
  wire T77;
  wire dmem_resp_valid;
  wire T78;
  wire T79;
  wire[4:0] T80;
  wire[4:0] T81;
  wire[4:0] wb_waddr;
  wire T82;
  wire T83;
  wire wb_wen;
  wire[4:0] T84;
  wire[4:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  reg [61:0] ex_reg_rs_msb_1;
  wire[61:0] T90;
  wire[61:0] T91;
  wire T92;
  wire T93;
  wire[63:0] T94;
  wire[63:0] T95;
  wire[63:0] T96;
  wire bypass_0;
  wire[63:0] bypass_1;
  wire T97;
  wire[1:0] T98;
  wire[63:0] T99;
  wire[63:0] bypass_2;
  wire[63:0] bypass_3;
  wire T100;
  wire T101;
  reg  ex_reg_rs_bypass_1;
  wire T102;
  wire[4:0] T103;
  wire[4:0] T104;
  wire[63:0] T105;
  reg [63:0] R106;
  reg [63:0] R107;
  wire[63:0] ex_rs_0;
  wire[63:0] T108;
  reg [1:0] ex_reg_rs_lsb_0;
  wire[1:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[63:0] id_rs_0;
  wire[63:0] T112;
  wire[63:0] T113;
  wire[4:0] T114;
  wire[4:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  reg [61:0] ex_reg_rs_msb_0;
  wire[61:0] T120;
  wire[61:0] T121;
  wire T122;
  wire T123;
  wire[63:0] T124;
  wire[63:0] T125;
  wire[63:0] T126;
  wire T127;
  wire[1:0] T128;
  wire[63:0] T129;
  wire T130;
  wire T131;
  reg  ex_reg_rs_bypass_0;
  wire T132;
  wire[4:0] T133;
  wire[4:0] T134;
  wire T135;
  wire[63:0] T136;
  wire[4:0] T137;
  wire[4:0] T138;
  wire[43:0] T139;
  reg [43:0] wb_reg_pc;
  wire[43:0] T140;
  wire T141;
  wire[32:0] T142;
  wire[32:0] T143;
  wire[63:0] pcr_io_time;
  wire T144;
  wire[1135:0] T145;
  wire[63:0] T146;
  wire[63:0] T147;
  wire[63:0] T148;
  wire[63:0] T149;
  wire T150;
  wire[63:0] T151;
  wire T152;
  wire[1:0] T153;
  wire[11:0] T154;
  wire T155;
  wire T156;
  wire dmem_resp_replay;
  reg  ex_reg_ctrl_fn_dw;
  wire T157;
  wire T158;
  reg [3:0] ex_reg_ctrl_fn_alu;
  wire[3:0] T159;
  wire[63:0] ex_op1;
  wire[63:0] T160;
  wire[43:0] T161;
  wire[43:0] T162;
  wire T163;
  reg [1:0] ex_reg_sel_alu1;
  wire[1:0] T164;
  wire[19:0] T165;
  wire T166;
  wire[63:0] T167;
  wire T168;
  wire[63:0] T169;
  wire[63:0] ex_op2;
  wire[63:0] T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[3:0] T173;
  wire T174;
  reg [2:0] ex_reg_sel_alu2;
  wire[2:0] T175;
  wire[27:0] T176;
  wire T177;
  wire[31:0] ex_imm;
  wire[31:0] T178;
  wire[11:0] T179;
  wire[4:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  reg [2:0] ex_reg_sel_imm;
  wire[2:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire[3:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire T196;
  wire[3:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire[6:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire[19:0] T222;
  wire[18:0] T223;
  wire[7:0] T224;
  wire[7:0] T225;
  wire[7:0] T226;
  wire[7:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire[10:0] T231;
  wire[10:0] T232;
  wire[10:0] T233;
  wire[10:0] T234;
  wire T235;
  wire T236;
  wire[31:0] T237;
  wire T238;
  wire[63:0] T239;
  wire T240;
  reg [63:0] wb_reg_rs2;
  wire[63:0] T241;
  reg [63:0] mem_reg_rs2;
  wire[63:0] T242;
  wire[6:0] T243;
  wire[4:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire[4:0] T248;
  wire[4:0] T249;
  wire[6:0] T250;
  wire[4:0] T251;
  wire[6:0] dmem_resp_waddr;
  wire[7:0] T252;
  wire T253;
  wire dmem_resp_fpu;
  wire T254;
  wire[2:0] pcr_io_fcsr_rm;
  wire[42:0] T255;
  wire[42:0] T256;
  wire[42:0] T257;
  wire[43:0] T258;
  wire[44:0] T259;
  wire[44:0] T260;
  wire[44:0] T261;
  wire[43:0] T262;
  wire[43:0] pcr_io_evec;
  wire T263;
  wire[44:0] mem_npc;
  wire[44:0] T264;
  wire[43:0] T265;
  wire[42:0] T266;
  wire T267;
  wire T268;
  wire T269;
  wire[1:0] T270;
  wire T271;
  wire T272;
  wire T273;
  wire[21:0] T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire pcr_io_status_s;
  wire pcr_io_status_ps;
  wire pcr_io_status_ei;
  wire pcr_io_status_pei;
  wire pcr_io_status_ef;
  wire pcr_io_status_u64;
  wire pcr_io_status_s64;
  wire pcr_io_status_vm;
  wire pcr_io_status_er;
  wire[6:0] pcr_io_status_zero;
  wire[7:0] pcr_io_status_im;
  wire[7:0] pcr_io_status_ip;
  wire pcr_io_fatc;
  wire[31:0] pcr_io_ptbr;
  wire[7:0] T281;
  wire[5:0] T282;
  wire[63:0] T283;
  wire[43:0] T284;
  wire[43:0] T285;
  wire[42:0] T286;
  wire[63:0] alu_io_adder_out;
  wire T287;
  wire T288;
  wire T289;
  wire[1:0] T290;
  wire T291;
  wire T292;
  wire T293;
  wire[21:0] T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire pcr_io_replay;
  wire[4:0] T300;
  wire T301;
  wire[4:0] T302;
  wire[4:0] T303;
  wire T304;
  wire[4:0] T305;
  wire[4:0] T306;
  wire[4:0] T307;
  wire[6:0] T308;
  wire[6:0] T309;
  wire[4:0] div_io_resp_bits_tag;
  wire T310;
  wire T311;
  wire div_io_resp_valid;
  wire div_io_req_ready;
  wire T312;
  wire T313;
  wire T314;
  wire[44:0] T315;
  wire T316;
  wire pcr_io_host_debug_stats_pcr;
  wire pcr_io_host_ipi_rep_ready;
  wire pcr_io_host_ipi_req_bits;
  wire pcr_io_host_ipi_req_valid;
  wire[63:0] pcr_io_host_pcr_rep_bits;
  wire pcr_io_host_pcr_rep_valid;
  wire pcr_io_host_pcr_req_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    wb_reg_inst = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_kill = {1{$random}};
    mem_reg_kill = {1{$random}};
    R10 = {2{$random}};
    R11 = {2{$random}};
    ex_reg_rs_lsb_1 = {1{$random}};
    for (initvar = 0; initvar < 31; initvar = initvar+1)
      T18[initvar] = {2{$random}};
    wb_reg_wdata = {2{$random}};
    mem_reg_wdata = {2{$random}};
    mem_reg_pc = {2{$random}};
    ex_reg_pc = {2{$random}};
    ex_reg_rs_msb_1 = {2{$random}};
    ex_reg_rs_bypass_1 = {1{$random}};
    R106 = {2{$random}};
    R107 = {2{$random}};
    ex_reg_rs_lsb_0 = {1{$random}};
    ex_reg_rs_msb_0 = {2{$random}};
    ex_reg_rs_bypass_0 = {1{$random}};
    wb_reg_pc = {2{$random}};
    ex_reg_ctrl_fn_dw = {1{$random}};
    ex_reg_ctrl_fn_alu = {1{$random}};
    ex_reg_sel_alu1 = {1{$random}};
    ex_reg_sel_alu2 = {1{$random}};
    ex_reg_sel_imm = {1{$random}};
    wb_reg_rs2 = {2{$random}};
    mem_reg_rs2 = {2{$random}};
  end
`endif

  assign T0 = reset ^ 1'h1;
  assign T1 = wb_reg_inst;
  assign T2 = T7 ? mem_reg_inst : wb_reg_inst;
  assign T3 = T6 ? ex_reg_inst : mem_reg_inst;
  assign T4 = T5 ? io_imem_resp_bits_data : ex_reg_inst;
  assign T5 = io_ctrl_killd ^ 1'h1;
  assign T6 = ex_reg_kill ^ 1'h1;
  assign T7 = mem_reg_kill ^ 1'h1;
  assign T8 = wb_reg_inst;
  assign T9 = R10;
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? T94 : T12;
  assign T12 = {ex_reg_rs_msb_1, ex_reg_rs_lsb_1};
  assign T13 = T89 ? io_ctrl_bypass_src_1 : T14;
  assign T14 = T88 ? T15 : ex_reg_rs_lsb_1;
  assign T15 = id_rs_1[1'h1:1'h0];
  assign id_rs_1 = T16;
  assign T16 = T86 ? wb_wdata : T17;
  assign T17 = T18[T84];
  assign wb_wdata = T20;
  assign T20 = T75 ? io_dmem_resp_bits_data_subword : T21;
  assign T21 = io_ctrl_ll_wen ? ll_wdata : T22;
  assign T22 = T74 ? pcr_io_rw_rdata : wb_reg_wdata;
  assign T23 = T7 ? T24 : wb_reg_wdata;
  assign T24 = T73 ? io_fpu_toint_data : mem_int_wdata;
  assign mem_int_wdata = io_ctrl_mem_jalr ? T26 : mem_reg_wdata;
  assign T25 = T6 ? alu_io_out : mem_reg_wdata;
  assign T26 = {T71, mem_br_target};
  assign mem_br_target = T31 + T27;
  assign T27 = T28;
  assign T28 = {1'h0, mem_reg_pc};
  assign T29 = T6 ? ex_reg_pc : mem_reg_pc;
  assign T30 = T5 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T31 = {T69, T32};
  assign T32 = T68 ? T52 : T33;
  assign T33 = T49 ? T34 : 22'h4;
  assign T34 = T35;
  assign T35 = {T43, T36};
  assign T36 = {T39, T37};
  assign T37 = {T38, 1'h0};
  assign T38 = mem_reg_inst[5'h18:5'h15];
  assign T39 = {T41, T40};
  assign T40 = mem_reg_inst[5'h1e:5'h19];
  assign T41 = T42;
  assign T42 = mem_reg_inst[5'h14:5'h14];
  assign T43 = {T47, T44};
  assign T44 = {T47, T45};
  assign T45 = T46;
  assign T46 = mem_reg_inst[5'h13:4'hc];
  assign T47 = T48;
  assign T48 = mem_reg_inst[5'h1f:5'h1f];
  assign T49 = T51 & T50;
  assign T50 = io_ctrl_mem_branch ^ 1'h1;
  assign T51 = io_ctrl_mem_jalr ^ 1'h1;
  assign T52 = {T66, T53};
  assign T53 = T54;
  assign T54 = {T62, T55};
  assign T55 = {T58, T56};
  assign T56 = {T57, 1'h0};
  assign T57 = mem_reg_inst[4'hb:4'h8];
  assign T58 = {T60, T59};
  assign T59 = mem_reg_inst[5'h1e:5'h19];
  assign T60 = T61;
  assign T61 = mem_reg_inst[3'h7:3'h7];
  assign T62 = {T64, T63};
  assign T63 = {T64, T64};
  assign T64 = T65;
  assign T65 = mem_reg_inst[5'h1f:5'h1f];
  assign T66 = T67 ? 7'h7f : 7'h0;
  assign T67 = T53[4'he:4'he];
  assign T68 = io_ctrl_mem_branch & io_ctrl_mem_br_taken;
  assign T69 = T70 ? 23'h7fffff : 23'h0;
  assign T70 = T32[5'h15:5'h15];
  assign T71 = T72 ? 19'h7ffff : 19'h0;
  assign T72 = mem_br_target[6'h2c:6'h2c];
  assign T73 = io_ctrl_mem_fp_val & io_ctrl_mem_wen;
  assign T74 = io_ctrl_csr != 3'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign T75 = dmem_resp_valid & dmem_resp_xpu;
  assign dmem_resp_xpu = T76 ^ 1'h1;
  assign T76 = T77;
  assign T77 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign T78 = T82 & T79;
  assign T79 = T80 < 5'h1f;
  assign T80 = T81[3'h4:1'h0];
  assign T81 = ~ wb_waddr;
  assign wb_waddr = io_ctrl_ll_wen ? io_ctrl_ll_waddr : io_ctrl_wb_waddr;
  assign T82 = wb_wen & T83;
  assign T83 = wb_waddr != 5'h0;
  assign wb_wen = io_ctrl_ll_wen | io_ctrl_wb_wen;
  assign T84 = ~ T85;
  assign T85 = io_imem_resp_bits_data[5'h18:5'h14];
  assign T86 = T82 & T87;
  assign T87 = wb_waddr == T85;
  assign T88 = T5 & io_ctrl_ren_1;
  assign T89 = T5 & io_ctrl_bypass_1;
  assign T90 = T92 ? T91 : ex_reg_rs_msb_1;
  assign T91 = id_rs_1 >> 2'h2;
  assign T92 = T88 & T93;
  assign T93 = io_ctrl_bypass_1 ^ 1'h1;
  assign T94 = T101 ? T99 : T95;
  assign T95 = T97 ? bypass_1 : T96;
  assign T96 = {63'h0, bypass_0};
  assign bypass_0 = 1'h0;
  assign bypass_1 = mem_reg_wdata;
  assign T97 = T98[1'h0:1'h0];
  assign T98 = ex_reg_rs_lsb_1;
  assign T99 = T100 ? bypass_3 : bypass_2;
  assign bypass_2 = wb_reg_wdata;
  assign bypass_3 = io_dmem_resp_bits_data;
  assign T100 = T98[1'h0:1'h0];
  assign T101 = T98[1'h1:1'h1];
  assign T102 = T5 ? io_ctrl_bypass_1 : ex_reg_rs_bypass_1;
  assign T103 = T104;
  assign T104 = wb_reg_inst[5'h18:5'h14];
  assign T105 = R106;
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? T124 : T108;
  assign T108 = {ex_reg_rs_msb_0, ex_reg_rs_lsb_0};
  assign T109 = T119 ? io_ctrl_bypass_src_0 : T110;
  assign T110 = T118 ? T111 : ex_reg_rs_lsb_0;
  assign T111 = id_rs_0[1'h1:1'h0];
  assign id_rs_0 = T112;
  assign T112 = T116 ? wb_wdata : T113;
  assign T113 = T18[T114];
  assign T114 = ~ T115;
  assign T115 = io_imem_resp_bits_data[5'h13:4'hf];
  assign T116 = T82 & T117;
  assign T117 = wb_waddr == T115;
  assign T118 = T5 & io_ctrl_ren_0;
  assign T119 = T5 & io_ctrl_bypass_0;
  assign T120 = T122 ? T121 : ex_reg_rs_msb_0;
  assign T121 = id_rs_0 >> 2'h2;
  assign T122 = T118 & T123;
  assign T123 = io_ctrl_bypass_0 ^ 1'h1;
  assign T124 = T131 ? T129 : T125;
  assign T125 = T127 ? bypass_1 : T126;
  assign T126 = {63'h0, bypass_0};
  assign T127 = T128[1'h0:1'h0];
  assign T128 = ex_reg_rs_lsb_0;
  assign T129 = T130 ? bypass_3 : bypass_2;
  assign T130 = T128[1'h0:1'h0];
  assign T131 = T128[1'h1:1'h1];
  assign T132 = T5 ? io_ctrl_bypass_0 : ex_reg_rs_bypass_0;
  assign T133 = T134;
  assign T134 = wb_reg_inst[5'h13:4'hf];
  assign T135 = wb_wen;
  assign T136 = wb_wdata;
  assign T137 = T138;
  assign T138 = wb_wen ? wb_waddr : 5'h0;
  assign T139 = wb_reg_pc;
  assign T140 = T7 ? mem_reg_pc : wb_reg_pc;
  assign T141 = io_ctrl_retire;
  assign T142 = T143;
  assign T143 = pcr_io_time[6'h20:1'h0];
  assign T144 = io_host_id;
  assign T146 = T152 ? T151 : T147;
  assign T147 = T150 ? T148 : wb_reg_wdata;
  assign T148 = pcr_io_rw_rdata & T149;
  assign T149 = ~ wb_reg_wdata;
  assign T150 = io_ctrl_csr == 3'h3;
  assign T151 = pcr_io_rw_rdata | wb_reg_wdata;
  assign T152 = io_ctrl_csr == 3'h2;
  assign T153 = io_ctrl_csr[1'h1:1'h0];
  assign T154 = wb_reg_inst[5'h1f:5'h14];
  assign T155 = T156 ? 1'h0 : io_ctrl_ll_ready;
  assign T156 = dmem_resp_replay & dmem_resp_xpu;
  assign dmem_resp_replay = io_dmem_resp_bits_replay & io_dmem_resp_bits_has_data;
  assign T157 = T5 ? T158 : ex_reg_ctrl_fn_dw;
  assign T158 = io_ctrl_fn_dw;
  assign T159 = T5 ? io_ctrl_fn_alu : ex_reg_ctrl_fn_alu;
  assign ex_op1 = T168 ? T167 : T160;
  assign T160 = {T165, T161};
  assign T161 = T163 ? T162 : 44'h0;
  assign T162 = ex_reg_pc;
  assign T163 = ex_reg_sel_alu1 == 2'h2;
  assign T164 = T5 ? io_ctrl_sel_alu1 : ex_reg_sel_alu1;
  assign T165 = T166 ? 20'hfffff : 20'h0;
  assign T166 = T161[6'h2b:6'h2b];
  assign T167 = ex_rs_0;
  assign T168 = ex_reg_sel_alu1 == 2'h1;
  assign T169 = ex_op2;
  assign ex_op2 = T240 ? T239 : T170;
  assign T170 = {T237, T171};
  assign T171 = T236 ? ex_imm : T172;
  assign T172 = {T176, T173};
  assign T173 = T174 ? 4'h4 : 4'h0;
  assign T174 = ex_reg_sel_alu2 == 3'h1;
  assign T175 = T5 ? io_ctrl_sel_alu2 : ex_reg_sel_alu2;
  assign T176 = T177 ? 28'hfffffff : 28'h0;
  assign T177 = T173[2'h3:2'h3];
  assign ex_imm = T178;
  assign T178 = {T222, T179};
  assign T179 = {T202, T180};
  assign T180 = {T191, T181};
  assign T181 = T190 ? T189 : T182;
  assign T182 = T188 ? T187 : T183;
  assign T183 = T185 ? T184 : 1'h0;
  assign T184 = ex_reg_inst[4'hf:4'hf];
  assign T185 = ex_reg_sel_imm == 3'h5;
  assign T186 = T5 ? io_ctrl_sel_imm : ex_reg_sel_imm;
  assign T187 = ex_reg_inst[5'h14:5'h14];
  assign T188 = ex_reg_sel_imm == 3'h4;
  assign T189 = ex_reg_inst[3'h7:3'h7];
  assign T190 = ex_reg_sel_imm == 3'h0;
  assign T191 = T201 ? 4'h0 : T192;
  assign T192 = T198 ? T197 : T193;
  assign T193 = T196 ? T195 : T194;
  assign T194 = ex_reg_inst[5'h18:5'h15];
  assign T195 = ex_reg_inst[5'h13:5'h10];
  assign T196 = ex_reg_sel_imm == 3'h5;
  assign T197 = ex_reg_inst[4'hb:4'h8];
  assign T198 = T200 | T199;
  assign T199 = ex_reg_sel_imm == 3'h1;
  assign T200 = ex_reg_sel_imm == 3'h0;
  assign T201 = ex_reg_sel_imm == 3'h2;
  assign T202 = {T208, T203};
  assign T203 = T205 ? 6'h0 : T204;
  assign T204 = ex_reg_inst[5'h1e:5'h19];
  assign T205 = T207 | T206;
  assign T206 = ex_reg_sel_imm == 3'h5;
  assign T207 = ex_reg_sel_imm == 3'h2;
  assign T208 = T219 ? 1'h0 : T209;
  assign T209 = T218 ? T216 : T210;
  assign T210 = T215 ? T213 : T211;
  assign T211 = T212;
  assign T212 = ex_reg_inst[5'h1f:5'h1f];
  assign T213 = T214;
  assign T214 = ex_reg_inst[3'h7:3'h7];
  assign T215 = ex_reg_sel_imm == 3'h1;
  assign T216 = T217;
  assign T217 = ex_reg_inst[5'h14:5'h14];
  assign T218 = ex_reg_sel_imm == 3'h3;
  assign T219 = T221 | T220;
  assign T220 = ex_reg_sel_imm == 3'h5;
  assign T221 = ex_reg_sel_imm == 3'h2;
  assign T222 = {T211, T223};
  assign T223 = {T231, T224};
  assign T224 = T228 ? T227 : T225;
  assign T225 = T226;
  assign T226 = ex_reg_inst[5'h13:4'hc];
  assign T227 = T211 ? 8'hff : 8'h0;
  assign T228 = T230 & T229;
  assign T229 = ex_reg_sel_imm != 3'h3;
  assign T230 = ex_reg_sel_imm != 3'h2;
  assign T231 = T235 ? T233 : T232;
  assign T232 = T211 ? 11'h7ff : 11'h0;
  assign T233 = T234;
  assign T234 = ex_reg_inst[5'h1e:5'h14];
  assign T235 = ex_reg_sel_imm == 3'h2;
  assign T236 = ex_reg_sel_alu2 == 3'h3;
  assign T237 = T238 ? 32'hffffffff : 32'h0;
  assign T238 = T171[5'h1f:5'h1f];
  assign T239 = ex_rs_1;
  assign T240 = ex_reg_sel_alu2 == 3'h2;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign T241 = io_ctrl_mem_rocc_val ? mem_reg_rs2 : wb_reg_rs2;
  assign T242 = io_ctrl_ex_rs2_val ? ex_rs_1 : mem_reg_rs2;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_inst_opcode = T243;
  assign T243 = wb_reg_inst[3'h6:1'h0];
  assign io_rocc_cmd_bits_inst_rd = T244;
  assign T244 = wb_reg_inst[4'hb:3'h7];
  assign io_rocc_cmd_bits_inst_xs2 = T245;
  assign T245 = wb_reg_inst[4'hc:4'hc];
  assign io_rocc_cmd_bits_inst_xs1 = T246;
  assign T246 = wb_reg_inst[4'hd:4'hd];
  assign io_rocc_cmd_bits_inst_xd = T247;
  assign T247 = wb_reg_inst[4'he:4'he];
  assign io_rocc_cmd_bits_inst_rs1 = T248;
  assign T248 = wb_reg_inst[5'h13:4'hf];
  assign io_rocc_cmd_bits_inst_rs2 = T249;
  assign T249 = wb_reg_inst[5'h18:5'h14];
  assign io_rocc_cmd_bits_inst_funct = T250;
  assign T250 = wb_reg_inst[5'h1f:5'h19];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data;
  assign io_fpu_dmem_resp_tag = T251;
  assign T251 = dmem_resp_waddr[3'h4:1'h0];
  assign dmem_resp_waddr = T252 >> 1'h1;
  assign T252 = io_dmem_resp_bits_tag;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_val = T253;
  assign T253 = dmem_resp_valid & dmem_resp_fpu;
  assign dmem_resp_fpu = T254;
  assign T254 = io_dmem_resp_bits_tag[1'h0:1'h0];
  assign io_fpu_fcsr_rm = pcr_io_fcsr_rm;
  assign io_fpu_fromint_data = ex_rs_0;
  assign io_fpu_inst = io_imem_resp_bits_data;
  assign io_imem_btb_update_bits_returnAddr = T255;
  assign T255 = mem_int_wdata[6'h2a:1'h0];
  assign io_imem_btb_update_bits_target = T256;
  assign T256 = io_imem_req_bits_pc[6'h2a:1'h0];
  assign io_imem_btb_update_bits_pc = T257;
  assign T257 = mem_reg_pc[6'h2a:1'h0];
  assign io_imem_req_bits_pc = T258;
  assign T258 = T259[6'h2b:1'h0];
  assign T259 = T260;
  assign T260 = T280 ? mem_npc : T261;
  assign T261 = {1'h0, T262};
  assign T262 = T263 ? pcr_io_evec : wb_reg_pc;
  assign T263 = io_ctrl_sel_pc == 3'h3;
  assign mem_npc = io_ctrl_mem_jalr ? T264 : mem_br_target;
  assign T264 = {1'h0, T265};
  assign T265 = {T267, T266};
  assign T266 = mem_reg_wdata[6'h2a:1'h0];
  assign T267 = T277 ? T276 : T268;
  assign T268 = T272 ? T271 : T269;
  assign T269 = T270[1'h0:1'h0];
  assign T270 = mem_reg_wdata[6'h2b:6'h2a];
  assign T271 = T270 == 2'h3;
  assign T272 = T275 | T273;
  assign T273 = T274 == 22'h3ffffe;
  assign T274 = mem_reg_wdata >> 6'h2a;
  assign T275 = T274 == 22'h3fffff;
  assign T276 = T270 != 2'h0;
  assign T277 = T279 | T278;
  assign T278 = T274 == 22'h1;
  assign T279 = T274 == 22'h0;
  assign T280 = io_ctrl_sel_pc == 3'h1;
  assign io_ptw_status_s = pcr_io_status_s;
  assign io_ptw_status_ps = pcr_io_status_ps;
  assign io_ptw_status_ei = pcr_io_status_ei;
  assign io_ptw_status_pei = pcr_io_status_pei;
  assign io_ptw_status_ef = pcr_io_status_ef;
  assign io_ptw_status_u64 = pcr_io_status_u64;
  assign io_ptw_status_s64 = pcr_io_status_s64;
  assign io_ptw_status_vm = pcr_io_status_vm;
  assign io_ptw_status_er = pcr_io_status_er;
  assign io_ptw_status_zero = pcr_io_status_zero;
  assign io_ptw_status_im = pcr_io_status_im;
  assign io_ptw_status_ip = pcr_io_status_ip;
  assign io_ptw_sret = io_ctrl_sret;
  assign io_ptw_invalidate = pcr_io_fatc;
  assign io_ptw_ptbr = pcr_io_ptbr;
  assign io_dmem_req_bits_tag = T281;
  assign T281 = {2'h0, T282};
  assign T282 = {io_ctrl_ex_waddr, io_ctrl_ex_fp_val};
  assign io_dmem_req_bits_data = T283;
  assign T283 = io_ctrl_mem_fp_val ? io_fpu_store_data : mem_reg_rs2;
  assign io_dmem_req_bits_addr = T284;
  assign T284 = T285;
  assign T285 = {T287, T286};
  assign T286 = alu_io_adder_out[6'h2a:1'h0];
  assign T287 = T297 ? T296 : T288;
  assign T288 = T292 ? T291 : T289;
  assign T289 = T290[1'h0:1'h0];
  assign T290 = alu_io_adder_out[6'h2b:6'h2a];
  assign T291 = T290 == 2'h3;
  assign T292 = T295 | T293;
  assign T293 = T294 == 22'h3ffffe;
  assign T294 = ex_rs_0 >> 6'h2a;
  assign T295 = T294 == 22'h3fffff;
  assign T296 = T290 != 2'h0;
  assign T297 = T299 | T298;
  assign T298 = T294 == 22'h1;
  assign T299 = T294 == 22'h0;
  assign io_ctrl_csr_replay = pcr_io_replay;
  assign io_ctrl_fp_sboard_clra = T300;
  assign T300 = dmem_resp_waddr[3'h4:1'h0];
  assign io_ctrl_fp_sboard_clr = T301;
  assign T301 = dmem_resp_replay & dmem_resp_fpu;
  assign io_ctrl_status_s = pcr_io_status_s;
  assign io_ctrl_status_ps = pcr_io_status_ps;
  assign io_ctrl_status_ei = pcr_io_status_ei;
  assign io_ctrl_status_pei = pcr_io_status_pei;
  assign io_ctrl_status_ef = pcr_io_status_ef;
  assign io_ctrl_status_u64 = pcr_io_status_u64;
  assign io_ctrl_status_s64 = pcr_io_status_s64;
  assign io_ctrl_status_vm = pcr_io_status_vm;
  assign io_ctrl_status_er = pcr_io_status_er;
  assign io_ctrl_status_zero = pcr_io_status_zero;
  assign io_ctrl_status_im = pcr_io_status_im;
  assign io_ctrl_status_ip = pcr_io_status_ip;
  assign io_ctrl_wb_waddr = T302;
  assign T302 = wb_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_waddr = T303;
  assign T303 = mem_reg_inst[4'hb:3'h7];
  assign io_ctrl_mem_rs1_ra = T304;
  assign T304 = T305 == 5'h1;
  assign T305 = mem_reg_inst[5'h13:4'hf];
  assign io_ctrl_ex_waddr = T306;
  assign T306 = ex_reg_inst[4'hb:3'h7];
  assign io_ctrl_ll_waddr = T307;
  assign T307 = T308[3'h4:1'h0];
  assign T308 = T156 ? dmem_resp_waddr : T309;
  assign T309 = {2'h0, div_io_resp_bits_tag};
  assign io_ctrl_ll_wen = T310;
  assign T310 = T156 ? 1'h1 : T311;
  assign T311 = T155 & div_io_resp_valid;
  assign io_ctrl_div_mul_rdy = div_io_req_ready;
  assign io_ctrl_mem_misprediction = T312;
  assign T312 = T314 | T313;
  assign T313 = io_ctrl_ex_valid ^ 1'h1;
  assign T314 = mem_npc != T315;
  assign T315 = {1'h0, ex_reg_pc};
  assign io_ctrl_mem_br_taken = T316;
  assign T316 = mem_reg_wdata[1'h0:1'h0];
  assign io_ctrl_inst = io_imem_resp_bits_data;
  assign io_host_debug_stats_pcr = pcr_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = pcr_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = pcr_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = pcr_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = pcr_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = pcr_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = pcr_io_host_pcr_req_ready;
  ALU alu(
       .io_dw( ex_reg_ctrl_fn_dw ),
       .io_fn( ex_reg_ctrl_fn_alu ),
       .io_in2( T169 ),
       .io_in1( ex_op1 ),
       .io_out( alu_io_out ),
       .io_adder_out( alu_io_adder_out )
  );
  MulDiv div(.clk(clk), .reset(reset),
       .io_req_ready( div_io_req_ready ),
       .io_req_valid( io_ctrl_div_mul_val ),
       .io_req_bits_fn( ex_reg_ctrl_fn_alu ),
       .io_req_bits_dw( ex_reg_ctrl_fn_dw ),
       .io_req_bits_in1( ex_rs_0 ),
       .io_req_bits_in2( ex_rs_1 ),
       .io_req_bits_tag( io_ctrl_ex_waddr ),
       .io_kill( io_ctrl_div_mul_kill ),
       .io_resp_ready( T155 ),
       .io_resp_valid( div_io_resp_valid ),
       .io_resp_bits_data( div_io_resp_bits_data ),
       .io_resp_bits_tag( div_io_resp_bits_tag )
  );
  CSRFile pcr(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( pcr_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( pcr_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( pcr_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( pcr_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( pcr_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( pcr_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( pcr_io_host_debug_stats_pcr ),
       .io_rw_addr( T154 ),
       .io_rw_cmd( T153 ),
       .io_rw_rdata( pcr_io_rw_rdata ),
       .io_rw_wdata( T146 ),
       .io_status_ip( pcr_io_status_ip ),
       .io_status_im( pcr_io_status_im ),
       .io_status_zero( pcr_io_status_zero ),
       .io_status_er( pcr_io_status_er ),
       .io_status_vm( pcr_io_status_vm ),
       .io_status_s64( pcr_io_status_s64 ),
       .io_status_u64( pcr_io_status_u64 ),
       .io_status_ef( pcr_io_status_ef ),
       .io_status_pei( pcr_io_status_pei ),
       .io_status_ei( pcr_io_status_ei ),
       .io_status_ps( pcr_io_status_ps ),
       .io_status_s( pcr_io_status_s ),
       .io_ptbr( pcr_io_ptbr ),
       .io_evec( pcr_io_evec ),
       .io_exception( io_ctrl_exception ),
       .io_retire( io_ctrl_retire ),
       .io_uarch_counters_15( 1'h0 ),
       .io_uarch_counters_14( 1'h0 ),
       .io_uarch_counters_13( 1'h0 ),
       .io_uarch_counters_12( 1'h0 ),
       .io_uarch_counters_11( 1'h0 ),
       .io_uarch_counters_10( 1'h0 ),
       .io_uarch_counters_9( 1'h0 ),
       .io_uarch_counters_8( 1'h0 ),
       .io_uarch_counters_7( 1'h0 ),
       .io_uarch_counters_6( 1'h0 ),
       .io_uarch_counters_5( 1'h0 ),
       .io_uarch_counters_4( 1'h0 ),
       .io_uarch_counters_3( 1'h0 ),
       .io_uarch_counters_2( 1'h0 ),
       .io_uarch_counters_1( 1'h0 ),
       .io_uarch_counters_0( 1'h0 ),
       .io_cause( io_ctrl_cause ),
       .io_badvaddr_wen( io_ctrl_badvaddr_wen ),
       .io_pc( wb_reg_pc ),
       .io_sret( io_ctrl_sret ),
       .io_fatc( pcr_io_fatc ),
       .io_replay( pcr_io_replay ),
       .io_time( pcr_io_time ),
       .io_fcsr_rm( pcr_io_fcsr_rm ),
       .io_fcsr_flags_valid( io_fpu_fcsr_flags_valid ),
       .io_fcsr_flags_bits( io_fpu_fcsr_flags_bits ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );

  always @(posedge clk) begin
    if(T7) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if(T6) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(T5) begin
      ex_reg_inst <= io_imem_resp_bits_data;
    end
    ex_reg_kill <= io_ctrl_killd;
    mem_reg_kill <= ex_reg_kill;
    R10 <= R11;
    if(ex_reg_rs_bypass_1) begin
      R11 <= T94;
    end else begin
      R11 <= T12;
    end
    if(T89) begin
      ex_reg_rs_lsb_1 <= io_ctrl_bypass_src_1;
    end else if(T88) begin
      ex_reg_rs_lsb_1 <= T15;
    end
    if (T78)
      T18[T81] <= wb_wdata;
    if(T7) begin
      wb_reg_wdata <= T24;
    end
    if(T6) begin
      mem_reg_wdata <= alu_io_out;
    end
    if(T6) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if(T5) begin
      ex_reg_pc <= io_imem_resp_bits_pc;
    end
    if(T92) begin
      ex_reg_rs_msb_1 <= T91;
    end
    if(T5) begin
      ex_reg_rs_bypass_1 <= io_ctrl_bypass_1;
    end
    R106 <= R107;
    if(ex_reg_rs_bypass_0) begin
      R107 <= T124;
    end else begin
      R107 <= T108;
    end
    if(T119) begin
      ex_reg_rs_lsb_0 <= io_ctrl_bypass_src_0;
    end else if(T118) begin
      ex_reg_rs_lsb_0 <= T111;
    end
    if(T122) begin
      ex_reg_rs_msb_0 <= T121;
    end
    if(T5) begin
      ex_reg_rs_bypass_0 <= io_ctrl_bypass_0;
    end
    if(T7) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if(T5) begin
      ex_reg_ctrl_fn_dw <= T158;
    end
    if(T5) begin
      ex_reg_ctrl_fn_alu <= io_ctrl_fn_alu;
    end
    if(T5) begin
      ex_reg_sel_alu1 <= io_ctrl_sel_alu1;
    end
    if(T5) begin
      ex_reg_sel_alu2 <= io_ctrl_sel_alu2;
    end
    if(T5) begin
      ex_reg_sel_imm <= io_ctrl_sel_imm;
    end
    if(io_ctrl_mem_rocc_val) begin
      wb_reg_rs2 <= mem_reg_rs2;
    end
    if(io_ctrl_ex_rs2_val) begin
      mem_reg_rs2 <= ex_rs_1;
    end
`ifndef SYNTHESIS
`ifdef PRINTF_COND
    if (`PRINTF_COND)
`endif
      if (T0)
        $fwrite(32'h80000002, "C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n", T144, T142, T141, T139, T137, T136, T135, T133, T105, T103, T9, T8, T1);
`endif
  end
endmodule

module FPUDecoder(
    input [31:0] io_inst,
    output[4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_round
);

  wire T0;
  wire T1;
  wire[31:0] T2;
  wire T3;
  wire T4;
  wire[31:0] T5;
  wire T6;
  wire T7;
  wire[31:0] T8;
  wire T9;
  wire T10;
  wire[31:0] T11;
  wire T12;
  wire T13;
  wire[31:0] T14;
  wire T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire T19;
  wire[31:0] T20;
  wire T21;
  wire[31:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire T29;
  wire[31:0] T30;
  wire T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire[31:0] T35;
  wire T36;
  wire T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire T41;
  wire[31:0] T42;
  wire T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire T53;
  wire T54;
  wire[31:0] T55;
  wire T56;
  wire T57;
  wire[31:0] T58;
  wire T59;
  wire T60;
  wire[31:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[31:0] T65;
  wire T66;
  wire T67;
  wire[31:0] T68;
  wire T69;
  wire T70;
  wire[31:0] T71;
  wire T72;
  wire T73;
  wire[31:0] T74;
  wire T75;
  wire T76;
  wire[31:0] T77;
  wire T78;
  wire T79;
  wire[31:0] T80;
  wire T81;
  wire[31:0] T82;
  wire T83;
  wire T84;
  wire[31:0] T85;
  wire T86;
  wire T87;
  wire[31:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire[31:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire[31:0] T114;
  wire[4:0] T115;
  wire[3:0] T116;
  wire[2:0] T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[31:0] T121;
  wire T122;
  wire[31:0] T123;
  wire T124;
  wire T125;
  wire[31:0] T126;
  wire T127;
  wire[31:0] T128;
  wire T129;
  wire T130;
  wire[31:0] T131;
  wire T132;
  wire[31:0] T133;
  wire T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire[31:0] T138;


  assign io_sigs_round = T0;
  assign T0 = T3 | T1;
  assign T1 = T2 == 32'he0000053;
  assign T2 = io_inst & 32'hedf0707f;
  assign T3 = T6 | T4;
  assign T4 = T5 == 32'he0000053;
  assign T5 = io_inst & 32'hfdf0607f;
  assign T6 = T9 | T7;
  assign T7 = T8 == 32'hc0000053;
  assign T8 = io_inst & 32'hedc0007f;
  assign T9 = T12 | T10;
  assign T10 = T11 == 32'h42000053;
  assign T11 = io_inst & 32'h7ff0007f;
  assign T12 = T15 | T13;
  assign T13 = T14 == 32'h40100053;
  assign T14 = io_inst & 32'h7ff0007f;
  assign T15 = T18 | T16;
  assign T16 = T17 == 32'h53;
  assign T17 = io_inst & 32'hec00007f;
  assign T18 = T21 | T19;
  assign T19 = T20 == 32'h53;
  assign T20 = io_inst & 32'hf400007f;
  assign T21 = T22 == 32'h43;
  assign T22 = io_inst & 32'h4000073;
  assign io_sigs_fma = T23;
  assign T23 = T24 | T16;
  assign T24 = T21 | T19;
  assign io_sigs_fastpipe = T25;
  assign T25 = T28 | T26;
  assign T26 = T27 == 32'h42000053;
  assign T27 = io_inst & 32'hfff0007f;
  assign T28 = T31 | T29;
  assign T29 = T30 == 32'h40100053;
  assign T30 = io_inst & 32'hfff0007f;
  assign T31 = T34 | T32;
  assign T32 = T33 == 32'h20000053;
  assign T33 = io_inst & 32'hf400607f;
  assign T34 = T35 == 32'h20000053;
  assign T35 = io_inst & 32'hfc00507f;
  assign io_sigs_toint = T36;
  assign T36 = T37 | T4;
  assign T37 = T40 | T38;
  assign T38 = T39 == 32'hc0000053;
  assign T39 = io_inst & 32'hfdc0007f;
  assign T40 = T43 | T41;
  assign T41 = T42 == 32'ha0000053;
  assign T42 = io_inst & 32'hfc00507f;
  assign T43 = T46 | T44;
  assign T44 = T45 == 32'ha0000053;
  assign T45 = io_inst & 32'hfc00607f;
  assign T46 = T47 == 32'h2027;
  assign T47 = io_inst & 32'h607f;
  assign io_sigs_fromint = T48;
  assign T48 = T51 | T49;
  assign T49 = T50 == 32'hf0000053;
  assign T50 = io_inst & 32'hfdf0707f;
  assign T51 = T52 == 32'hd0000053;
  assign T52 = io_inst & 32'hfdc0007f;
  assign io_sigs_single = T53;
  assign T53 = T56 | T54;
  assign T54 = T55 == 32'he0000053;
  assign T55 = io_inst & 32'heff0707f;
  assign T56 = T59 | T57;
  assign T57 = T58 == 32'he0000053;
  assign T58 = io_inst & 32'hfff0607f;
  assign T59 = T62 | T60;
  assign T60 = T61 == 32'hc0000053;
  assign T61 = io_inst & 32'hefc0007f;
  assign T62 = T63 | T13;
  assign T63 = T66 | T64;
  assign T64 = T65 == 32'h20000053;
  assign T65 = io_inst & 32'h7e00507f;
  assign T66 = T69 | T67;
  assign T67 = T68 == 32'h20000053;
  assign T68 = io_inst & 32'h7e00607f;
  assign T69 = T72 | T70;
  assign T70 = T71 == 32'h20000053;
  assign T71 = io_inst & 32'hf600607f;
  assign T72 = T75 | T73;
  assign T73 = T74 == 32'h2007;
  assign T74 = io_inst & 32'h705f;
  assign T75 = T78 | T76;
  assign T76 = T77 == 32'h53;
  assign T77 = io_inst & 32'hee00007f;
  assign T78 = T81 | T79;
  assign T79 = T80 == 32'h53;
  assign T80 = io_inst & 32'hf600007f;
  assign T81 = T82 == 32'h43;
  assign T82 = io_inst & 32'h6000073;
  assign io_sigs_swap23 = T19;
  assign io_sigs_ren3 = T21;
  assign io_sigs_ren2 = T83;
  assign T83 = T86 | T84;
  assign T84 = T85 == 32'h20000053;
  assign T85 = io_inst & 32'h7c00507f;
  assign T86 = T89 | T87;
  assign T87 = T88 == 32'h20000053;
  assign T88 = io_inst & 32'h7c00607f;
  assign T89 = T90 | T32;
  assign T90 = T91 | T46;
  assign T91 = T92 | T16;
  assign T92 = T21 | T19;
  assign io_sigs_ren1 = T93;
  assign T93 = T94 | T4;
  assign T94 = T95 | T38;
  assign T95 = T96 | T10;
  assign T96 = T97 | T13;
  assign T97 = T98 | T84;
  assign T98 = T99 | T87;
  assign T99 = T100 | T32;
  assign T100 = T101 | T16;
  assign T101 = T21 | T19;
  assign io_sigs_wen = T102;
  assign T102 = T103 | T49;
  assign T103 = T104 | T51;
  assign T104 = T105 | T26;
  assign T105 = T106 | T29;
  assign T106 = T107 | T32;
  assign T107 = T108 | T34;
  assign T108 = T111 | T109;
  assign T109 = T110 == 32'h2007;
  assign T110 = io_inst & 32'h607f;
  assign T111 = T112 | T16;
  assign T112 = T21 | T19;
  assign io_sigs_ldst = T113;
  assign T113 = T114 == 32'h2007;
  assign T114 = io_inst & 32'h605f;
  assign io_sigs_cmd = T115;
  assign T115 = {T137, T116};
  assign T116 = {T134, T117};
  assign T117 = {T129, T118};
  assign T118 = {T124, T119};
  assign T119 = T122 | T120;
  assign T120 = T121 == 32'h8000010;
  assign T121 = io_inst & 32'h8000010;
  assign T122 = T123 == 32'h4;
  assign T123 = io_inst & 32'h4;
  assign T124 = T127 | T125;
  assign T125 = T126 == 32'h10000010;
  assign T126 = io_inst & 32'h10000010;
  assign T127 = T128 == 32'h8;
  assign T128 = io_inst & 32'h8;
  assign T129 = T132 | T130;
  assign T130 = T131 == 32'h20000000;
  assign T131 = io_inst & 32'h20000000;
  assign T132 = T133 == 32'h0;
  assign T133 = io_inst & 32'h40;
  assign T134 = T132 | T135;
  assign T135 = T136 == 32'h40000000;
  assign T136 = io_inst & 32'h40000000;
  assign T137 = T138 == 32'h0;
  assign T138 = io_inst & 32'h10;
endmodule

module mulAddSubRecodedFloatN_0(
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output[32:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire roundInexact;
  wire anyRound;
  wire T4;
  wire[27:0] T5;
  wire[27:0] T6;
  wire[25:0] T7;
  wire[26:0] roundMask;
  wire[26:0] T8;
  wire[24:0] T9;
  wire[24:0] T10;
  wire T11;
  wire[27:0] T12;
  wire[42:0] T13;
  wire T14;
  wire T15;
  wire[15:0] T16;
  wire[15:0] absSigSumExtraMask;
  wire[14:0] T17;
  wire[6:0] T18;
  wire[2:0] T19;
  wire T20;
  wire[2:0] T21;
  wire[6:0] T22;
  wire[14:0] T23;
  wire[16:0] T24;
  wire[3:0] normTo2ShiftDist;
  wire[3:0] estNormDist_5;
  wire[3:0] T25;
  wire[6:0] estNormDist;
  wire[6:0] T26;
  wire[6:0] estNormPos_dist;
  wire[6:0] T27;
  wire[6:0] T28;
  wire[6:0] T29;
  wire[6:0] T30;
  wire[6:0] T31;
  wire[6:0] T32;
  wire[6:0] T33;
  wire[6:0] T34;
  wire[6:0] T35;
  wire[6:0] T36;
  wire[6:0] T37;
  wire[6:0] T38;
  wire[6:0] T39;
  wire[6:0] T40;
  wire[6:0] T41;
  wire[6:0] T42;
  wire[6:0] T43;
  wire[6:0] T44;
  wire[6:0] T45;
  wire[6:0] T46;
  wire[6:0] T47;
  wire[6:0] T48;
  wire[6:0] T49;
  wire[6:0] T50;
  wire[6:0] T51;
  wire[6:0] T52;
  wire[6:0] T53;
  wire[6:0] T54;
  wire[6:0] T55;
  wire[6:0] T56;
  wire[6:0] T57;
  wire[6:0] T58;
  wire[6:0] T59;
  wire[6:0] T60;
  wire[6:0] T61;
  wire[6:0] T62;
  wire[6:0] T63;
  wire[6:0] T64;
  wire[6:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[6:0] T68;
  wire[6:0] T69;
  wire[6:0] T70;
  wire[6:0] T71;
  wire[6:0] T72;
  wire[6:0] T73;
  wire[6:0] T74;
  wire T75;
  wire[50:0] T76;
  wire[50:0] T77;
  wire[49:0] T78;
  wire[49:0] T79;
  wire[74:0] sigSum;
  wire[74:0] T80;
  wire[75:0] T81;
  wire T82;
  wire doSubMags;
  wire opSignC;
  wire T83;
  wire T84;
  wire signProd;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire[23:0] T90;
  wire[23:0] CExtraMask;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[6:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[5:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[3:0] T102;
  wire[7:0] T103;
  wire[23:0] T104;
  wire[128:0] T105;
  wire[6:0] T106;
  wire[10:0] T107;
  wire[10:0] T108;
  wire[10:0] sNatCAlignDist;
  wire[10:0] T109;
  wire[8:0] T110;
  wire[10:0] sExpAlignedProd;
  wire[10:0] T111;
  wire[10:0] T112;
  wire[8:0] T113;
  wire[10:0] T114;
  wire[7:0] T115;
  wire[8:0] T116;
  wire[2:0] T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire[9:0] T122;
  wire CAlignDist_floor;
  wire T123;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T124;
  wire isZeroA;
  wire[2:0] T125;
  wire[7:0] T126;
  wire[7:0] T127;
  wire[3:0] T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[5:0] T131;
  wire[7:0] T132;
  wire[7:0] T133;
  wire[6:0] T134;
  wire[15:0] T135;
  wire[15:0] T136;
  wire[15:0] T137;
  wire[14:0] T138;
  wire[15:0] T139;
  wire[15:0] T140;
  wire[15:0] T141;
  wire[13:0] T142;
  wire[15:0] T143;
  wire[15:0] T144;
  wire[15:0] T145;
  wire[11:0] T146;
  wire[15:0] T147;
  wire[15:0] T148;
  wire[15:0] T149;
  wire[7:0] T150;
  wire[15:0] T151;
  wire[15:0] T152;
  wire[15:0] T153;
  wire[7:0] T154;
  wire[15:0] T155;
  wire[15:0] T156;
  wire[11:0] T157;
  wire[15:0] T158;
  wire[15:0] T159;
  wire[13:0] T160;
  wire[15:0] T161;
  wire[15:0] T162;
  wire[14:0] T163;
  wire[23:0] sigC;
  wire[22:0] T164;
  wire T165;
  wire isZeroC;
  wire[2:0] T166;
  wire[74:0] T167;
  wire[74:0] T168;
  wire[74:0] T169;
  wire[73:0] T170;
  wire[49:0] T171;
  wire[49:0] T172;
  wire[23:0] negSigC;
  wire[23:0] T173;
  wire[74:0] T174;
  wire[48:0] T175;
  wire[47:0] T176;
  wire[23:0] sigB;
  wire[22:0] T177;
  wire T178;
  wire[23:0] sigA;
  wire[22:0] T179;
  wire T180;
  wire[50:0] T181;
  wire[49:0] T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire[6:0] CDom_estNormDist;
  wire[6:0] T232;
  wire[4:0] T233;
  wire[6:0] T234;
  wire T235;
  wire CAlignDist_0;
  wire T236;
  wire[9:0] T237;
  wire isCDominant;
  wire T238;
  wire T239;
  wire[9:0] T240;
  wire T241;
  wire[1:0] T242;
  wire T243;
  wire[1:0] T244;
  wire T245;
  wire[3:0] T246;
  wire[1:0] T247;
  wire T248;
  wire[1:0] T249;
  wire[3:0] T250;
  wire T251;
  wire[1:0] T252;
  wire T253;
  wire[1:0] T254;
  wire T255;
  wire[7:0] T256;
  wire[7:0] T257;
  wire[7:0] T258;
  wire[6:0] T259;
  wire[7:0] T260;
  wire[7:0] T261;
  wire[7:0] T262;
  wire[5:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[7:0] T266;
  wire[3:0] T267;
  wire[7:0] T268;
  wire[7:0] T269;
  wire[7:0] T270;
  wire[3:0] T271;
  wire[7:0] T272;
  wire[7:0] T273;
  wire[5:0] T274;
  wire[7:0] T275;
  wire[7:0] T276;
  wire[6:0] T277;
  wire[15:0] T278;
  wire[42:0] cFirstNormAbsSigSum;
  wire[42:0] T279;
  wire[41:0] T280;
  wire[41:0] notCDom_pos_firstNormAbsSigSum;
  wire[41:0] T281;
  wire[41:0] T282;
  wire[31:0] T283;
  wire[31:0] T284;
  wire[9:0] T285;
  wire[41:0] T286;
  wire[33:0] T287;
  wire T288;
  wire T289;
  wire[1:0] firstReduceSigSum;
  wire T290;
  wire[17:0] T291;
  wire T292;
  wire[15:0] T293;
  wire T294;
  wire T295;
  wire[1:0] firstReduceNotSigSum;
  wire T296;
  wire[17:0] T297;
  wire[74:0] notSigSum;
  wire T298;
  wire[15:0] T299;
  wire[32:0] T300;
  wire T301;
  wire[41:0] T302;
  wire[41:0] T303;
  wire[41:0] T304;
  wire[15:0] T305;
  wire[15:0] T306;
  wire[25:0] T307;
  wire T308;
  wire T309;
  wire[41:0] CDom_firstNormAbsSigSum;
  wire[41:0] T310;
  wire[41:0] T311;
  wire[41:0] T312;
  wire T313;
  wire[40:0] T314;
  wire[41:0] T315;
  wire T316;
  wire T317;
  wire T318;
  wire[41:0] T319;
  wire[41:0] T320;
  wire[41:0] T321;
  wire T322;
  wire[40:0] T323;
  wire[41:0] T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire[41:0] T329;
  wire[41:0] T330;
  wire[41:0] T331;
  wire T332;
  wire[40:0] T333;
  wire[41:0] T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire[41:0] T339;
  wire[41:0] T340;
  wire T341;
  wire[40:0] T342;
  wire[41:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire[42:0] T349;
  wire[42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[42:0] T350;
  wire[42:0] T351;
  wire[10:0] T352;
  wire[42:0] T353;
  wire[32:0] T354;
  wire T355;
  wire[31:0] T356;
  wire T357;
  wire[42:0] T358;
  wire[42:0] T359;
  wire[41:0] T360;
  wire[42:0] T361;
  wire[26:0] T362;
  wire T363;
  wire T364;
  wire[42:0] T365;
  wire T366;
  wire[15:0] T367;
  wire[15:0] T368;
  wire[15:0] T369;
  wire doIncrSig;
  wire T370;
  wire T371;
  wire T372;
  wire[41:0] T373;
  wire[41:0] T374;
  wire[24:0] T375;
  wire[8:0] T376;
  wire T377;
  wire[8:0] T378;
  wire[24:0] T379;
  wire[1024:0] T380;
  wire[9:0] T381;
  wire[9:0] T382;
  wire[10:0] sExpX3;
  wire[10:0] T383;
  wire[10:0] sExpSum;
  wire[10:0] T384;
  wire[7:0] T385;
  wire[7:0] T386;
  wire[7:0] T387;
  wire[6:0] T388;
  wire[7:0] T389;
  wire[7:0] T390;
  wire[7:0] T391;
  wire[5:0] T392;
  wire[7:0] T393;
  wire[7:0] T394;
  wire[7:0] T395;
  wire[3:0] T396;
  wire[7:0] T397;
  wire[7:0] T398;
  wire[7:0] T399;
  wire[3:0] T400;
  wire[7:0] T401;
  wire[7:0] T402;
  wire[5:0] T403;
  wire[7:0] T404;
  wire[7:0] T405;
  wire[6:0] T406;
  wire[15:0] T407;
  wire[15:0] T408;
  wire[15:0] T409;
  wire[14:0] T410;
  wire[15:0] T411;
  wire[15:0] T412;
  wire[15:0] T413;
  wire[13:0] T414;
  wire[15:0] T415;
  wire[15:0] T416;
  wire[15:0] T417;
  wire[11:0] T418;
  wire[15:0] T419;
  wire[15:0] T420;
  wire[15:0] T421;
  wire[7:0] T422;
  wire[15:0] T423;
  wire[15:0] T424;
  wire[15:0] T425;
  wire[7:0] T426;
  wire[15:0] T427;
  wire[15:0] T428;
  wire[11:0] T429;
  wire[15:0] T430;
  wire[15:0] T431;
  wire[13:0] T432;
  wire[15:0] T433;
  wire[15:0] T434;
  wire[14:0] T435;
  wire[26:0] T436;
  wire[26:0] T437;
  wire T438;
  wire T439;
  wire[27:0] T440;
  wire[27:0] T441;
  wire[26:0] roundPosMask;
  wire[26:0] T442;
  wire[25:0] T443;
  wire[25:0] T444;
  wire T445;
  wire allRound;
  wire allRoundExtra;
  wire[27:0] T446;
  wire[27:0] T447;
  wire[25:0] T448;
  wire[27:0] T449;
  wire commonCase;
  wire T450;
  wire notSpecial_addZeros;
  wire T451;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T452;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T453;
  wire isSpecialA;
  wire[1:0] T454;
  wire overflow;
  wire overflowY;
  wire[2:0] T455;
  wire[10:0] sExpY;
  wire[10:0] T456;
  wire[10:0] T457;
  wire T458;
  wire[1:0] T459;
  wire[25:0] sigY3;
  wire[25:0] T460;
  wire[25:0] T461;
  wire[25:0] T462;
  wire[25:0] T463;
  wire[25:0] T464;
  wire[25:0] T465;
  wire[25:0] T466;
  wire[27:0] T467;
  wire[27:0] T468;
  wire roundEven;
  wire T469;
  wire T470;
  wire T471;
  wire roundingMode_nearest_even;
  wire T472;
  wire T473;
  wire T474;
  wire[25:0] T475;
  wire[25:0] T476;
  wire roundUp;
  wire T477;
  wire T478;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T479;
  wire doNegSignSum;
  wire T480;
  wire T481;
  wire T482;
  wire isZeroY;
  wire[2:0] T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire[25:0] T497;
  wire[25:0] T498;
  wire[27:0] T499;
  wire[27:0] T500;
  wire[26:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[10:0] T505;
  wire[10:0] T506;
  wire T507;
  wire[10:0] T508;
  wire[10:0] T509;
  wire T510;
  wire underflow;
  wire underflowY;
  wire T511;
  wire T512;
  wire[9:0] T513;
  wire[7:0] T514;
  wire sigX3Shift1;
  wire[1:0] T515;
  wire T516;
  wire[1:0] T517;
  wire invalid;
  wire notSigNaN_invalid;
  wire T518;
  wire T519;
  wire isInfC;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire isInfB;
  wire T524;
  wire T525;
  wire isInfA;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire isNaNB;
  wire T530;
  wire T531;
  wire isNaNA;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire isSigNaNC;
  wire T537;
  wire T538;
  wire isNaNC;
  wire T539;
  wire T540;
  wire isSigNaNB;
  wire T541;
  wire T542;
  wire isSigNaNA;
  wire T543;
  wire T544;
  wire[32:0] T545;
  wire[31:0] T546;
  wire[22:0] fractOut;
  wire[22:0] T547;
  wire[22:0] T548;
  wire T549;
  wire isSatOut;
  wire T550;
  wire overflowY_roundMagUp;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire isNaNOut;
  wire T555;
  wire T556;
  wire[22:0] fractY;
  wire[22:0] T557;
  wire[22:0] T558;
  wire[8:0] expOut;
  wire[8:0] T559;
  wire[8:0] T560;
  wire[8:0] T561;
  wire notNaN_isInfOut;
  wire T562;
  wire T563;
  wire T564;
  wire[8:0] T565;
  wire[8:0] T566;
  wire[8:0] T567;
  wire[8:0] T568;
  wire[8:0] T569;
  wire[8:0] T570;
  wire[8:0] T571;
  wire[8:0] T572;
  wire[8:0] T573;
  wire[8:0] T574;
  wire[8:0] T575;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T576;
  wire[8:0] T577;
  wire T578;
  wire T579;
  wire[8:0] T580;
  wire signOut;
  wire T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;


  assign io_exceptionFlags = T0;
  assign T0 = {T517, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & roundInexact;
  assign roundInexact = doIncrSig ? T445 : anyRound;
  assign anyRound = T439 | T4;
  assign T4 = T5 != 28'h0;
  assign T5 = T12 & T6;
  assign T6 = {2'h0, T7};
  assign T7 = roundMask >> 1'h1;
  assign roundMask = T436 | T8;
  assign T8 = {T9, 2'h3};
  assign T9 = T375 | T10;
  assign T10 = {24'h0, T11};
  assign T11 = T12[5'h1a:5'h1a];
  assign T12 = T13[5'h1b:1'h0];
  assign T13 = {T373, T14};
  assign T14 = doIncrSig ? T366 : T15;
  assign T15 = T16 != 16'h0;
  assign T16 = T278 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T17, 1'h1};
  assign T17 = {T256, T18};
  assign T18 = {T246, T19};
  assign T19 = {T242, T20};
  assign T20 = T21[2'h2:2'h2];
  assign T21 = T22[3'h6:3'h4];
  assign T22 = T23[4'he:4'h8];
  assign T23 = T24[4'hf:1'h1];
  assign T24 = $signed(17'h10000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T25;
  assign T25 = estNormDist[2'h3:1'h0];
  assign estNormDist = isCDominant ? CDom_estNormDist : T26;
  assign T26 = T231 ? estNormPos_dist : estNormPos_dist;
  assign estNormPos_dist = T230 ? 7'h18 : T27;
  assign T27 = T229 ? 7'h19 : T28;
  assign T28 = T228 ? 7'h1a : T29;
  assign T29 = T227 ? 7'h1b : T30;
  assign T30 = T226 ? 7'h1c : T31;
  assign T31 = T225 ? 7'h1d : T32;
  assign T32 = T224 ? 7'h1e : T33;
  assign T33 = T223 ? 7'h1f : T34;
  assign T34 = T222 ? 7'h20 : T35;
  assign T35 = T221 ? 7'h21 : T36;
  assign T36 = T220 ? 7'h22 : T37;
  assign T37 = T219 ? 7'h23 : T38;
  assign T38 = T218 ? 7'h24 : T39;
  assign T39 = T217 ? 7'h25 : T40;
  assign T40 = T216 ? 7'h26 : T41;
  assign T41 = T215 ? 7'h27 : T42;
  assign T42 = T214 ? 7'h28 : T43;
  assign T43 = T213 ? 7'h29 : T44;
  assign T44 = T212 ? 7'h2a : T45;
  assign T45 = T211 ? 7'h2b : T46;
  assign T46 = T210 ? 7'h2c : T47;
  assign T47 = T209 ? 7'h2d : T48;
  assign T48 = T208 ? 7'h2e : T49;
  assign T49 = T207 ? 7'h2f : T50;
  assign T50 = T206 ? 7'h30 : T51;
  assign T51 = T205 ? 7'h31 : T52;
  assign T52 = T204 ? 7'h32 : T53;
  assign T53 = T203 ? 7'h33 : T54;
  assign T54 = T202 ? 7'h34 : T55;
  assign T55 = T201 ? 7'h35 : T56;
  assign T56 = T200 ? 7'h36 : T57;
  assign T57 = T199 ? 7'h37 : T58;
  assign T58 = T198 ? 7'h38 : T59;
  assign T59 = T197 ? 7'h39 : T60;
  assign T60 = T196 ? 7'h3a : T61;
  assign T61 = T195 ? 7'h3b : T62;
  assign T62 = T194 ? 7'h3c : T63;
  assign T63 = T193 ? 7'h3d : T64;
  assign T64 = T192 ? 7'h3e : T65;
  assign T65 = T191 ? 7'h3f : T66;
  assign T66 = T190 ? 7'h40 : T67;
  assign T67 = T189 ? 7'h41 : T68;
  assign T68 = T188 ? 7'h42 : T69;
  assign T69 = T187 ? 7'h43 : T70;
  assign T70 = T186 ? 7'h44 : T71;
  assign T71 = T185 ? 7'h45 : T72;
  assign T72 = T184 ? 7'h46 : T73;
  assign T73 = T183 ? 7'h47 : T74;
  assign T74 = T75 ? 7'h48 : 7'h49;
  assign T75 = T76[1'h1:1'h1];
  assign T76 = T181 ^ T77;
  assign T77 = T78 << 1'h1;
  assign T78 = 50'h0 | T79;
  assign T79 = sigSum[6'h32:1'h1];
  assign sigSum = T174 + T80;
  assign T80 = T81[7'h4a:1'h0];
  assign T81 = {T167, T82};
  assign T82 = T89 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T84 ^ T83;
  assign T83 = io_op[1'h0:1'h0];
  assign T84 = io_c[6'h20:6'h20];
  assign signProd = T86 ^ T85;
  assign T85 = io_op[1'h1:1'h1];
  assign T86 = T88 ^ T87;
  assign T87 = io_b[6'h20:6'h20];
  assign T88 = io_a[6'h20:6'h20];
  assign T89 = T90 != 24'h0;
  assign T90 = sigC & CExtraMask;
  assign CExtraMask = {T135, T91};
  assign T91 = T132 | T92;
  assign T92 = T93 & 8'haa;
  assign T93 = T94 << 1'h1;
  assign T94 = T95[3'h6:1'h0];
  assign T95 = T129 | T96;
  assign T96 = T97 & 8'hcc;
  assign T97 = T98 << 2'h2;
  assign T98 = T99[3'h5:1'h0];
  assign T99 = T126 | T100;
  assign T100 = T101 & 8'hf0;
  assign T101 = T102 << 3'h4;
  assign T102 = T103[2'h3:1'h0];
  assign T103 = T104[5'h17:5'h10];
  assign T104 = T105[7'h4d:6'h36];
  assign T105 = $signed(129'h100000000000000000000000000000000) >>> T106;
  assign T106 = T107[3'h6:1'h0];
  assign T107 = CAlignDist_floor ? 11'h0 : T108;
  assign T108 = T121 ? sNatCAlignDist : 11'h4a;
  assign sNatCAlignDist = sExpAlignedProd - T109;
  assign T109 = {2'h0, T110};
  assign T110 = io_c[5'h1f:5'h17];
  assign sExpAlignedProd = T111 + 11'h1b;
  assign T111 = T114 + T112;
  assign T112 = {2'h0, T113};
  assign T113 = io_a[5'h1f:5'h17];
  assign T114 = {T117, T115};
  assign T115 = T116[3'h7:1'h0];
  assign T116 = io_b[5'h1f:5'h17];
  assign T117 = 3'h0 - T118;
  assign T118 = {2'h0, T119};
  assign T119 = T120 ^ 1'h1;
  assign T120 = T116[4'h8:4'h8];
  assign T121 = T122 < 10'h4a;
  assign T122 = sNatCAlignDist[4'h9:1'h0];
  assign CAlignDist_floor = isZeroProd | T123;
  assign T123 = sNatCAlignDist[4'ha:4'ha];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T124 == 3'h0;
  assign T124 = T116[4'h8:3'h6];
  assign isZeroA = T125 == 3'h0;
  assign T125 = T113[4'h8:3'h6];
  assign T126 = T127 & 8'hf;
  assign T127 = {4'h0, T128};
  assign T128 = T103 >> 3'h4;
  assign T129 = T130 & 8'h33;
  assign T130 = {2'h0, T131};
  assign T131 = T99 >> 2'h2;
  assign T132 = T133 & 8'h55;
  assign T133 = {1'h0, T134};
  assign T134 = T95 >> 1'h1;
  assign T135 = T161 | T136;
  assign T136 = T137 & 16'haaaa;
  assign T137 = T138 << 1'h1;
  assign T138 = T139[4'he:1'h0];
  assign T139 = T158 | T140;
  assign T140 = T141 & 16'hcccc;
  assign T141 = T142 << 2'h2;
  assign T142 = T143[4'hd:1'h0];
  assign T143 = T155 | T144;
  assign T144 = T145 & 16'hf0f0;
  assign T145 = T146 << 3'h4;
  assign T146 = T147[4'hb:1'h0];
  assign T147 = T152 | T148;
  assign T148 = T149 & 16'hff00;
  assign T149 = T150 << 4'h8;
  assign T150 = T151[3'h7:1'h0];
  assign T151 = T104[4'hf:1'h0];
  assign T152 = T153 & 16'hff;
  assign T153 = {8'h0, T154};
  assign T154 = T151 >> 4'h8;
  assign T155 = T156 & 16'hf0f;
  assign T156 = {4'h0, T157};
  assign T157 = T147 >> 3'h4;
  assign T158 = T159 & 16'h3333;
  assign T159 = {2'h0, T160};
  assign T160 = T143 >> 2'h2;
  assign T161 = T162 & 16'h5555;
  assign T162 = {1'h0, T163};
  assign T163 = T139 >> 1'h1;
  assign sigC = {T165, T164};
  assign T164 = io_c[5'h16:1'h0];
  assign T165 = isZeroC ^ 1'h1;
  assign isZeroC = T166 == 3'h0;
  assign T166 = T110[4'h8:3'h6];
  assign T167 = $signed(T168) >>> T106;
  assign T168 = T169;
  assign T169 = {doSubMags, T170};
  assign T170 = {negSigC, T171};
  assign T171 = 50'h0 - T172;
  assign T172 = {49'h0, doSubMags};
  assign negSigC = doSubMags ? T173 : sigC;
  assign T173 = ~ sigC;
  assign T174 = {26'h0, T175};
  assign T175 = T176 << 1'h1;
  assign T176 = sigA * sigB;
  assign sigB = {T178, T177};
  assign T177 = io_b[5'h16:1'h0];
  assign T178 = isZeroB ^ 1'h1;
  assign sigA = {T180, T179};
  assign T179 = io_a[5'h16:1'h0];
  assign T180 = isZeroA ^ 1'h1;
  assign T181 = {1'h0, T182};
  assign T182 = 50'h0 ^ T79;
  assign T183 = T76[2'h2:2'h2];
  assign T184 = T76[2'h3:2'h3];
  assign T185 = T76[3'h4:3'h4];
  assign T186 = T76[3'h5:3'h5];
  assign T187 = T76[3'h6:3'h6];
  assign T188 = T76[3'h7:3'h7];
  assign T189 = T76[4'h8:4'h8];
  assign T190 = T76[4'h9:4'h9];
  assign T191 = T76[4'ha:4'ha];
  assign T192 = T76[4'hb:4'hb];
  assign T193 = T76[4'hc:4'hc];
  assign T194 = T76[4'hd:4'hd];
  assign T195 = T76[4'he:4'he];
  assign T196 = T76[4'hf:4'hf];
  assign T197 = T76[5'h10:5'h10];
  assign T198 = T76[5'h11:5'h11];
  assign T199 = T76[5'h12:5'h12];
  assign T200 = T76[5'h13:5'h13];
  assign T201 = T76[5'h14:5'h14];
  assign T202 = T76[5'h15:5'h15];
  assign T203 = T76[5'h16:5'h16];
  assign T204 = T76[5'h17:5'h17];
  assign T205 = T76[5'h18:5'h18];
  assign T206 = T76[5'h19:5'h19];
  assign T207 = T76[5'h1a:5'h1a];
  assign T208 = T76[5'h1b:5'h1b];
  assign T209 = T76[5'h1c:5'h1c];
  assign T210 = T76[5'h1d:5'h1d];
  assign T211 = T76[5'h1e:5'h1e];
  assign T212 = T76[5'h1f:5'h1f];
  assign T213 = T76[6'h20:6'h20];
  assign T214 = T76[6'h21:6'h21];
  assign T215 = T76[6'h22:6'h22];
  assign T216 = T76[6'h23:6'h23];
  assign T217 = T76[6'h24:6'h24];
  assign T218 = T76[6'h25:6'h25];
  assign T219 = T76[6'h26:6'h26];
  assign T220 = T76[6'h27:6'h27];
  assign T221 = T76[6'h28:6'h28];
  assign T222 = T76[6'h29:6'h29];
  assign T223 = T76[6'h2a:6'h2a];
  assign T224 = T76[6'h2b:6'h2b];
  assign T225 = T76[6'h2c:6'h2c];
  assign T226 = T76[6'h2d:6'h2d];
  assign T227 = T76[6'h2e:6'h2e];
  assign T228 = T76[6'h2f:6'h2f];
  assign T229 = T76[6'h30:6'h30];
  assign T230 = T76[6'h31:6'h31];
  assign T231 = sigSum[6'h33:6'h33];
  assign CDom_estNormDist = T235 ? T106 : T232;
  assign T232 = {2'h0, T233};
  assign T233 = T234[3'h4:1'h0];
  assign T234 = T106 - 7'h1;
  assign T235 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T236;
  assign T236 = T237 == 10'h0;
  assign T237 = sNatCAlignDist[4'h9:1'h0];
  assign isCDominant = T241 & T238;
  assign T238 = CAlignDist_floor | T239;
  assign T239 = T240 < 10'h19;
  assign T240 = sNatCAlignDist[4'h9:1'h0];
  assign T241 = isZeroC ^ 1'h1;
  assign T242 = {T245, T243};
  assign T243 = T244[1'h1:1'h1];
  assign T244 = T21[1'h1:1'h0];
  assign T245 = T244[1'h0:1'h0];
  assign T246 = {T252, T247};
  assign T247 = {T251, T248};
  assign T248 = T249[1'h1:1'h1];
  assign T249 = T250[2'h3:2'h2];
  assign T250 = T22[2'h3:1'h0];
  assign T251 = T249[1'h0:1'h0];
  assign T252 = {T255, T253};
  assign T253 = T254[1'h1:1'h1];
  assign T254 = T250[1'h1:1'h0];
  assign T255 = T254[1'h0:1'h0];
  assign T256 = T275 | T257;
  assign T257 = T258 & 8'haa;
  assign T258 = T259 << 1'h1;
  assign T259 = T260[3'h6:1'h0];
  assign T260 = T272 | T261;
  assign T261 = T262 & 8'hcc;
  assign T262 = T263 << 2'h2;
  assign T263 = T264[3'h5:1'h0];
  assign T264 = T269 | T265;
  assign T265 = T266 & 8'hf0;
  assign T266 = T267 << 3'h4;
  assign T267 = T268[2'h3:1'h0];
  assign T268 = T23[3'h7:1'h0];
  assign T269 = T270 & 8'hf;
  assign T270 = {4'h0, T271};
  assign T271 = T268 >> 3'h4;
  assign T272 = T273 & 8'h33;
  assign T273 = {2'h0, T274};
  assign T274 = T264 >> 2'h2;
  assign T275 = T276 & 8'h55;
  assign T276 = {1'h0, T277};
  assign T277 = T260 >> 1'h1;
  assign T278 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign cFirstNormAbsSigSum = T231 ? T349 : T279;
  assign T279 = {1'h0, T280};
  assign T280 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T309 ? T302 : T281;
  assign T281 = T301 ? T286 : T282;
  assign T282 = {T285, T283};
  assign T283 = 32'h0 - T284;
  assign T284 = {31'h0, doSubMags};
  assign T285 = sigSum[4'ha:1'h1];
  assign T286 = {8'h0, T287};
  assign T287 = {T300, T288};
  assign T288 = doSubMags ? T294 : T289;
  assign T289 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T292, T290};
  assign T290 = T291 != 18'h0;
  assign T291 = sigSum[5'h11:1'h0];
  assign T292 = T293 != 16'h0;
  assign T293 = sigSum[6'h21:5'h12];
  assign T294 = ~ T295;
  assign T295 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T298, T296};
  assign T296 = T297 != 18'h0;
  assign T297 = notSigSum[5'h11:1'h0];
  assign notSigSum = ~ sigSum;
  assign T298 = T299 != 16'h0;
  assign T299 = notSigSum[6'h21:5'h12];
  assign T300 = sigSum[6'h32:5'h12];
  assign T301 = estNormPos_dist[3'h4:3'h4];
  assign T302 = T308 ? T304 : T303;
  assign T303 = sigSum[6'h2a:1'h1];
  assign T304 = {T307, T305};
  assign T305 = 16'h0 - T306;
  assign T306 = {15'h0, doSubMags};
  assign T307 = sigSum[5'h1a:1'h1];
  assign T308 = estNormPos_dist[3'h4:3'h4];
  assign T309 = estNormPos_dist[3'h5:3'h5];
  assign CDom_firstNormAbsSigSum = T310;
  assign T310 = T319 | T311;
  assign T311 = T315 & T312;
  assign T312 = {T314, T313};
  assign T313 = firstReduceNotSigSum[1'h0:1'h0];
  assign T314 = notSigSum[6'h3a:5'h12];
  assign T315 = T316 ? 42'h3ffffffffff : 42'h0;
  assign T316 = T317;
  assign T317 = doSubMags & T318;
  assign T318 = CDom_estNormDist[3'h4:3'h4];
  assign T319 = T329 | T320;
  assign T320 = T324 & T321;
  assign T321 = {T323, T322};
  assign T322 = firstReduceNotSigSum != 2'h0;
  assign T323 = notSigSum[7'h4a:6'h22];
  assign T324 = T325 ? 42'h3ffffffffff : 42'h0;
  assign T325 = T326;
  assign T326 = doSubMags & T327;
  assign T327 = ~ T328;
  assign T328 = CDom_estNormDist[3'h4:3'h4];
  assign T329 = T339 | T330;
  assign T330 = T334 & T331;
  assign T331 = {T333, T332};
  assign T332 = firstReduceSigSum[1'h0:1'h0];
  assign T333 = sigSum[6'h3a:5'h12];
  assign T334 = T335 ? 42'h3ffffffffff : 42'h0;
  assign T335 = T336;
  assign T336 = T338 & T337;
  assign T337 = CDom_estNormDist[3'h4:3'h4];
  assign T338 = ~ doSubMags;
  assign T339 = T343 & T340;
  assign T340 = {T342, T341};
  assign T341 = firstReduceSigSum != 2'h0;
  assign T342 = sigSum[7'h4a:6'h22];
  assign T343 = T344 ? 42'h3ffffffffff : 42'h0;
  assign T344 = T345;
  assign T345 = T348 & T346;
  assign T346 = ~ T347;
  assign T347 = CDom_estNormDist[3'h4:3'h4];
  assign T348 = ~ doSubMags;
  assign T349 = isCDominant ? T365 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T364 ? T358 : T350;
  assign T350 = T357 ? T353 : T351;
  assign T351 = T352 << 6'h20;
  assign T352 = notSigSum[4'hb:1'h1];
  assign T353 = {10'h0, T354};
  assign T354 = {T356, T355};
  assign T355 = firstReduceNotSigSum[1'h0:1'h0];
  assign T356 = notSigSum[6'h31:5'h12];
  assign T357 = estNormPos_dist[3'h4:3'h4];
  assign T358 = T363 ? T361 : T359;
  assign T359 = {1'h0, T360};
  assign T360 = notSigSum[6'h2a:1'h1];
  assign T361 = T362 << 5'h10;
  assign T362 = notSigSum[5'h1b:1'h1];
  assign T363 = estNormPos_dist[3'h4:3'h4];
  assign T364 = estNormPos_dist[3'h5:3'h5];
  assign T365 = {1'h0, CDom_firstNormAbsSigSum};
  assign T366 = T367 == 16'h0;
  assign T367 = T368 & absSigSumExtraMask;
  assign T368 = ~ T369;
  assign T369 = cFirstNormAbsSigSum[4'hf:1'h0];
  assign doIncrSig = T370 & doSubMags;
  assign T370 = T372 & T371;
  assign T371 = ~ T231;
  assign T372 = ~ isCDominant;
  assign T373 = T374 >> normTo2ShiftDist;
  assign T374 = cFirstNormAbsSigSum[6'h2a:1'h1];
  assign T375 = {T407, T376};
  assign T376 = {T385, T377};
  assign T377 = T378[4'h8:4'h8];
  assign T378 = T379[5'h18:5'h10];
  assign T379 = T380[8'h83:7'h6b];
  assign T380 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T381;
  assign T381 = ~ T382;
  assign T382 = sExpX3[4'h9:1'h0];
  assign sExpX3 = sExpSum - T383;
  assign T383 = {4'h0, estNormDist};
  assign sExpSum = CAlignDist_floor ? T384 : sExpAlignedProd;
  assign T384 = {2'h0, T110};
  assign T385 = T404 | T386;
  assign T386 = T387 & 8'haa;
  assign T387 = T388 << 1'h1;
  assign T388 = T389[3'h6:1'h0];
  assign T389 = T401 | T390;
  assign T390 = T391 & 8'hcc;
  assign T391 = T392 << 2'h2;
  assign T392 = T393[3'h5:1'h0];
  assign T393 = T398 | T394;
  assign T394 = T395 & 8'hf0;
  assign T395 = T396 << 3'h4;
  assign T396 = T397[2'h3:1'h0];
  assign T397 = T378[3'h7:1'h0];
  assign T398 = T399 & 8'hf;
  assign T399 = {4'h0, T400};
  assign T400 = T397 >> 3'h4;
  assign T401 = T402 & 8'h33;
  assign T402 = {2'h0, T403};
  assign T403 = T393 >> 2'h2;
  assign T404 = T405 & 8'h55;
  assign T405 = {1'h0, T406};
  assign T406 = T389 >> 1'h1;
  assign T407 = T433 | T408;
  assign T408 = T409 & 16'haaaa;
  assign T409 = T410 << 1'h1;
  assign T410 = T411[4'he:1'h0];
  assign T411 = T430 | T412;
  assign T412 = T413 & 16'hcccc;
  assign T413 = T414 << 2'h2;
  assign T414 = T415[4'hd:1'h0];
  assign T415 = T427 | T416;
  assign T416 = T417 & 16'hf0f0;
  assign T417 = T418 << 3'h4;
  assign T418 = T419[4'hb:1'h0];
  assign T419 = T424 | T420;
  assign T420 = T421 & 16'hff00;
  assign T421 = T422 << 4'h8;
  assign T422 = T423[3'h7:1'h0];
  assign T423 = T379[4'hf:1'h0];
  assign T424 = T425 & 16'hff;
  assign T425 = {8'h0, T426};
  assign T426 = T423 >> 4'h8;
  assign T427 = T428 & 16'hf0f;
  assign T428 = {4'h0, T429};
  assign T429 = T419 >> 3'h4;
  assign T430 = T431 & 16'h3333;
  assign T431 = {2'h0, T432};
  assign T432 = T415 >> 2'h2;
  assign T433 = T434 & 16'h5555;
  assign T434 = {1'h0, T435};
  assign T435 = T411 >> 1'h1;
  assign T436 = 27'h0 - T437;
  assign T437 = {26'h0, T438};
  assign T438 = sExpX3[4'ha:4'ha];
  assign T439 = T440 != 28'h0;
  assign T440 = T12 & T441;
  assign T441 = {1'h0, roundPosMask};
  assign roundPosMask = T442 & roundMask;
  assign T442 = {1'h0, T443};
  assign T443 = ~ T444;
  assign T444 = roundMask >> 1'h1;
  assign T445 = ~ allRound;
  assign allRound = T439 & allRoundExtra;
  assign allRoundExtra = T446 == 28'h0;
  assign T446 = T449 & T447;
  assign T447 = {2'h0, T448};
  assign T448 = roundMask >> 1'h1;
  assign T449 = ~ T12;
  assign commonCase = T451 & T450;
  assign T450 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T451 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T452 == 2'h3;
  assign T452 = T110[4'h8:3'h7];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T453 == 2'h3;
  assign T453 = T116[4'h8:3'h7];
  assign isSpecialA = T454 == 2'h3;
  assign T454 = T113[4'h8:3'h7];
  assign overflow = commonCase & overflowY;
  assign overflowY = T455 == 3'h3;
  assign T455 = sExpY[4'h9:3'h7];
  assign sExpY = T505 | T456;
  assign T456 = T458 ? T457 : 11'h0;
  assign T457 = sExpX3 - 11'h1;
  assign T458 = T459 == 2'h0;
  assign T459 = sigY3[5'h19:5'h18];
  assign sigY3 = T475 | T460;
  assign T460 = roundEven ? T461 : 26'h0;
  assign T461 = T464 & T462;
  assign T462 = ~ T463;
  assign T463 = roundMask >> 1'h1;
  assign T464 = T465[5'h19:1'h0];
  assign T465 = T466 + 26'h1;
  assign T466 = T467 >> 2'h2;
  assign T467 = T12 | T468;
  assign T468 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T472 : T469;
  assign T469 = T471 & T470;
  assign T470 = ~ T4;
  assign T471 = roundingMode_nearest_even & T439;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T472 = T473 & allRoundExtra;
  assign T473 = roundingMode_nearest_even & T474;
  assign T474 = ~ T439;
  assign T475 = T497 | T476;
  assign T476 = roundUp ? T464 : 26'h0;
  assign roundUp = T484 | T477;
  assign T477 = T478 & 1'h1;
  assign T478 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T482 & T479;
  assign T479 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T480 : T231;
  assign T480 = doSubMags & T481;
  assign T481 = ~ isZeroC;
  assign T482 = ~ isZeroY;
  assign isZeroY = T483 == 3'h0;
  assign T483 = T12[5'h1b:5'h19];
  assign T484 = T487 | T485;
  assign T485 = T486 & T439;
  assign T486 = doIncrSig & roundingMode_nearest_even;
  assign T487 = T489 | T488;
  assign T488 = doIncrSig & allRound;
  assign T489 = T493 | T490;
  assign T490 = T491 & anyRound;
  assign T491 = T492 & roundDirectUp;
  assign T492 = ~ doIncrSig;
  assign T493 = T494 & T4;
  assign T494 = T495 & T439;
  assign T495 = T496 & roundingMode_nearest_even;
  assign T496 = ~ doIncrSig;
  assign T497 = T502 ? T498 : 26'h0;
  assign T498 = T499 >> 2'h2;
  assign T499 = T12 & T500;
  assign T500 = {1'h0, T501};
  assign T501 = ~ roundMask;
  assign T502 = T504 & T503;
  assign T503 = ~ roundEven;
  assign T504 = ~ roundUp;
  assign T505 = T508 | T506;
  assign T506 = T507 ? sExpX3 : 11'h0;
  assign T507 = sigY3[5'h18:5'h18];
  assign T508 = T510 ? T509 : 11'h0;
  assign T509 = sExpX3 + 11'h1;
  assign T510 = sigY3[5'h19:5'h19];
  assign underflow = commonCase & underflowY;
  assign underflowY = roundInexact & T511;
  assign T511 = T516 | T512;
  assign T512 = T382 <= T513;
  assign T513 = {2'h0, T514};
  assign T514 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign sigX3Shift1 = T515 == 2'h0;
  assign T515 = T12[5'h1b:5'h1a];
  assign T516 = sExpX3[4'ha:4'ha];
  assign T517 = {invalid, 1'h0};
  assign invalid = T536 | notSigNaN_invalid;
  assign notSigNaN_invalid = T533 | T518;
  assign T518 = T519 & doSubMags;
  assign T519 = T522 & isInfC;
  assign isInfC = isSpecialC & T520;
  assign T520 = T521 ^ 1'h1;
  assign T521 = T110[3'h6:3'h6];
  assign T522 = T528 & T523;
  assign T523 = isInfA | isInfB;
  assign isInfB = isSpecialB & T524;
  assign T524 = T525 ^ 1'h1;
  assign T525 = T116[3'h6:3'h6];
  assign isInfA = isSpecialA & T526;
  assign T526 = T527 ^ 1'h1;
  assign T527 = T113[3'h6:3'h6];
  assign T528 = T531 & T529;
  assign T529 = ~ isNaNB;
  assign isNaNB = isSpecialB & T530;
  assign T530 = T116[3'h6:3'h6];
  assign T531 = ~ isNaNA;
  assign isNaNA = isSpecialA & T532;
  assign T532 = T113[3'h6:3'h6];
  assign T533 = T535 | T534;
  assign T534 = isZeroA & isInfB;
  assign T535 = isInfA & isZeroB;
  assign T536 = T540 | isSigNaNC;
  assign isSigNaNC = isNaNC & T537;
  assign T537 = T538 ^ 1'h1;
  assign T538 = T164[5'h16:5'h16];
  assign isNaNC = isSpecialC & T539;
  assign T539 = T110[3'h6:3'h6];
  assign T540 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T541;
  assign T541 = T542 ^ 1'h1;
  assign T542 = T177[5'h16:5'h16];
  assign isSigNaNA = isNaNA & T543;
  assign T543 = T544 ^ 1'h1;
  assign T544 = T179[5'h16:5'h16];
  assign io_out = T545;
  assign T545 = {signOut, T546};
  assign T546 = {expOut, fractOut};
  assign fractOut = fractY | T547;
  assign T547 = 23'h0 - T548;
  assign T548 = {22'h0, T549};
  assign T549 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T550;
  assign T550 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T553 | T551;
  assign T551 = roundingMode_max & T552;
  assign T552 = ~ signY;
  assign T553 = roundingMode_nearest_even | T554;
  assign T554 = roundingMode_min & signY;
  assign isNaNOut = T555 | notSigNaN_invalid;
  assign T555 = T556 | isNaNC;
  assign T556 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T558 : T557;
  assign T557 = sigY3[5'h17:1'h1];
  assign T558 = sigY3[5'h16:1'h0];
  assign expOut = T560 | T559;
  assign T559 = isNaNOut ? 9'h1c0 : 9'h0;
  assign T560 = T565 | T561;
  assign T561 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign notNaN_isInfOut = T563 | T562;
  assign T562 = overflow & overflowY_roundMagUp;
  assign T563 = T564 | isInfC;
  assign T564 = isInfA | isInfB;
  assign T565 = T567 | T566;
  assign T566 = isSatOut ? 9'h17f : 9'h0;
  assign T567 = T570 & T568;
  assign T568 = ~ T569;
  assign T569 = notNaN_isInfOut ? 9'h40 : 9'h0;
  assign T570 = T573 & T571;
  assign T571 = ~ T572;
  assign T572 = isSatOut ? 9'h80 : 9'h0;
  assign T573 = T580 & T574;
  assign T574 = ~ T575;
  assign T575 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign notSpecial_isZeroOut = T579 | totalUnderflowY;
  assign totalUnderflowY = T578 | T576;
  assign T576 = T577 < 9'h6b;
  assign T577 = sExpY[4'h8:1'h0];
  assign T578 = sExpY[4'h9:4'h9];
  assign T579 = notSpecial_addZeros | isZeroY;
  assign T580 = sExpY[4'h8:1'h0];
  assign signOut = T582 | T581;
  assign T581 = commonCase & signY;
  assign T582 = T586 | T583;
  assign T583 = T584 & opSignC;
  assign T584 = T585 & isSpecialC;
  assign T585 = mulSpecial ^ 1'h1;
  assign T586 = T590 | T587;
  assign T587 = T588 & signProd;
  assign T588 = mulSpecial & T589;
  assign T589 = isSpecialC ^ 1'h1;
  assign T590 = T591 | isNaNOut;
  assign T591 = T592 & opSignC;
  assign T592 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_0(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T0;
  reg [2:0] in_rm;
  wire[2:0] T1;
  wire[32:0] T2;
  reg [64:0] in_in3;
  wire[64:0] T3;
  wire[64:0] T4;
  wire[64:0] T5;
  wire[32:0] zero;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[32:0] T12;
  reg [64:0] in_in2;
  wire[64:0] T13;
  wire[64:0] T14;
  wire T15;
  wire[32:0] T16;
  reg [64:0] in_in1;
  wire[64:0] T17;
  wire[1:0] T18;
  reg [4:0] in_cmd;
  wire[4:0] T19;
  wire[4:0] T20;
  wire[4:0] T21;
  wire[1:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  reg [4:0] R27;
  wire[4:0] T28;
  wire[4:0] res_exc;
  wire[4:0] fma_io_exceptionFlags;
  reg  valid;
  reg [64:0] R29;
  wire[64:0] T30;
  wire[64:0] res_data;
  wire[64:0] T31;
  wire[32:0] fma_io_out;
  reg  R32;
  wire T33;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R27 = {1{$random}};
    valid = {1{$random}};
    R29 = {3{$random}};
    R32 = {1{$random}};
  end
`endif

  assign T0 = in_rm[1'h1:1'h0];
  assign T1 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T2 = in_in3[6'h20:1'h0];
  assign T3 = T9 ? T5 : T4;
  assign T4 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T5 = {32'h0, zero};
  assign zero = T6 << 6'h20;
  assign T6 = T8 ^ T7;
  assign T7 = io_in_bits_in2[6'h20:6'h20];
  assign T8 = io_in_bits_in1[6'h20:6'h20];
  assign T9 = io_in_valid & T10;
  assign T10 = T11 ^ 1'h1;
  assign T11 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T12 = in_in2[6'h20:1'h0];
  assign T13 = T15 ? 65'h80000000 : T14;
  assign T14 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T15 = io_in_valid & io_in_bits_swap23;
  assign T16 = in_in1[6'h20:1'h0];
  assign T17 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T18 = in_cmd[1'h1:1'h0];
  assign T19 = io_in_valid ? T21 : T20;
  assign T20 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T21 = {3'h0, T22};
  assign T22 = {T24, T23};
  assign T23 = io_in_bits_cmd[1'h0:1'h0];
  assign T24 = T26 & T25;
  assign T25 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T26 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R27;
  assign T28 = valid ? res_exc : R27;
  assign res_exc = fma_io_exceptionFlags;
  assign io_out_bits_data = R29;
  assign T30 = valid ? res_data : R29;
  assign res_data = T31;
  assign T31 = {32'h0, fma_io_out};
  assign io_out_valid = R32;
  assign T33 = reset ? 1'h0 : valid;
  mulAddSubRecodedFloatN_0 fma(
       .io_op( T18 ),
       .io_a( T16 ),
       .io_b( T12 ),
       .io_c( T2 ),
       .io_roundingMode( T0 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T9) begin
      in_in3 <= T5;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T15) begin
      in_in2 <= 65'h80000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T21;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(valid) begin
      R27 <= res_exc;
    end
    valid <= io_in_valid;
    if(valid) begin
      R29 <= res_data;
    end
    if(reset) begin
      R32 <= 1'h0;
    end else begin
      R32 <= valid;
    end
  end
endmodule

module mulAddSubRecodedFloatN_1(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire roundInexact;
  wire anyRound;
  wire T4;
  wire[56:0] T5;
  wire[56:0] T6;
  wire[54:0] T7;
  wire[55:0] roundMask;
  wire[55:0] T8;
  wire[53:0] T9;
  wire[53:0] T10;
  wire T11;
  wire[56:0] T12;
  wire[87:0] T13;
  wire T14;
  wire T15;
  wire[31:0] T16;
  wire[31:0] absSigSumExtraMask;
  wire[30:0] T17;
  wire[14:0] T18;
  wire[6:0] T19;
  wire[2:0] T20;
  wire T21;
  wire[2:0] T22;
  wire[6:0] T23;
  wire[14:0] T24;
  wire[30:0] T25;
  wire[32:0] T26;
  wire[4:0] normTo2ShiftDist;
  wire[4:0] estNormDist_5;
  wire[4:0] T27;
  wire[7:0] estNormDist;
  wire[7:0] T28;
  wire[7:0] estNormPos_dist;
  wire[7:0] T29;
  wire[7:0] T30;
  wire[7:0] T31;
  wire[7:0] T32;
  wire[7:0] T33;
  wire[7:0] T34;
  wire[7:0] T35;
  wire[7:0] T36;
  wire[7:0] T37;
  wire[7:0] T38;
  wire[7:0] T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[7:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[7:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[7:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T54;
  wire[7:0] T55;
  wire[7:0] T56;
  wire[7:0] T57;
  wire[7:0] T58;
  wire[7:0] T59;
  wire[7:0] T60;
  wire[7:0] T61;
  wire[7:0] T62;
  wire[7:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[7:0] T66;
  wire[7:0] T67;
  wire[7:0] T68;
  wire[7:0] T69;
  wire[7:0] T70;
  wire[7:0] T71;
  wire[7:0] T72;
  wire[7:0] T73;
  wire[7:0] T74;
  wire[7:0] T75;
  wire[7:0] T76;
  wire[7:0] T77;
  wire[7:0] T78;
  wire[7:0] T79;
  wire[7:0] T80;
  wire[7:0] T81;
  wire[7:0] T82;
  wire[7:0] T83;
  wire[7:0] T84;
  wire[7:0] T85;
  wire[7:0] T86;
  wire[7:0] T87;
  wire[7:0] T88;
  wire[7:0] T89;
  wire[7:0] T90;
  wire[7:0] T91;
  wire[7:0] T92;
  wire[7:0] T93;
  wire[7:0] T94;
  wire[7:0] T95;
  wire[7:0] T96;
  wire[7:0] T97;
  wire[7:0] T98;
  wire[7:0] T99;
  wire[7:0] T100;
  wire[7:0] T101;
  wire[7:0] T102;
  wire[7:0] T103;
  wire[7:0] T104;
  wire[7:0] T105;
  wire[7:0] T106;
  wire[7:0] T107;
  wire[7:0] T108;
  wire[7:0] T109;
  wire[7:0] T110;
  wire[7:0] T111;
  wire[7:0] T112;
  wire[7:0] T113;
  wire[7:0] T114;
  wire[7:0] T115;
  wire[7:0] T116;
  wire[7:0] T117;
  wire[7:0] T118;
  wire[7:0] T119;
  wire[7:0] T120;
  wire[7:0] T121;
  wire[7:0] T122;
  wire[7:0] T123;
  wire[7:0] T124;
  wire[7:0] T125;
  wire[7:0] T126;
  wire[7:0] T127;
  wire[7:0] T128;
  wire[7:0] T129;
  wire[7:0] T130;
  wire[7:0] T131;
  wire[7:0] T132;
  wire[7:0] T133;
  wire[7:0] T134;
  wire T135;
  wire[108:0] T136;
  wire[108:0] T137;
  wire[107:0] T138;
  wire[107:0] T139;
  wire[161:0] sigSum;
  wire[161:0] T140;
  wire[162:0] T141;
  wire T142;
  wire doSubMags;
  wire opSignC;
  wire T143;
  wire T144;
  wire signProd;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire[52:0] T150;
  wire[52:0] CExtraMask;
  wire[20:0] T151;
  wire[4:0] T152;
  wire T153;
  wire[4:0] T154;
  wire[20:0] T155;
  wire[52:0] T156;
  wire[256:0] T157;
  wire[7:0] T158;
  wire[13:0] T159;
  wire[13:0] T160;
  wire[13:0] sNatCAlignDist;
  wire[13:0] T161;
  wire[11:0] T162;
  wire[13:0] sExpAlignedProd;
  wire[13:0] T163;
  wire[13:0] T164;
  wire[11:0] T165;
  wire[13:0] T166;
  wire[10:0] T167;
  wire[11:0] T168;
  wire[2:0] T169;
  wire[2:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire[12:0] T174;
  wire CAlignDist_floor;
  wire T175;
  wire isZeroProd;
  wire isZeroB;
  wire[2:0] T176;
  wire isZeroA;
  wire[2:0] T177;
  wire[3:0] T178;
  wire[1:0] T179;
  wire T180;
  wire[1:0] T181;
  wire[3:0] T182;
  wire T183;
  wire[1:0] T184;
  wire T185;
  wire[1:0] T186;
  wire T187;
  wire[15:0] T188;
  wire[15:0] T189;
  wire[15:0] T190;
  wire[14:0] T191;
  wire[15:0] T192;
  wire[15:0] T193;
  wire[15:0] T194;
  wire[13:0] T195;
  wire[15:0] T196;
  wire[15:0] T197;
  wire[15:0] T198;
  wire[11:0] T199;
  wire[15:0] T200;
  wire[15:0] T201;
  wire[15:0] T202;
  wire[7:0] T203;
  wire[15:0] T204;
  wire[15:0] T205;
  wire[15:0] T206;
  wire[7:0] T207;
  wire[15:0] T208;
  wire[15:0] T209;
  wire[11:0] T210;
  wire[15:0] T211;
  wire[15:0] T212;
  wire[13:0] T213;
  wire[15:0] T214;
  wire[15:0] T215;
  wire[14:0] T216;
  wire[31:0] T217;
  wire[31:0] T218;
  wire[31:0] T219;
  wire[30:0] T220;
  wire[31:0] T221;
  wire[31:0] T222;
  wire[31:0] T223;
  wire[29:0] T224;
  wire[31:0] T225;
  wire[31:0] T226;
  wire[31:0] T227;
  wire[27:0] T228;
  wire[31:0] T229;
  wire[31:0] T230;
  wire[31:0] T231;
  wire[23:0] T232;
  wire[31:0] T233;
  wire[31:0] T234;
  wire[31:0] T235;
  wire[15:0] T236;
  wire[31:0] T237;
  wire[31:0] T238;
  wire[31:0] T239;
  wire[15:0] T240;
  wire[31:0] T241;
  wire[31:0] T242;
  wire[23:0] T243;
  wire[31:0] T244;
  wire[31:0] T245;
  wire[27:0] T246;
  wire[31:0] T247;
  wire[31:0] T248;
  wire[29:0] T249;
  wire[31:0] T250;
  wire[31:0] T251;
  wire[30:0] T252;
  wire[52:0] sigC;
  wire[51:0] T253;
  wire T254;
  wire isZeroC;
  wire[2:0] T255;
  wire[161:0] T256;
  wire[161:0] T257;
  wire[161:0] T258;
  wire[160:0] T259;
  wire[107:0] T260;
  wire[107:0] T261;
  wire[52:0] negSigC;
  wire[52:0] T262;
  wire[161:0] T263;
  wire[106:0] T264;
  wire[105:0] T265;
  wire[52:0] sigB;
  wire[51:0] T266;
  wire T267;
  wire[52:0] sigA;
  wire[51:0] T268;
  wire T269;
  wire[108:0] T270;
  wire[107:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire[7:0] CDom_estNormDist;
  wire[7:0] T379;
  wire[5:0] T380;
  wire[7:0] T381;
  wire T382;
  wire CAlignDist_0;
  wire T383;
  wire[12:0] T384;
  wire isCDominant;
  wire T385;
  wire T386;
  wire[12:0] T387;
  wire T388;
  wire[1:0] T389;
  wire T390;
  wire[1:0] T391;
  wire T392;
  wire[3:0] T393;
  wire[1:0] T394;
  wire T395;
  wire[1:0] T396;
  wire[3:0] T397;
  wire T398;
  wire[1:0] T399;
  wire T400;
  wire[1:0] T401;
  wire T402;
  wire[7:0] T403;
  wire[7:0] T404;
  wire[7:0] T405;
  wire[6:0] T406;
  wire[7:0] T407;
  wire[7:0] T408;
  wire[7:0] T409;
  wire[5:0] T410;
  wire[7:0] T411;
  wire[7:0] T412;
  wire[7:0] T413;
  wire[3:0] T414;
  wire[7:0] T415;
  wire[7:0] T416;
  wire[7:0] T417;
  wire[3:0] T418;
  wire[7:0] T419;
  wire[7:0] T420;
  wire[5:0] T421;
  wire[7:0] T422;
  wire[7:0] T423;
  wire[6:0] T424;
  wire[15:0] T425;
  wire[15:0] T426;
  wire[15:0] T427;
  wire[14:0] T428;
  wire[15:0] T429;
  wire[15:0] T430;
  wire[15:0] T431;
  wire[13:0] T432;
  wire[15:0] T433;
  wire[15:0] T434;
  wire[15:0] T435;
  wire[11:0] T436;
  wire[15:0] T437;
  wire[15:0] T438;
  wire[15:0] T439;
  wire[7:0] T440;
  wire[15:0] T441;
  wire[15:0] T442;
  wire[15:0] T443;
  wire[7:0] T444;
  wire[15:0] T445;
  wire[15:0] T446;
  wire[11:0] T447;
  wire[15:0] T448;
  wire[15:0] T449;
  wire[13:0] T450;
  wire[15:0] T451;
  wire[15:0] T452;
  wire[14:0] T453;
  wire[31:0] T454;
  wire[87:0] cFirstNormAbsSigSum;
  wire[87:0] T455;
  wire[86:0] T456;
  wire[86:0] notCDom_pos_firstNormAbsSigSum;
  wire[86:0] T457;
  wire[86:0] T458;
  wire[53:0] T459;
  wire[53:0] T460;
  wire[32:0] T461;
  wire[86:0] T462;
  wire[86:0] T463;
  wire[85:0] T464;
  wire[85:0] T465;
  wire T466;
  wire[86:0] T467;
  wire[65:0] T468;
  wire T469;
  wire T470;
  wire[1:0] firstReduceSigSum;
  wire T471;
  wire[43:0] T472;
  wire T473;
  wire[31:0] T474;
  wire T475;
  wire T476;
  wire[1:0] firstReduceNotSigSum;
  wire T477;
  wire[43:0] T478;
  wire[161:0] notSigSum;
  wire T479;
  wire[31:0] T480;
  wire[64:0] T481;
  wire T482;
  wire T483;
  wire[86:0] T484;
  wire[86:0] T485;
  wire T486;
  wire T487;
  wire[10:0] T488;
  wire T489;
  wire[10:0] T490;
  wire[85:0] T491;
  wire[86:0] T492;
  wire[21:0] T493;
  wire[21:0] T494;
  wire[64:0] T495;
  wire T496;
  wire T497;
  wire[86:0] CDom_firstNormAbsSigSum;
  wire[86:0] T498;
  wire[86:0] T499;
  wire[86:0] T500;
  wire T501;
  wire[85:0] T502;
  wire[86:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[86:0] T507;
  wire[86:0] T508;
  wire[86:0] T509;
  wire T510;
  wire[85:0] T511;
  wire[86:0] T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire[86:0] T517;
  wire[86:0] T518;
  wire[86:0] T519;
  wire T520;
  wire[85:0] T521;
  wire[86:0] T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire[86:0] T527;
  wire[86:0] T528;
  wire T529;
  wire[85:0] T530;
  wire[86:0] T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire[87:0] T537;
  wire[87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire[87:0] T538;
  wire[87:0] T539;
  wire[33:0] T540;
  wire[87:0] T541;
  wire[87:0] T542;
  wire[1:0] T543;
  wire[87:0] T544;
  wire[64:0] T545;
  wire T546;
  wire[63:0] T547;
  wire T548;
  wire T549;
  wire[87:0] T550;
  wire[87:0] T551;
  wire T552;
  wire[10:0] T553;
  wire[86:0] T554;
  wire[87:0] T555;
  wire[65:0] T556;
  wire T557;
  wire T558;
  wire[87:0] T559;
  wire T560;
  wire[31:0] T561;
  wire[31:0] T562;
  wire[31:0] T563;
  wire doIncrSig;
  wire T564;
  wire T565;
  wire T566;
  wire[86:0] T567;
  wire[86:0] T568;
  wire[53:0] T569;
  wire[21:0] T570;
  wire[5:0] T571;
  wire[1:0] T572;
  wire T573;
  wire[1:0] T574;
  wire[5:0] T575;
  wire[21:0] T576;
  wire[53:0] T577;
  wire[8192:0] T578;
  wire[12:0] T579;
  wire[12:0] T580;
  wire[13:0] sExpX3;
  wire[13:0] T581;
  wire[13:0] sExpSum;
  wire[13:0] T582;
  wire T583;
  wire[3:0] T584;
  wire[1:0] T585;
  wire T586;
  wire[1:0] T587;
  wire[3:0] T588;
  wire T589;
  wire[1:0] T590;
  wire T591;
  wire[1:0] T592;
  wire T593;
  wire[15:0] T594;
  wire[15:0] T595;
  wire[15:0] T596;
  wire[14:0] T597;
  wire[15:0] T598;
  wire[15:0] T599;
  wire[15:0] T600;
  wire[13:0] T601;
  wire[15:0] T602;
  wire[15:0] T603;
  wire[15:0] T604;
  wire[11:0] T605;
  wire[15:0] T606;
  wire[15:0] T607;
  wire[15:0] T608;
  wire[7:0] T609;
  wire[15:0] T610;
  wire[15:0] T611;
  wire[15:0] T612;
  wire[7:0] T613;
  wire[15:0] T614;
  wire[15:0] T615;
  wire[11:0] T616;
  wire[15:0] T617;
  wire[15:0] T618;
  wire[13:0] T619;
  wire[15:0] T620;
  wire[15:0] T621;
  wire[14:0] T622;
  wire[31:0] T623;
  wire[31:0] T624;
  wire[31:0] T625;
  wire[30:0] T626;
  wire[31:0] T627;
  wire[31:0] T628;
  wire[31:0] T629;
  wire[29:0] T630;
  wire[31:0] T631;
  wire[31:0] T632;
  wire[31:0] T633;
  wire[27:0] T634;
  wire[31:0] T635;
  wire[31:0] T636;
  wire[31:0] T637;
  wire[23:0] T638;
  wire[31:0] T639;
  wire[31:0] T640;
  wire[31:0] T641;
  wire[15:0] T642;
  wire[31:0] T643;
  wire[31:0] T644;
  wire[31:0] T645;
  wire[15:0] T646;
  wire[31:0] T647;
  wire[31:0] T648;
  wire[23:0] T649;
  wire[31:0] T650;
  wire[31:0] T651;
  wire[27:0] T652;
  wire[31:0] T653;
  wire[31:0] T654;
  wire[29:0] T655;
  wire[31:0] T656;
  wire[31:0] T657;
  wire[30:0] T658;
  wire[55:0] T659;
  wire[55:0] T660;
  wire T661;
  wire T662;
  wire[56:0] T663;
  wire[56:0] T664;
  wire[55:0] roundPosMask;
  wire[55:0] T665;
  wire[54:0] T666;
  wire[54:0] T667;
  wire T668;
  wire allRound;
  wire allRoundExtra;
  wire[56:0] T669;
  wire[56:0] T670;
  wire[54:0] T671;
  wire[56:0] T672;
  wire commonCase;
  wire T673;
  wire notSpecial_addZeros;
  wire T674;
  wire addSpecial;
  wire isSpecialC;
  wire[1:0] T675;
  wire mulSpecial;
  wire isSpecialB;
  wire[1:0] T676;
  wire isSpecialA;
  wire[1:0] T677;
  wire overflow;
  wire overflowY;
  wire[2:0] T678;
  wire[13:0] sExpY;
  wire[13:0] T679;
  wire[13:0] T680;
  wire T681;
  wire[1:0] T682;
  wire[54:0] sigY3;
  wire[54:0] T683;
  wire[54:0] T684;
  wire[54:0] T685;
  wire[54:0] T686;
  wire[54:0] T687;
  wire[54:0] T688;
  wire[54:0] T689;
  wire[56:0] T690;
  wire[56:0] T691;
  wire roundEven;
  wire T692;
  wire T693;
  wire T694;
  wire roundingMode_nearest_even;
  wire T695;
  wire T696;
  wire T697;
  wire[54:0] T698;
  wire[54:0] T699;
  wire roundUp;
  wire T700;
  wire T701;
  wire roundDirectUp;
  wire roundingMode_max;
  wire roundingMode_min;
  wire signY;
  wire T702;
  wire doNegSignSum;
  wire T703;
  wire T704;
  wire T705;
  wire isZeroY;
  wire[2:0] T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[54:0] T720;
  wire[54:0] T721;
  wire[56:0] T722;
  wire[56:0] T723;
  wire[55:0] T724;
  wire T725;
  wire T726;
  wire T727;
  wire[13:0] T728;
  wire[13:0] T729;
  wire T730;
  wire[13:0] T731;
  wire[13:0] T732;
  wire T733;
  wire underflow;
  wire underflowY;
  wire T734;
  wire T735;
  wire[12:0] T736;
  wire[10:0] T737;
  wire sigX3Shift1;
  wire[1:0] T738;
  wire T739;
  wire[1:0] T740;
  wire invalid;
  wire notSigNaN_invalid;
  wire T741;
  wire T742;
  wire isInfC;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire isInfB;
  wire T747;
  wire T748;
  wire isInfA;
  wire T749;
  wire T750;
  wire T751;
  wire T752;
  wire isNaNB;
  wire T753;
  wire T754;
  wire isNaNA;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire isSigNaNC;
  wire T760;
  wire T761;
  wire isNaNC;
  wire T762;
  wire T763;
  wire isSigNaNB;
  wire T764;
  wire T765;
  wire isSigNaNA;
  wire T766;
  wire T767;
  wire[64:0] T768;
  wire[63:0] T769;
  wire[51:0] fractOut;
  wire[51:0] T770;
  wire[51:0] T771;
  wire T772;
  wire isSatOut;
  wire T773;
  wire overflowY_roundMagUp;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire isNaNOut;
  wire T778;
  wire T779;
  wire[51:0] fractY;
  wire[51:0] T780;
  wire[51:0] T781;
  wire[11:0] expOut;
  wire[11:0] T782;
  wire[11:0] T783;
  wire[11:0] T784;
  wire notNaN_isInfOut;
  wire T785;
  wire T786;
  wire T787;
  wire[11:0] T788;
  wire[11:0] T789;
  wire[11:0] T790;
  wire[11:0] T791;
  wire[11:0] T792;
  wire[11:0] T793;
  wire[11:0] T794;
  wire[11:0] T795;
  wire[11:0] T796;
  wire[11:0] T797;
  wire[11:0] T798;
  wire notSpecial_isZeroOut;
  wire totalUnderflowY;
  wire T799;
  wire[11:0] T800;
  wire T801;
  wire T802;
  wire[11:0] T803;
  wire signOut;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;


  assign io_exceptionFlags = T0;
  assign T0 = {T740, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & roundInexact;
  assign roundInexact = doIncrSig ? T668 : anyRound;
  assign anyRound = T662 | T4;
  assign T4 = T5 != 57'h0;
  assign T5 = T12 & T6;
  assign T6 = {2'h0, T7};
  assign T7 = roundMask >> 1'h1;
  assign roundMask = T659 | T8;
  assign T8 = {T9, 2'h3};
  assign T9 = T569 | T10;
  assign T10 = {53'h0, T11};
  assign T11 = T12[6'h37:6'h37];
  assign T12 = T13[6'h38:1'h0];
  assign T13 = {T567, T14};
  assign T14 = doIncrSig ? T560 : T15;
  assign T15 = T16 != 32'h0;
  assign T16 = T454 & absSigSumExtraMask;
  assign absSigSumExtraMask = {T17, 1'h1};
  assign T17 = {T425, T18};
  assign T18 = {T403, T19};
  assign T19 = {T393, T20};
  assign T20 = {T389, T21};
  assign T21 = T22[2'h2:2'h2];
  assign T22 = T23[3'h6:3'h4];
  assign T23 = T24[4'he:4'h8];
  assign T24 = T25[5'h1e:5'h10];
  assign T25 = T26[5'h1f:1'h1];
  assign T26 = $signed(33'h100000000) >>> normTo2ShiftDist;
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign estNormDist_5 = T27;
  assign T27 = estNormDist[3'h4:1'h0];
  assign estNormDist = isCDominant ? CDom_estNormDist : T28;
  assign T28 = T378 ? estNormPos_dist : estNormPos_dist;
  assign estNormPos_dist = T377 ? 8'h35 : T29;
  assign T29 = T376 ? 8'h36 : T30;
  assign T30 = T375 ? 8'h37 : T31;
  assign T31 = T374 ? 8'h38 : T32;
  assign T32 = T373 ? 8'h39 : T33;
  assign T33 = T372 ? 8'h3a : T34;
  assign T34 = T371 ? 8'h3b : T35;
  assign T35 = T370 ? 8'h3c : T36;
  assign T36 = T369 ? 8'h3d : T37;
  assign T37 = T368 ? 8'h3e : T38;
  assign T38 = T367 ? 8'h3f : T39;
  assign T39 = T366 ? 8'h40 : T40;
  assign T40 = T365 ? 8'h41 : T41;
  assign T41 = T364 ? 8'h42 : T42;
  assign T42 = T363 ? 8'h43 : T43;
  assign T43 = T362 ? 8'h44 : T44;
  assign T44 = T361 ? 8'h45 : T45;
  assign T45 = T360 ? 8'h46 : T46;
  assign T46 = T359 ? 8'h47 : T47;
  assign T47 = T358 ? 8'h48 : T48;
  assign T48 = T357 ? 8'h49 : T49;
  assign T49 = T356 ? 8'h4a : T50;
  assign T50 = T355 ? 8'h4b : T51;
  assign T51 = T354 ? 8'h4c : T52;
  assign T52 = T353 ? 8'h4d : T53;
  assign T53 = T352 ? 8'h4e : T54;
  assign T54 = T351 ? 8'h4f : T55;
  assign T55 = T350 ? 8'h50 : T56;
  assign T56 = T349 ? 8'h51 : T57;
  assign T57 = T348 ? 8'h52 : T58;
  assign T58 = T347 ? 8'h53 : T59;
  assign T59 = T346 ? 8'h54 : T60;
  assign T60 = T345 ? 8'h55 : T61;
  assign T61 = T344 ? 8'h56 : T62;
  assign T62 = T343 ? 8'h57 : T63;
  assign T63 = T342 ? 8'h58 : T64;
  assign T64 = T341 ? 8'h59 : T65;
  assign T65 = T340 ? 8'h5a : T66;
  assign T66 = T339 ? 8'h5b : T67;
  assign T67 = T338 ? 8'h5c : T68;
  assign T68 = T337 ? 8'h5d : T69;
  assign T69 = T336 ? 8'h5e : T70;
  assign T70 = T335 ? 8'h5f : T71;
  assign T71 = T334 ? 8'h60 : T72;
  assign T72 = T333 ? 8'h61 : T73;
  assign T73 = T332 ? 8'h62 : T74;
  assign T74 = T331 ? 8'h63 : T75;
  assign T75 = T330 ? 8'h64 : T76;
  assign T76 = T329 ? 8'h65 : T77;
  assign T77 = T328 ? 8'h66 : T78;
  assign T78 = T327 ? 8'h67 : T79;
  assign T79 = T326 ? 8'h68 : T80;
  assign T80 = T325 ? 8'h69 : T81;
  assign T81 = T324 ? 8'h6a : T82;
  assign T82 = T323 ? 8'h6b : T83;
  assign T83 = T322 ? 8'h6c : T84;
  assign T84 = T321 ? 8'h6d : T85;
  assign T85 = T320 ? 8'h6e : T86;
  assign T86 = T319 ? 8'h6f : T87;
  assign T87 = T318 ? 8'h70 : T88;
  assign T88 = T317 ? 8'h71 : T89;
  assign T89 = T316 ? 8'h72 : T90;
  assign T90 = T315 ? 8'h73 : T91;
  assign T91 = T314 ? 8'h74 : T92;
  assign T92 = T313 ? 8'h75 : T93;
  assign T93 = T312 ? 8'h76 : T94;
  assign T94 = T311 ? 8'h77 : T95;
  assign T95 = T310 ? 8'h78 : T96;
  assign T96 = T309 ? 8'h79 : T97;
  assign T97 = T308 ? 8'h7a : T98;
  assign T98 = T307 ? 8'h7b : T99;
  assign T99 = T306 ? 8'h7c : T100;
  assign T100 = T305 ? 8'h7d : T101;
  assign T101 = T304 ? 8'h7e : T102;
  assign T102 = T303 ? 8'h7f : T103;
  assign T103 = T302 ? 8'h80 : T104;
  assign T104 = T301 ? 8'h81 : T105;
  assign T105 = T300 ? 8'h82 : T106;
  assign T106 = T299 ? 8'h83 : T107;
  assign T107 = T298 ? 8'h84 : T108;
  assign T108 = T297 ? 8'h85 : T109;
  assign T109 = T296 ? 8'h86 : T110;
  assign T110 = T295 ? 8'h87 : T111;
  assign T111 = T294 ? 8'h88 : T112;
  assign T112 = T293 ? 8'h89 : T113;
  assign T113 = T292 ? 8'h8a : T114;
  assign T114 = T291 ? 8'h8b : T115;
  assign T115 = T290 ? 8'h8c : T116;
  assign T116 = T289 ? 8'h8d : T117;
  assign T117 = T288 ? 8'h8e : T118;
  assign T118 = T287 ? 8'h8f : T119;
  assign T119 = T286 ? 8'h90 : T120;
  assign T120 = T285 ? 8'h91 : T121;
  assign T121 = T284 ? 8'h92 : T122;
  assign T122 = T283 ? 8'h93 : T123;
  assign T123 = T282 ? 8'h94 : T124;
  assign T124 = T281 ? 8'h95 : T125;
  assign T125 = T280 ? 8'h96 : T126;
  assign T126 = T279 ? 8'h97 : T127;
  assign T127 = T278 ? 8'h98 : T128;
  assign T128 = T277 ? 8'h99 : T129;
  assign T129 = T276 ? 8'h9a : T130;
  assign T130 = T275 ? 8'h9b : T131;
  assign T131 = T274 ? 8'h9c : T132;
  assign T132 = T273 ? 8'h9d : T133;
  assign T133 = T272 ? 8'h9e : T134;
  assign T134 = T135 ? 8'h9f : 8'ha0;
  assign T135 = T136[1'h1:1'h1];
  assign T136 = T270 ^ T137;
  assign T137 = T138 << 1'h1;
  assign T138 = 108'h0 | T139;
  assign T139 = sigSum[7'h6c:1'h1];
  assign sigSum = T263 + T140;
  assign T140 = T141[8'ha1:1'h0];
  assign T141 = {T256, T142};
  assign T142 = T149 ^ doSubMags;
  assign doSubMags = signProd ^ opSignC;
  assign opSignC = T144 ^ T143;
  assign T143 = io_op[1'h0:1'h0];
  assign T144 = io_c[7'h40:7'h40];
  assign signProd = T146 ^ T145;
  assign T145 = io_op[1'h1:1'h1];
  assign T146 = T148 ^ T147;
  assign T147 = io_b[7'h40:7'h40];
  assign T148 = io_a[7'h40:7'h40];
  assign T149 = T150 != 53'h0;
  assign T150 = sigC & CExtraMask;
  assign CExtraMask = {T217, T151};
  assign T151 = {T188, T152};
  assign T152 = {T178, T153};
  assign T153 = T154[3'h4:3'h4];
  assign T154 = T155[5'h14:5'h10];
  assign T155 = T156[6'h34:6'h20];
  assign T156 = T157[8'h93:7'h5f];
  assign T157 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000) >>> T158;
  assign T158 = T159[3'h7:1'h0];
  assign T159 = CAlignDist_floor ? 14'h0 : T160;
  assign T160 = T173 ? sNatCAlignDist : 14'ha1;
  assign sNatCAlignDist = sExpAlignedProd - T161;
  assign T161 = {2'h0, T162};
  assign T162 = io_c[6'h3f:6'h34];
  assign sExpAlignedProd = T163 + 14'h38;
  assign T163 = T166 + T164;
  assign T164 = {2'h0, T165};
  assign T165 = io_a[6'h3f:6'h34];
  assign T166 = {T169, T167};
  assign T167 = T168[4'ha:1'h0];
  assign T168 = io_b[6'h3f:6'h34];
  assign T169 = 3'h0 - T170;
  assign T170 = {2'h0, T171};
  assign T171 = T172 ^ 1'h1;
  assign T172 = T168[4'hb:4'hb];
  assign T173 = T174 < 13'ha1;
  assign T174 = sNatCAlignDist[4'hc:1'h0];
  assign CAlignDist_floor = isZeroProd | T175;
  assign T175 = sNatCAlignDist[4'hd:4'hd];
  assign isZeroProd = isZeroA | isZeroB;
  assign isZeroB = T176 == 3'h0;
  assign T176 = T168[4'hb:4'h9];
  assign isZeroA = T177 == 3'h0;
  assign T177 = T165[4'hb:4'h9];
  assign T178 = {T184, T179};
  assign T179 = {T183, T180};
  assign T180 = T181[1'h1:1'h1];
  assign T181 = T182[2'h3:2'h2];
  assign T182 = T154[2'h3:1'h0];
  assign T183 = T181[1'h0:1'h0];
  assign T184 = {T187, T185};
  assign T185 = T186[1'h1:1'h1];
  assign T186 = T182[1'h1:1'h0];
  assign T187 = T186[1'h0:1'h0];
  assign T188 = T214 | T189;
  assign T189 = T190 & 16'haaaa;
  assign T190 = T191 << 1'h1;
  assign T191 = T192[4'he:1'h0];
  assign T192 = T211 | T193;
  assign T193 = T194 & 16'hcccc;
  assign T194 = T195 << 2'h2;
  assign T195 = T196[4'hd:1'h0];
  assign T196 = T208 | T197;
  assign T197 = T198 & 16'hf0f0;
  assign T198 = T199 << 3'h4;
  assign T199 = T200[4'hb:1'h0];
  assign T200 = T205 | T201;
  assign T201 = T202 & 16'hff00;
  assign T202 = T203 << 4'h8;
  assign T203 = T204[3'h7:1'h0];
  assign T204 = T155[4'hf:1'h0];
  assign T205 = T206 & 16'hff;
  assign T206 = {8'h0, T207};
  assign T207 = T204 >> 4'h8;
  assign T208 = T209 & 16'hf0f;
  assign T209 = {4'h0, T210};
  assign T210 = T200 >> 3'h4;
  assign T211 = T212 & 16'h3333;
  assign T212 = {2'h0, T213};
  assign T213 = T196 >> 2'h2;
  assign T214 = T215 & 16'h5555;
  assign T215 = {1'h0, T216};
  assign T216 = T192 >> 1'h1;
  assign T217 = T250 | T218;
  assign T218 = T219 & 32'haaaaaaaa;
  assign T219 = T220 << 1'h1;
  assign T220 = T221[5'h1e:1'h0];
  assign T221 = T247 | T222;
  assign T222 = T223 & 32'hcccccccc;
  assign T223 = T224 << 2'h2;
  assign T224 = T225[5'h1d:1'h0];
  assign T225 = T244 | T226;
  assign T226 = T227 & 32'hf0f0f0f0;
  assign T227 = T228 << 3'h4;
  assign T228 = T229[5'h1b:1'h0];
  assign T229 = T241 | T230;
  assign T230 = T231 & 32'hff00ff00;
  assign T231 = T232 << 4'h8;
  assign T232 = T233[5'h17:1'h0];
  assign T233 = T238 | T234;
  assign T234 = T235 & 32'hffff0000;
  assign T235 = T236 << 5'h10;
  assign T236 = T237[4'hf:1'h0];
  assign T237 = T156[5'h1f:1'h0];
  assign T238 = T239 & 32'hffff;
  assign T239 = {16'h0, T240};
  assign T240 = T237 >> 5'h10;
  assign T241 = T242 & 32'hff00ff;
  assign T242 = {8'h0, T243};
  assign T243 = T233 >> 4'h8;
  assign T244 = T245 & 32'hf0f0f0f;
  assign T245 = {4'h0, T246};
  assign T246 = T229 >> 3'h4;
  assign T247 = T248 & 32'h33333333;
  assign T248 = {2'h0, T249};
  assign T249 = T225 >> 2'h2;
  assign T250 = T251 & 32'h55555555;
  assign T251 = {1'h0, T252};
  assign T252 = T221 >> 1'h1;
  assign sigC = {T254, T253};
  assign T253 = io_c[6'h33:1'h0];
  assign T254 = isZeroC ^ 1'h1;
  assign isZeroC = T255 == 3'h0;
  assign T255 = T162[4'hb:4'h9];
  assign T256 = $signed(T257) >>> T158;
  assign T257 = T258;
  assign T258 = {doSubMags, T259};
  assign T259 = {negSigC, T260};
  assign T260 = 108'h0 - T261;
  assign T261 = {107'h0, doSubMags};
  assign negSigC = doSubMags ? T262 : sigC;
  assign T262 = ~ sigC;
  assign T263 = {55'h0, T264};
  assign T264 = T265 << 1'h1;
  assign T265 = sigA * sigB;
  assign sigB = {T267, T266};
  assign T266 = io_b[6'h33:1'h0];
  assign T267 = isZeroB ^ 1'h1;
  assign sigA = {T269, T268};
  assign T268 = io_a[6'h33:1'h0];
  assign T269 = isZeroA ^ 1'h1;
  assign T270 = {1'h0, T271};
  assign T271 = 108'h0 ^ T139;
  assign T272 = T136[2'h2:2'h2];
  assign T273 = T136[2'h3:2'h3];
  assign T274 = T136[3'h4:3'h4];
  assign T275 = T136[3'h5:3'h5];
  assign T276 = T136[3'h6:3'h6];
  assign T277 = T136[3'h7:3'h7];
  assign T278 = T136[4'h8:4'h8];
  assign T279 = T136[4'h9:4'h9];
  assign T280 = T136[4'ha:4'ha];
  assign T281 = T136[4'hb:4'hb];
  assign T282 = T136[4'hc:4'hc];
  assign T283 = T136[4'hd:4'hd];
  assign T284 = T136[4'he:4'he];
  assign T285 = T136[4'hf:4'hf];
  assign T286 = T136[5'h10:5'h10];
  assign T287 = T136[5'h11:5'h11];
  assign T288 = T136[5'h12:5'h12];
  assign T289 = T136[5'h13:5'h13];
  assign T290 = T136[5'h14:5'h14];
  assign T291 = T136[5'h15:5'h15];
  assign T292 = T136[5'h16:5'h16];
  assign T293 = T136[5'h17:5'h17];
  assign T294 = T136[5'h18:5'h18];
  assign T295 = T136[5'h19:5'h19];
  assign T296 = T136[5'h1a:5'h1a];
  assign T297 = T136[5'h1b:5'h1b];
  assign T298 = T136[5'h1c:5'h1c];
  assign T299 = T136[5'h1d:5'h1d];
  assign T300 = T136[5'h1e:5'h1e];
  assign T301 = T136[5'h1f:5'h1f];
  assign T302 = T136[6'h20:6'h20];
  assign T303 = T136[6'h21:6'h21];
  assign T304 = T136[6'h22:6'h22];
  assign T305 = T136[6'h23:6'h23];
  assign T306 = T136[6'h24:6'h24];
  assign T307 = T136[6'h25:6'h25];
  assign T308 = T136[6'h26:6'h26];
  assign T309 = T136[6'h27:6'h27];
  assign T310 = T136[6'h28:6'h28];
  assign T311 = T136[6'h29:6'h29];
  assign T312 = T136[6'h2a:6'h2a];
  assign T313 = T136[6'h2b:6'h2b];
  assign T314 = T136[6'h2c:6'h2c];
  assign T315 = T136[6'h2d:6'h2d];
  assign T316 = T136[6'h2e:6'h2e];
  assign T317 = T136[6'h2f:6'h2f];
  assign T318 = T136[6'h30:6'h30];
  assign T319 = T136[6'h31:6'h31];
  assign T320 = T136[6'h32:6'h32];
  assign T321 = T136[6'h33:6'h33];
  assign T322 = T136[6'h34:6'h34];
  assign T323 = T136[6'h35:6'h35];
  assign T324 = T136[6'h36:6'h36];
  assign T325 = T136[6'h37:6'h37];
  assign T326 = T136[6'h38:6'h38];
  assign T327 = T136[6'h39:6'h39];
  assign T328 = T136[6'h3a:6'h3a];
  assign T329 = T136[6'h3b:6'h3b];
  assign T330 = T136[6'h3c:6'h3c];
  assign T331 = T136[6'h3d:6'h3d];
  assign T332 = T136[6'h3e:6'h3e];
  assign T333 = T136[6'h3f:6'h3f];
  assign T334 = T136[7'h40:7'h40];
  assign T335 = T136[7'h41:7'h41];
  assign T336 = T136[7'h42:7'h42];
  assign T337 = T136[7'h43:7'h43];
  assign T338 = T136[7'h44:7'h44];
  assign T339 = T136[7'h45:7'h45];
  assign T340 = T136[7'h46:7'h46];
  assign T341 = T136[7'h47:7'h47];
  assign T342 = T136[7'h48:7'h48];
  assign T343 = T136[7'h49:7'h49];
  assign T344 = T136[7'h4a:7'h4a];
  assign T345 = T136[7'h4b:7'h4b];
  assign T346 = T136[7'h4c:7'h4c];
  assign T347 = T136[7'h4d:7'h4d];
  assign T348 = T136[7'h4e:7'h4e];
  assign T349 = T136[7'h4f:7'h4f];
  assign T350 = T136[7'h50:7'h50];
  assign T351 = T136[7'h51:7'h51];
  assign T352 = T136[7'h52:7'h52];
  assign T353 = T136[7'h53:7'h53];
  assign T354 = T136[7'h54:7'h54];
  assign T355 = T136[7'h55:7'h55];
  assign T356 = T136[7'h56:7'h56];
  assign T357 = T136[7'h57:7'h57];
  assign T358 = T136[7'h58:7'h58];
  assign T359 = T136[7'h59:7'h59];
  assign T360 = T136[7'h5a:7'h5a];
  assign T361 = T136[7'h5b:7'h5b];
  assign T362 = T136[7'h5c:7'h5c];
  assign T363 = T136[7'h5d:7'h5d];
  assign T364 = T136[7'h5e:7'h5e];
  assign T365 = T136[7'h5f:7'h5f];
  assign T366 = T136[7'h60:7'h60];
  assign T367 = T136[7'h61:7'h61];
  assign T368 = T136[7'h62:7'h62];
  assign T369 = T136[7'h63:7'h63];
  assign T370 = T136[7'h64:7'h64];
  assign T371 = T136[7'h65:7'h65];
  assign T372 = T136[7'h66:7'h66];
  assign T373 = T136[7'h67:7'h67];
  assign T374 = T136[7'h68:7'h68];
  assign T375 = T136[7'h69:7'h69];
  assign T376 = T136[7'h6a:7'h6a];
  assign T377 = T136[7'h6b:7'h6b];
  assign T378 = sigSum[7'h6d:7'h6d];
  assign CDom_estNormDist = T382 ? T158 : T379;
  assign T379 = {2'h0, T380};
  assign T380 = T381[3'h5:1'h0];
  assign T381 = T158 - 8'h1;
  assign T382 = CAlignDist_0 | doSubMags;
  assign CAlignDist_0 = CAlignDist_floor | T383;
  assign T383 = T384 == 13'h0;
  assign T384 = sNatCAlignDist[4'hc:1'h0];
  assign isCDominant = T388 & T385;
  assign T385 = CAlignDist_floor | T386;
  assign T386 = T387 < 13'h36;
  assign T387 = sNatCAlignDist[4'hc:1'h0];
  assign T388 = isZeroC ^ 1'h1;
  assign T389 = {T392, T390};
  assign T390 = T391[1'h1:1'h1];
  assign T391 = T22[1'h1:1'h0];
  assign T392 = T391[1'h0:1'h0];
  assign T393 = {T399, T394};
  assign T394 = {T398, T395};
  assign T395 = T396[1'h1:1'h1];
  assign T396 = T397[2'h3:2'h2];
  assign T397 = T23[2'h3:1'h0];
  assign T398 = T396[1'h0:1'h0];
  assign T399 = {T402, T400};
  assign T400 = T401[1'h1:1'h1];
  assign T401 = T397[1'h1:1'h0];
  assign T402 = T401[1'h0:1'h0];
  assign T403 = T422 | T404;
  assign T404 = T405 & 8'haa;
  assign T405 = T406 << 1'h1;
  assign T406 = T407[3'h6:1'h0];
  assign T407 = T419 | T408;
  assign T408 = T409 & 8'hcc;
  assign T409 = T410 << 2'h2;
  assign T410 = T411[3'h5:1'h0];
  assign T411 = T416 | T412;
  assign T412 = T413 & 8'hf0;
  assign T413 = T414 << 3'h4;
  assign T414 = T415[2'h3:1'h0];
  assign T415 = T24[3'h7:1'h0];
  assign T416 = T417 & 8'hf;
  assign T417 = {4'h0, T418};
  assign T418 = T415 >> 3'h4;
  assign T419 = T420 & 8'h33;
  assign T420 = {2'h0, T421};
  assign T421 = T411 >> 2'h2;
  assign T422 = T423 & 8'h55;
  assign T423 = {1'h0, T424};
  assign T424 = T407 >> 1'h1;
  assign T425 = T451 | T426;
  assign T426 = T427 & 16'haaaa;
  assign T427 = T428 << 1'h1;
  assign T428 = T429[4'he:1'h0];
  assign T429 = T448 | T430;
  assign T430 = T431 & 16'hcccc;
  assign T431 = T432 << 2'h2;
  assign T432 = T433[4'hd:1'h0];
  assign T433 = T445 | T434;
  assign T434 = T435 & 16'hf0f0;
  assign T435 = T436 << 3'h4;
  assign T436 = T437[4'hb:1'h0];
  assign T437 = T442 | T438;
  assign T438 = T439 & 16'hff00;
  assign T439 = T440 << 4'h8;
  assign T440 = T441[3'h7:1'h0];
  assign T441 = T25[4'hf:1'h0];
  assign T442 = T443 & 16'hff;
  assign T443 = {8'h0, T444};
  assign T444 = T441 >> 4'h8;
  assign T445 = T446 & 16'hf0f;
  assign T446 = {4'h0, T447};
  assign T447 = T437 >> 3'h4;
  assign T448 = T449 & 16'h3333;
  assign T449 = {2'h0, T450};
  assign T450 = T433 >> 2'h2;
  assign T451 = T452 & 16'h5555;
  assign T452 = {1'h0, T453};
  assign T453 = T429 >> 1'h1;
  assign T454 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign cFirstNormAbsSigSum = T378 ? T537 : T455;
  assign T455 = {1'h0, T456};
  assign T456 = isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign notCDom_pos_firstNormAbsSigSum = T497 ? T484 : T457;
  assign T457 = T483 ? T462 : T458;
  assign T458 = {T461, T459};
  assign T459 = 54'h0 - T460;
  assign T460 = {53'h0, doSubMags};
  assign T461 = sigSum[6'h21:1'h1];
  assign T462 = T482 ? T467 : T463;
  assign T463 = {T466, T464};
  assign T464 = 86'h0 - T465;
  assign T465 = {85'h0, doSubMags};
  assign T466 = sigSum[1'h1:1'h1];
  assign T467 = {21'h0, T468};
  assign T468 = {T481, T469};
  assign T469 = doSubMags ? T475 : T470;
  assign T470 = firstReduceSigSum[1'h0:1'h0];
  assign firstReduceSigSum = {T473, T471};
  assign T471 = T472 != 44'h0;
  assign T472 = sigSum[6'h2b:1'h0];
  assign T473 = T474 != 32'h0;
  assign T474 = sigSum[7'h4b:6'h2c];
  assign T475 = ~ T476;
  assign T476 = firstReduceNotSigSum[1'h0:1'h0];
  assign firstReduceNotSigSum = {T479, T477};
  assign T477 = T478 != 44'h0;
  assign T478 = notSigSum[6'h2b:1'h0];
  assign notSigSum = ~ sigSum;
  assign T479 = T480 != 32'h0;
  assign T480 = notSigSum[7'h4b:6'h2c];
  assign T481 = sigSum[7'h6c:6'h2c];
  assign T482 = estNormPos_dist[3'h4:3'h4];
  assign T483 = estNormPos_dist[3'h5:3'h5];
  assign T484 = T496 ? T492 : T485;
  assign T485 = {T491, T486};
  assign T486 = doSubMags ? T489 : T487;
  assign T487 = T488 != 11'h0;
  assign T488 = sigSum[4'hb:1'h1];
  assign T489 = T490 == 11'h0;
  assign T490 = notSigSum[4'hb:1'h1];
  assign T491 = sigSum[7'h61:4'hc];
  assign T492 = {T495, T493};
  assign T493 = 22'h0 - T494;
  assign T494 = {21'h0, doSubMags};
  assign T495 = sigSum[7'h41:1'h1];
  assign T496 = estNormPos_dist[3'h5:3'h5];
  assign T497 = estNormPos_dist[3'h6:3'h6];
  assign CDom_firstNormAbsSigSum = T498;
  assign T498 = T507 | T499;
  assign T499 = T503 & T500;
  assign T500 = {T502, T501};
  assign T501 = firstReduceNotSigSum[1'h0:1'h0];
  assign T502 = notSigSum[8'h81:6'h2c];
  assign T503 = T504 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T504 = T505;
  assign T505 = doSubMags & T506;
  assign T506 = CDom_estNormDist[3'h5:3'h5];
  assign T507 = T517 | T508;
  assign T508 = T512 & T509;
  assign T509 = {T511, T510};
  assign T510 = firstReduceNotSigSum != 2'h0;
  assign T511 = notSigSum[8'ha1:7'h4c];
  assign T512 = T513 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T513 = T514;
  assign T514 = doSubMags & T515;
  assign T515 = ~ T516;
  assign T516 = CDom_estNormDist[3'h5:3'h5];
  assign T517 = T527 | T518;
  assign T518 = T522 & T519;
  assign T519 = {T521, T520};
  assign T520 = firstReduceSigSum[1'h0:1'h0];
  assign T521 = sigSum[8'h81:6'h2c];
  assign T522 = T523 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T523 = T524;
  assign T524 = T526 & T525;
  assign T525 = CDom_estNormDist[3'h5:3'h5];
  assign T526 = ~ doSubMags;
  assign T527 = T531 & T528;
  assign T528 = {T530, T529};
  assign T529 = firstReduceSigSum != 2'h0;
  assign T530 = sigSum[8'ha1:7'h4c];
  assign T531 = T532 ? 87'h7fffffffffffffffffffff : 87'h0;
  assign T532 = T533;
  assign T533 = T536 & T534;
  assign T534 = ~ T535;
  assign T535 = CDom_estNormDist[3'h5:3'h5];
  assign T536 = ~ doSubMags;
  assign T537 = isCDominant ? T559 : notCDom_neg_cFirstNormAbsSigSum;
  assign notCDom_neg_cFirstNormAbsSigSum = T558 ? T550 : T538;
  assign T538 = T549 ? T541 : T539;
  assign T539 = T540 << 6'h36;
  assign T540 = notSigSum[6'h22:1'h1];
  assign T541 = T548 ? T544 : T542;
  assign T542 = T543 << 7'h56;
  assign T543 = notSigSum[2'h2:1'h1];
  assign T544 = {23'h0, T545};
  assign T545 = {T547, T546};
  assign T546 = firstReduceNotSigSum[1'h0:1'h0];
  assign T547 = notSigSum[7'h6b:6'h2c];
  assign T548 = estNormPos_dist[3'h4:3'h4];
  assign T549 = estNormPos_dist[3'h5:3'h5];
  assign T550 = T557 ? T555 : T551;
  assign T551 = {T554, T552};
  assign T552 = T553 != 11'h0;
  assign T553 = notSigSum[4'hb:1'h1];
  assign T554 = notSigSum[7'h62:4'hc];
  assign T555 = T556 << 5'h16;
  assign T556 = notSigSum[7'h42:1'h1];
  assign T557 = estNormPos_dist[3'h5:3'h5];
  assign T558 = estNormPos_dist[3'h6:3'h6];
  assign T559 = {1'h0, CDom_firstNormAbsSigSum};
  assign T560 = T561 == 32'h0;
  assign T561 = T562 & absSigSumExtraMask;
  assign T562 = ~ T563;
  assign T563 = cFirstNormAbsSigSum[5'h1f:1'h0];
  assign doIncrSig = T564 & doSubMags;
  assign T564 = T566 & T565;
  assign T565 = ~ T378;
  assign T566 = ~ isCDominant;
  assign T567 = T568 >> normTo2ShiftDist;
  assign T568 = cFirstNormAbsSigSum[7'h57:1'h1];
  assign T569 = {T623, T570};
  assign T570 = {T594, T571};
  assign T571 = {T584, T572};
  assign T572 = {T583, T573};
  assign T573 = T574[1'h1:1'h1];
  assign T574 = T575[3'h5:3'h4];
  assign T575 = T576[5'h15:5'h10];
  assign T576 = T577[6'h35:6'h20];
  assign T577 = T578[11'h403:10'h3ce];
  assign T578 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000) >>> T579;
  assign T579 = ~ T580;
  assign T580 = sExpX3[4'hc:1'h0];
  assign sExpX3 = sExpSum - T581;
  assign T581 = {6'h0, estNormDist};
  assign sExpSum = CAlignDist_floor ? T582 : sExpAlignedProd;
  assign T582 = {2'h0, T162};
  assign T583 = T574[1'h0:1'h0];
  assign T584 = {T590, T585};
  assign T585 = {T589, T586};
  assign T586 = T587[1'h1:1'h1];
  assign T587 = T588[2'h3:2'h2];
  assign T588 = T575[2'h3:1'h0];
  assign T589 = T587[1'h0:1'h0];
  assign T590 = {T593, T591};
  assign T591 = T592[1'h1:1'h1];
  assign T592 = T588[1'h1:1'h0];
  assign T593 = T592[1'h0:1'h0];
  assign T594 = T620 | T595;
  assign T595 = T596 & 16'haaaa;
  assign T596 = T597 << 1'h1;
  assign T597 = T598[4'he:1'h0];
  assign T598 = T617 | T599;
  assign T599 = T600 & 16'hcccc;
  assign T600 = T601 << 2'h2;
  assign T601 = T602[4'hd:1'h0];
  assign T602 = T614 | T603;
  assign T603 = T604 & 16'hf0f0;
  assign T604 = T605 << 3'h4;
  assign T605 = T606[4'hb:1'h0];
  assign T606 = T611 | T607;
  assign T607 = T608 & 16'hff00;
  assign T608 = T609 << 4'h8;
  assign T609 = T610[3'h7:1'h0];
  assign T610 = T576[4'hf:1'h0];
  assign T611 = T612 & 16'hff;
  assign T612 = {8'h0, T613};
  assign T613 = T610 >> 4'h8;
  assign T614 = T615 & 16'hf0f;
  assign T615 = {4'h0, T616};
  assign T616 = T606 >> 3'h4;
  assign T617 = T618 & 16'h3333;
  assign T618 = {2'h0, T619};
  assign T619 = T602 >> 2'h2;
  assign T620 = T621 & 16'h5555;
  assign T621 = {1'h0, T622};
  assign T622 = T598 >> 1'h1;
  assign T623 = T656 | T624;
  assign T624 = T625 & 32'haaaaaaaa;
  assign T625 = T626 << 1'h1;
  assign T626 = T627[5'h1e:1'h0];
  assign T627 = T653 | T628;
  assign T628 = T629 & 32'hcccccccc;
  assign T629 = T630 << 2'h2;
  assign T630 = T631[5'h1d:1'h0];
  assign T631 = T650 | T632;
  assign T632 = T633 & 32'hf0f0f0f0;
  assign T633 = T634 << 3'h4;
  assign T634 = T635[5'h1b:1'h0];
  assign T635 = T647 | T636;
  assign T636 = T637 & 32'hff00ff00;
  assign T637 = T638 << 4'h8;
  assign T638 = T639[5'h17:1'h0];
  assign T639 = T644 | T640;
  assign T640 = T641 & 32'hffff0000;
  assign T641 = T642 << 5'h10;
  assign T642 = T643[4'hf:1'h0];
  assign T643 = T577[5'h1f:1'h0];
  assign T644 = T645 & 32'hffff;
  assign T645 = {16'h0, T646};
  assign T646 = T643 >> 5'h10;
  assign T647 = T648 & 32'hff00ff;
  assign T648 = {8'h0, T649};
  assign T649 = T639 >> 4'h8;
  assign T650 = T651 & 32'hf0f0f0f;
  assign T651 = {4'h0, T652};
  assign T652 = T635 >> 3'h4;
  assign T653 = T654 & 32'h33333333;
  assign T654 = {2'h0, T655};
  assign T655 = T631 >> 2'h2;
  assign T656 = T657 & 32'h55555555;
  assign T657 = {1'h0, T658};
  assign T658 = T627 >> 1'h1;
  assign T659 = 56'h0 - T660;
  assign T660 = {55'h0, T661};
  assign T661 = sExpX3[4'hd:4'hd];
  assign T662 = T663 != 57'h0;
  assign T663 = T12 & T664;
  assign T664 = {1'h0, roundPosMask};
  assign roundPosMask = T665 & roundMask;
  assign T665 = {1'h0, T666};
  assign T666 = ~ T667;
  assign T667 = roundMask >> 1'h1;
  assign T668 = ~ allRound;
  assign allRound = T662 & allRoundExtra;
  assign allRoundExtra = T669 == 57'h0;
  assign T669 = T672 & T670;
  assign T670 = {2'h0, T671};
  assign T671 = roundMask >> 1'h1;
  assign T672 = ~ T12;
  assign commonCase = T674 & T673;
  assign T673 = ~ notSpecial_addZeros;
  assign notSpecial_addZeros = isZeroProd & isZeroC;
  assign T674 = ~ addSpecial;
  assign addSpecial = mulSpecial | isSpecialC;
  assign isSpecialC = T675 == 2'h3;
  assign T675 = T162[4'hb:4'ha];
  assign mulSpecial = isSpecialA | isSpecialB;
  assign isSpecialB = T676 == 2'h3;
  assign T676 = T168[4'hb:4'ha];
  assign isSpecialA = T677 == 2'h3;
  assign T677 = T165[4'hb:4'ha];
  assign overflow = commonCase & overflowY;
  assign overflowY = T678 == 3'h3;
  assign T678 = sExpY[4'hc:4'ha];
  assign sExpY = T728 | T679;
  assign T679 = T681 ? T680 : 14'h0;
  assign T680 = sExpX3 - 14'h1;
  assign T681 = T682 == 2'h0;
  assign T682 = sigY3[6'h36:6'h35];
  assign sigY3 = T698 | T683;
  assign T683 = roundEven ? T684 : 55'h0;
  assign T684 = T687 & T685;
  assign T685 = ~ T686;
  assign T686 = roundMask >> 1'h1;
  assign T687 = T688[6'h36:1'h0];
  assign T688 = T689 + 55'h1;
  assign T689 = T690 >> 2'h2;
  assign T690 = T12 | T691;
  assign T691 = {1'h0, roundMask};
  assign roundEven = doIncrSig ? T695 : T692;
  assign T692 = T694 & T693;
  assign T693 = ~ T4;
  assign T694 = roundingMode_nearest_even & T662;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign T695 = T696 & allRoundExtra;
  assign T696 = roundingMode_nearest_even & T697;
  assign T697 = ~ T662;
  assign T698 = T720 | T699;
  assign T699 = roundUp ? T687 : 55'h0;
  assign roundUp = T707 | T700;
  assign T700 = T701 & 1'h1;
  assign T701 = doIncrSig & roundDirectUp;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign signY = T705 & T702;
  assign T702 = signProd ^ doNegSignSum;
  assign doNegSignSum = isCDominant ? T703 : T378;
  assign T703 = doSubMags & T704;
  assign T704 = ~ isZeroC;
  assign T705 = ~ isZeroY;
  assign isZeroY = T706 == 3'h0;
  assign T706 = T12[6'h38:6'h36];
  assign T707 = T710 | T708;
  assign T708 = T709 & T662;
  assign T709 = doIncrSig & roundingMode_nearest_even;
  assign T710 = T712 | T711;
  assign T711 = doIncrSig & allRound;
  assign T712 = T716 | T713;
  assign T713 = T714 & anyRound;
  assign T714 = T715 & roundDirectUp;
  assign T715 = ~ doIncrSig;
  assign T716 = T717 & T4;
  assign T717 = T718 & T662;
  assign T718 = T719 & roundingMode_nearest_even;
  assign T719 = ~ doIncrSig;
  assign T720 = T725 ? T721 : 55'h0;
  assign T721 = T722 >> 2'h2;
  assign T722 = T12 & T723;
  assign T723 = {1'h0, T724};
  assign T724 = ~ roundMask;
  assign T725 = T727 & T726;
  assign T726 = ~ roundEven;
  assign T727 = ~ roundUp;
  assign T728 = T731 | T729;
  assign T729 = T730 ? sExpX3 : 14'h0;
  assign T730 = sigY3[6'h35:6'h35];
  assign T731 = T733 ? T732 : 14'h0;
  assign T732 = sExpX3 + 14'h1;
  assign T733 = sigY3[6'h36:6'h36];
  assign underflow = commonCase & underflowY;
  assign underflowY = roundInexact & T734;
  assign T734 = T739 | T735;
  assign T735 = T580 <= T736;
  assign T736 = {2'h0, T737};
  assign T737 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign sigX3Shift1 = T738 == 2'h0;
  assign T738 = T12[6'h38:6'h37];
  assign T739 = sExpX3[4'hd:4'hd];
  assign T740 = {invalid, 1'h0};
  assign invalid = T759 | notSigNaN_invalid;
  assign notSigNaN_invalid = T756 | T741;
  assign T741 = T742 & doSubMags;
  assign T742 = T745 & isInfC;
  assign isInfC = isSpecialC & T743;
  assign T743 = T744 ^ 1'h1;
  assign T744 = T162[4'h9:4'h9];
  assign T745 = T751 & T746;
  assign T746 = isInfA | isInfB;
  assign isInfB = isSpecialB & T747;
  assign T747 = T748 ^ 1'h1;
  assign T748 = T168[4'h9:4'h9];
  assign isInfA = isSpecialA & T749;
  assign T749 = T750 ^ 1'h1;
  assign T750 = T165[4'h9:4'h9];
  assign T751 = T754 & T752;
  assign T752 = ~ isNaNB;
  assign isNaNB = isSpecialB & T753;
  assign T753 = T168[4'h9:4'h9];
  assign T754 = ~ isNaNA;
  assign isNaNA = isSpecialA & T755;
  assign T755 = T165[4'h9:4'h9];
  assign T756 = T758 | T757;
  assign T757 = isZeroA & isInfB;
  assign T758 = isInfA & isZeroB;
  assign T759 = T763 | isSigNaNC;
  assign isSigNaNC = isNaNC & T760;
  assign T760 = T761 ^ 1'h1;
  assign T761 = T253[6'h33:6'h33];
  assign isNaNC = isSpecialC & T762;
  assign T762 = T162[4'h9:4'h9];
  assign T763 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T764;
  assign T764 = T765 ^ 1'h1;
  assign T765 = T266[6'h33:6'h33];
  assign isSigNaNA = isNaNA & T766;
  assign T766 = T767 ^ 1'h1;
  assign T767 = T268[6'h33:6'h33];
  assign io_out = T768;
  assign T768 = {signOut, T769};
  assign T769 = {expOut, fractOut};
  assign fractOut = fractY | T770;
  assign T770 = 52'h0 - T771;
  assign T771 = {51'h0, T772};
  assign T772 = isNaNOut | isSatOut;
  assign isSatOut = overflow & T773;
  assign T773 = ~ overflowY_roundMagUp;
  assign overflowY_roundMagUp = T776 | T774;
  assign T774 = roundingMode_max & T775;
  assign T775 = ~ signY;
  assign T776 = roundingMode_nearest_even | T777;
  assign T777 = roundingMode_min & signY;
  assign isNaNOut = T778 | notSigNaN_invalid;
  assign T778 = T779 | isNaNC;
  assign T779 = isNaNA | isNaNB;
  assign fractY = sigX3Shift1 ? T781 : T780;
  assign T780 = sigY3[6'h34:1'h1];
  assign T781 = sigY3[6'h33:1'h0];
  assign expOut = T783 | T782;
  assign T782 = isNaNOut ? 12'he00 : 12'h0;
  assign T783 = T788 | T784;
  assign T784 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = T786 | T785;
  assign T785 = overflow & overflowY_roundMagUp;
  assign T786 = T787 | isInfC;
  assign T787 = isInfA | isInfB;
  assign T788 = T790 | T789;
  assign T789 = isSatOut ? 12'hbff : 12'h0;
  assign T790 = T793 & T791;
  assign T791 = ~ T792;
  assign T792 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T793 = T796 & T794;
  assign T794 = ~ T795;
  assign T795 = isSatOut ? 12'h400 : 12'h0;
  assign T796 = T803 & T797;
  assign T797 = ~ T798;
  assign T798 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign notSpecial_isZeroOut = T802 | totalUnderflowY;
  assign totalUnderflowY = T801 | T799;
  assign T799 = T800 < 12'h3ce;
  assign T800 = sExpY[4'hb:1'h0];
  assign T801 = sExpY[4'hc:4'hc];
  assign T802 = notSpecial_addZeros | isZeroY;
  assign T803 = sExpY[4'hb:1'h0];
  assign signOut = T805 | T804;
  assign T804 = commonCase & signY;
  assign T805 = T809 | T806;
  assign T806 = T807 & opSignC;
  assign T807 = T808 & isSpecialC;
  assign T808 = mulSpecial ^ 1'h1;
  assign T809 = T813 | T810;
  assign T810 = T811 & signProd;
  assign T811 = mulSpecial & T812;
  assign T812 = isSpecialC ^ 1'h1;
  assign T813 = T814 | isNaNOut;
  assign T814 = T815 & opSignC;
  assign T815 = doSubMags ^ 1'h1;
endmodule

module FPUFMAPipe_1(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  wire[1:0] T0;
  reg [2:0] in_rm;
  wire[2:0] T1;
  reg [64:0] in_in3;
  wire[64:0] T2;
  wire[64:0] T3;
  wire[64:0] zero;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg [64:0] in_in2;
  wire[64:0] T10;
  wire[64:0] T11;
  wire T12;
  reg [64:0] in_in1;
  wire[64:0] T13;
  wire[1:0] T14;
  reg [4:0] in_cmd;
  wire[4:0] T15;
  wire[4:0] T16;
  wire[4:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  reg [4:0] R23;
  wire[4:0] T24;
  reg [4:0] R25;
  wire[4:0] T26;
  wire[4:0] res_exc;
  wire[4:0] fma_io_exceptionFlags;
  reg  valid;
  reg  R27;
  wire T28;
  reg [64:0] R29;
  wire[64:0] T30;
  reg [64:0] R31;
  wire[64:0] T32;
  wire[64:0] res_data;
  wire[64:0] fma_io_out;
  reg  R33;
  wire T34;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_rm = {1{$random}};
    in_in3 = {3{$random}};
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_cmd = {1{$random}};
    R23 = {1{$random}};
    R25 = {1{$random}};
    valid = {1{$random}};
    R27 = {1{$random}};
    R29 = {3{$random}};
    R31 = {3{$random}};
    R33 = {1{$random}};
  end
`endif

  assign T0 = in_rm[1'h1:1'h0];
  assign T1 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T2 = T7 ? zero : T3;
  assign T3 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign zero = T4 << 7'h40;
  assign T4 = T6 ^ T5;
  assign T5 = io_in_bits_in2[7'h40:7'h40];
  assign T6 = io_in_bits_in1[7'h40:7'h40];
  assign T7 = io_in_valid & T8;
  assign T8 = T9 ^ 1'h1;
  assign T9 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T10 = T12 ? 65'h8000000000000000 : T11;
  assign T11 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T12 = io_in_valid & io_in_bits_swap23;
  assign T13 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T14 = in_cmd[1'h1:1'h0];
  assign T15 = io_in_valid ? T17 : T16;
  assign T16 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T17 = {3'h0, T18};
  assign T18 = {T20, T19};
  assign T19 = io_in_bits_cmd[1'h0:1'h0];
  assign T20 = T22 & T21;
  assign T21 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T22 = io_in_bits_cmd[1'h1:1'h1];
  assign io_out_bits_exc = R23;
  assign T24 = R27 ? R25 : R23;
  assign T26 = valid ? res_exc : R25;
  assign res_exc = fma_io_exceptionFlags;
  assign T28 = reset ? 1'h0 : valid;
  assign io_out_bits_data = R29;
  assign T30 = R27 ? R31 : R29;
  assign T32 = valid ? res_data : R31;
  assign res_data = fma_io_out;
  assign io_out_valid = R33;
  assign T34 = reset ? 1'h0 : R27;
  mulAddSubRecodedFloatN_1 fma(
       .io_op( T14 ),
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_c( in_in3 ),
       .io_roundingMode( T0 ),
       .io_out( fma_io_out ),
       .io_exceptionFlags( fma_io_exceptionFlags )
  );

  always @(posedge clk) begin
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(T7) begin
      in_in3 <= zero;
    end else if(io_in_valid) begin
      in_in3 <= io_in_bits_in3;
    end
    if(T12) begin
      in_in2 <= 65'h8000000000000000;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_cmd <= T17;
    end else if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(R27) begin
      R23 <= R25;
    end
    if(valid) begin
      R25 <= res_exc;
    end
    valid <= io_in_valid;
    if(reset) begin
      R27 <= 1'h0;
    end else begin
      R27 <= valid;
    end
    if(R27) begin
      R29 <= R31;
    end
    if(valid) begin
      R31 <= res_data;
    end
    if(reset) begin
      R33 <= 1'h0;
    end else begin
      R33 <= R27;
    end
  end
endmodule

module recodedFloatNCompare(
    input [64:0] io_a,
    input [64:0] io_b,
    output io_a_eq_b,
    output io_a_lt_b,
    output io_a_eq_b_invalid,
    output io_a_lt_b_invalid
);

  wire T0;
  wire T1;
  wire[2:0] T2;
  wire[11:0] T3;
  wire T4;
  wire[2:0] T5;
  wire[11:0] T6;
  wire T7;
  wire isSignalingNaNB;
  wire T8;
  wire T9;
  wire[51:0] T10;
  wire isSignalingNaNA;
  wire T11;
  wire T12;
  wire[51:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire magLess;
  wire T17;
  wire T18;
  wire expEqual;
  wire T19;
  wire T20;
  wire T21;
  wire isZeroB;
  wire T22;
  wire isZeroA;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire magEqual;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire signEqual;
  wire T34;
  wire T35;


  assign io_a_lt_b_invalid = T0;
  assign T0 = T4 | T1;
  assign T1 = T2 == 3'h7;
  assign T2 = T3[4'hb:4'h9];
  assign T3 = io_b[6'h3f:6'h34];
  assign T4 = T5 == 3'h7;
  assign T5 = T6[4'hb:4'h9];
  assign T6 = io_a[6'h3f:6'h34];
  assign io_a_eq_b_invalid = T7;
  assign T7 = isSignalingNaNA | isSignalingNaNB;
  assign isSignalingNaNB = T1 & T8;
  assign T8 = T9 ^ 1'h1;
  assign T9 = T10[6'h33:6'h33];
  assign T10 = io_b[6'h33:1'h0];
  assign isSignalingNaNA = T4 & T11;
  assign T11 = T12 ^ 1'h1;
  assign T12 = T13[6'h33:6'h33];
  assign T13 = io_a[6'h33:1'h0];
  assign io_a_lt_b = T14;
  assign T14 = T31 & T15;
  assign T15 = T30 ? T25 : T16;
  assign T16 = T24 ? T20 : magLess;
  assign magLess = T19 | T17;
  assign T17 = expEqual & T18;
  assign T18 = T13 < T10;
  assign expEqual = T6 == T3;
  assign T19 = T6 < T3;
  assign T20 = T21 ^ 1'h1;
  assign T21 = isZeroA & isZeroB;
  assign isZeroB = T22 ^ 1'h1;
  assign T22 = T2 != 3'h0;
  assign isZeroA = T23 ^ 1'h1;
  assign T23 = T5 != 3'h0;
  assign T24 = io_a[7'h40:7'h40];
  assign T25 = T28 & T26;
  assign T26 = magEqual ^ 1'h1;
  assign magEqual = expEqual & T27;
  assign T27 = T13 == T10;
  assign T28 = T24 & T29;
  assign T29 = magLess ^ 1'h1;
  assign T30 = io_b[7'h40:7'h40];
  assign T31 = io_a_lt_b_invalid ^ 1'h1;
  assign io_a_eq_b = T32;
  assign T32 = T34 & T33;
  assign T33 = isZeroA | signEqual;
  assign signEqual = T24 == T30;
  assign T34 = T35 & magEqual;
  assign T35 = T4 ^ 1'h1;
endmodule

module FPToInt(input clk,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output[63:0] io_out_bits_store,
    output[63:0] io_out_bits_toint,
    output[4:0] io_out_bits_exc
);

  reg [64:0] in_in2;
  wire[64:0] T0;
  wire[64:0] T1;
  wire[64:0] T2;
  wire[63:0] T3;
  wire[51:0] T4;
  wire[51:0] T5;
  wire[22:0] T6;
  wire[51:0] T7;
  wire[51:0] T8;
  wire T9;
  wire[2:0] T10;
  wire[11:0] T11;
  wire[11:0] T12;
  wire[11:0] T13;
  wire[11:0] T14;
  wire T15;
  wire[11:0] T16;
  wire[7:0] T17;
  wire T18;
  wire[11:0] T19;
  wire[10:0] T20;
  wire T21;
  wire[11:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire[4:0] T29;
  wire T30;
  wire T31;
  reg [64:0] in_in1;
  wire[64:0] T32;
  wire[64:0] T33;
  wire[64:0] T34;
  wire[63:0] T35;
  wire[51:0] T36;
  wire[51:0] T37;
  wire[22:0] T38;
  wire[51:0] T39;
  wire[51:0] T40;
  wire T41;
  wire[2:0] T42;
  wire[11:0] T43;
  wire[11:0] T44;
  wire[11:0] T45;
  wire[11:0] T46;
  wire T47;
  wire[11:0] T48;
  wire[7:0] T49;
  wire T50;
  wire[11:0] T51;
  wire[10:0] T52;
  wire T53;
  wire[11:0] T54;
  wire T55;
  wire T56;
  wire[4:0] T57;
  wire[4:0] T58;
  wire[4:0] dcmp_exc;
  wire T59;
  wire[2:0] T60;
  wire[2:0] T61;
  wire[1:0] T62;
  wire dcmp_io_a_eq_b_invalid;
  wire dcmp_io_a_lt_b_invalid;
  wire[2:0] T63;
  reg [2:0] in_rm;
  wire[2:0] T64;
  wire T65;
  wire[4:0] T66;
  reg [4:0] in_cmd;
  wire[4:0] T67;
  wire[4:0] T68;
  wire[3:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[10:0] T80;
  wire[11:0] T81;
  wire T82;
  wire T83;
  wire[63:0] T84;
  wire[115:0] T85;
  wire[5:0] T86;
  wire[5:0] T87;
  wire T88;
  wire T89;
  wire[52:0] T90;
  wire[51:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire[1:0] T100;
  wire[2:0] T101;
  wire T102;
  wire[50:0] T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[2:0] T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire[1:0] T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire[10:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[1:0] T139;
  reg [1:0] in_typ;
  wire[1:0] T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire[4:0] T158;
  wire[63:0] T159;
  wire[63:0] T160;
  wire[63:0] T161;
  wire[63:0] unrec_out;
  wire[63:0] unrec_d;
  wire[62:0] T162;
  wire[51:0] T163;
  wire[51:0] T164;
  wire[51:0] T165;
  wire[52:0] T166;
  wire[5:0] T167;
  wire[5:0] T168;
  wire[11:0] T169;
  wire[52:0] T170;
  wire[51:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire[9:0] T175;
  wire T176;
  wire[1:0] T177;
  wire T178;
  wire[2:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire T185;
  wire T186;
  wire[1:0] T187;
  wire T188;
  wire T189;
  wire T190;
  wire[1:0] T191;
  wire[10:0] T192;
  wire[10:0] T193;
  wire[10:0] T194;
  wire[10:0] T195;
  wire[10:0] T196;
  wire T197;
  wire[63:0] T198;
  wire[31:0] unrec_s;
  wire[30:0] T199;
  wire[22:0] T200;
  wire[22:0] T201;
  wire[22:0] T202;
  wire[23:0] T203;
  wire[4:0] T204;
  wire[4:0] T205;
  wire[8:0] T206;
  wire[23:0] T207;
  wire[22:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire[6:0] T212;
  wire T213;
  wire[1:0] T214;
  wire T215;
  wire[2:0] T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire[1:0] T221;
  wire T222;
  wire T223;
  wire[1:0] T224;
  wire T225;
  wire T226;
  wire T227;
  wire[1:0] T228;
  wire[7:0] T229;
  wire[7:0] T230;
  wire[7:0] T231;
  wire[7:0] T232;
  wire[7:0] T233;
  wire T234;
  wire[31:0] T235;
  wire[31:0] T236;
  wire T237;
  reg  in_single;
  wire T238;
  wire[63:0] T239;
  wire[9:0] classify_out;
  wire[9:0] classify_d;
  wire[4:0] T240;
  wire[2:0] T241;
  wire[1:0] T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire[11:0] T248;
  wire T249;
  wire[1:0] T250;
  wire[2:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire[9:0] T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire[1:0] T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[4:0] T270;
  wire[2:0] T271;
  wire[1:0] T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire[1:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[51:0] T283;
  wire T284;
  wire T285;
  wire T286;
  wire[9:0] classify_s;
  wire[4:0] T287;
  wire[2:0] T288;
  wire[1:0] T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire[8:0] T295;
  wire T296;
  wire[1:0] T297;
  wire[2:0] T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire[6:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire[1:0] T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire[4:0] T317;
  wire[2:0] T318;
  wire[1:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire[1:0] T326;
  wire T327;
  wire T328;
  wire T329;
  wire[22:0] T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[63:0] T335;
  wire T336;
  wire[2:0] T337;
  wire[2:0] T338;
  wire[1:0] T339;
  wire dcmp_io_a_eq_b;
  wire dcmp_io_a_lt_b;
  wire[2:0] T340;
  wire[63:0] T341;
  wire[63:0] T342;
  wire[31:0] T343;
  wire[31:0] T344;
  wire[63:0] T345;
  wire[63:0] T346;
  wire[63:0] T347;
  wire[63:0] T348;
  wire[63:0] T349;
  wire[63:0] T350;
  wire T351;
  wire[63:0] T352;
  wire[63:0] T353;
  wire[63:0] T354;
  wire[63:0] T355;
  wire[31:0] T356;
  wire T357;
  wire T358;
  wire T359;
  wire[31:0] T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire[31:0] T369;
  wire T370;
  wire T371;
  reg  valid;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    in_in2 = {3{$random}};
    in_in1 = {3{$random}};
    in_rm = {1{$random}};
    in_cmd = {1{$random}};
    in_typ = {1{$random}};
    in_single = {1{$random}};
    valid = {1{$random}};
  end
`endif

  assign T0 = T25 ? T2 : T1;
  assign T1 = io_in_valid ? io_in_bits_in2 : in_in2;
  assign T2 = {T24, T3};
  assign T3 = {T11, T4};
  assign T4 = T7 | T5;
  assign T5 = T6 << 5'h1d;
  assign T6 = io_in_bits_in2[5'h16:1'h0];
  assign T7 = 52'h0 - T8;
  assign T8 = {51'h0, T9};
  assign T9 = T10 == 3'h7;
  assign T10 = io_in_bits_in2[5'h1f:5'h1d];
  assign T11 = T23 ? T22 : T12;
  assign T12 = T21 ? T19 : T13;
  assign T13 = T18 ? T16 : T14;
  assign T14 = T15 ? 12'hc00 : 12'he00;
  assign T15 = T10 < 3'h7;
  assign T16 = {4'h8, T17};
  assign T17 = io_in_bits_in2[5'h1e:5'h17];
  assign T18 = T10 < 3'h6;
  assign T19 = {1'h0, T20};
  assign T20 = {3'h7, T17};
  assign T21 = T10 < 3'h4;
  assign T22 = {4'h0, T17};
  assign T23 = T10 < 3'h1;
  assign T24 = io_in_bits_in2[6'h20:6'h20];
  assign T25 = io_in_valid & T26;
  assign T26 = T30 & T27;
  assign T27 = T28 == 1'h0;
  assign T28 = T29 == 5'hc;
  assign T29 = io_in_bits_cmd & 5'hc;
  assign T30 = io_in_bits_single & T31;
  assign T31 = io_in_bits_ldst ^ 1'h1;
  assign T32 = T25 ? T34 : T33;
  assign T33 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign T34 = {T56, T35};
  assign T35 = {T43, T36};
  assign T36 = T39 | T37;
  assign T37 = T38 << 5'h1d;
  assign T38 = io_in_bits_in1[5'h16:1'h0];
  assign T39 = 52'h0 - T40;
  assign T40 = {51'h0, T41};
  assign T41 = T42 == 3'h7;
  assign T42 = io_in_bits_in1[5'h1f:5'h1d];
  assign T43 = T55 ? T54 : T44;
  assign T44 = T53 ? T51 : T45;
  assign T45 = T50 ? T48 : T46;
  assign T46 = T47 ? 12'hc00 : 12'he00;
  assign T47 = T42 < 3'h7;
  assign T48 = {4'h8, T49};
  assign T49 = io_in_bits_in1[5'h1e:5'h17];
  assign T50 = T42 < 3'h6;
  assign T51 = {1'h0, T52};
  assign T52 = {3'h7, T49};
  assign T53 = T42 < 3'h4;
  assign T54 = {4'h0, T49};
  assign T55 = T42 < 3'h1;
  assign T56 = io_in_bits_in1[6'h20:6'h20];
  assign io_out_bits_exc = T57;
  assign T57 = T157 ? T68 : T58;
  assign T58 = T65 ? dcmp_exc : 5'h0;
  assign dcmp_exc = T59 << 3'h4;
  assign T59 = T60 != 3'h0;
  assign T60 = T63 & T61;
  assign T61 = {1'h0, T62};
  assign T62 = {dcmp_io_a_lt_b_invalid, dcmp_io_a_eq_b_invalid};
  assign T63 = ~ in_rm;
  assign T64 = io_in_valid ? io_in_bits_rm : in_rm;
  assign T65 = T66 == 5'h4;
  assign T66 = in_cmd & 5'hc;
  assign T67 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign T68 = {T72, T69};
  assign T69 = {3'h0, T70};
  assign T70 = T99 & T71;
  assign T71 = T72 ^ 1'h1;
  assign T72 = T155 | T73;
  assign T73 = T154 ? T148 : T74;
  assign T74 = T147 ? T141 : T75;
  assign T75 = T138 ? T132 : T76;
  assign T76 = T88 ? 1'h0 : T77;
  assign T77 = T131 ? T127 : T78;
  assign T78 = T126 ? T82 : T79;
  assign T79 = 11'h40 <= T80;
  assign T80 = T81[4'ha:1'h0];
  assign T81 = in_in1[6'h3f:6'h34];
  assign T82 = T93 | T83;
  assign T83 = T84 != 64'h0;
  assign T84 = T85[7'h73:6'h34];
  assign T85 = T90 << T86;
  assign T86 = T88 ? 6'h0 : T87;
  assign T87 = T81[3'h5:1'h0];
  assign T88 = T89 ^ 1'h1;
  assign T89 = T81[4'hb:4'hb];
  assign T90 = {T92, T91};
  assign T91 = in_in1[6'h33:1'h0];
  assign T92 = T88 ^ 1'h1;
  assign T93 = T125 | T94;
  assign T94 = T124 ? T113 : T95;
  assign T95 = T112 ? T111 : T96;
  assign T96 = T110 ? T97 : 1'h0;
  assign T97 = T108 & T98;
  assign T98 = T88 ? T105 : T99;
  assign T99 = T100 != 2'h0;
  assign T100 = T101[1'h1:1'h0];
  assign T101 = {T104, T102};
  assign T102 = T103 != 51'h0;
  assign T103 = T85[6'h32:1'h0];
  assign T104 = T85[6'h34:6'h33];
  assign T105 = T106 ^ 1'h1;
  assign T106 = T107 == 3'h0;
  assign T107 = T81[4'hb:4'h9];
  assign T108 = T109 ^ 1'h1;
  assign T109 = in_in1[7'h40:7'h40];
  assign T110 = in_rm == 3'h3;
  assign T111 = T109 & T98;
  assign T112 = in_rm == 3'h2;
  assign T113 = T88 ? T119 : T114;
  assign T114 = T117 | T115;
  assign T115 = T116 == 2'h3;
  assign T116 = T101[1'h1:1'h0];
  assign T117 = T118 == 2'h3;
  assign T118 = T101[2'h2:1'h1];
  assign T119 = T120 & T99;
  assign T120 = T121 ^ 1'h1;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T123 == 11'h7ff;
  assign T123 = T81[4'ha:1'h0];
  assign T124 = in_rm == 3'h0;
  assign T125 = T109 ^ 1'h1;
  assign T126 = T80 == 11'h3f;
  assign T127 = T130 & T128;
  assign T128 = T94 & T129;
  assign T129 = T84 == 64'hffffffffffffffff;
  assign T130 = T109 ^ 1'h1;
  assign T131 = T80 == 11'h3e;
  assign T132 = T88 ? T137 : T133;
  assign T133 = T109 | T134;
  assign T134 = T136 ? T128 : T135;
  assign T135 = 11'h40 <= T80;
  assign T136 = T80 == 11'h3f;
  assign T137 = T109 & T94;
  assign T138 = T139 == 2'h2;
  assign T139 = in_typ ^ 2'h1;
  assign T140 = io_in_valid ? io_in_bits_typ : in_typ;
  assign T141 = T88 ? 1'h0 : T142;
  assign T142 = T146 ? T127 : T143;
  assign T143 = T145 ? T82 : T144;
  assign T144 = 11'h20 <= T80;
  assign T145 = T80 == 11'h1f;
  assign T146 = T80 == 11'h1e;
  assign T147 = T139 == 2'h1;
  assign T148 = T88 ? T153 : T149;
  assign T149 = T109 | T150;
  assign T150 = T152 ? T128 : T151;
  assign T151 = 11'h20 <= T80;
  assign T152 = T80 == 11'h1f;
  assign T153 = T109 & T94;
  assign T154 = T139 == 2'h0;
  assign T155 = T156 == 2'h3;
  assign T156 = T81[4'hb:4'ha];
  assign T157 = T158 == 5'h8;
  assign T158 = in_cmd & 5'hc;
  assign io_out_bits_toint = T159;
  assign T159 = T157 ? T341 : T160;
  assign T160 = T65 ? T335 : T161;
  assign T161 = T334 ? T239 : unrec_out;
  assign unrec_out = in_single ? T198 : unrec_d;
  assign unrec_d = {T197, T162};
  assign T162 = {T192, T163};
  assign T163 = T180 ? T171 : T164;
  assign T164 = T172 ? T165 : 52'h0;
  assign T165 = T166[6'h33:1'h0];
  assign T166 = T170 >> T167;
  assign T167 = 6'h2 - T168;
  assign T168 = T169[3'h5:1'h0];
  assign T169 = in_in1[6'h3f:6'h34];
  assign T170 = {1'h1, T171};
  assign T171 = in_in1[6'h33:1'h0];
  assign T172 = T178 | T173;
  assign T173 = T176 & T174;
  assign T174 = T175 < 10'h2;
  assign T175 = T169[4'h9:1'h0];
  assign T176 = T177 == 2'h1;
  assign T177 = T169[4'hb:4'ha];
  assign T178 = T179 == 3'h1;
  assign T179 = T169[4'hb:4'h9];
  assign T180 = T185 | T181;
  assign T181 = T183 & T182;
  assign T182 = T169[4'h9:4'h9];
  assign T183 = T184 == 2'h3;
  assign T184 = T169[4'hb:4'ha];
  assign T185 = T188 | T186;
  assign T186 = T187 == 2'h2;
  assign T187 = T169[4'hb:4'ha];
  assign T188 = T190 & T189;
  assign T189 = T174 ^ 1'h1;
  assign T190 = T191 == 2'h1;
  assign T191 = T169[4'hb:4'ha];
  assign T192 = T185 ? T195 : T193;
  assign T193 = 11'h0 - T194;
  assign T194 = {10'h0, T183};
  assign T195 = T196 - 11'h401;
  assign T196 = T169[4'ha:1'h0];
  assign T197 = in_in1[7'h40:7'h40];
  assign T198 = {T235, unrec_s};
  assign unrec_s = {T234, T199};
  assign T199 = {T229, T200};
  assign T200 = T217 ? T208 : T201;
  assign T201 = T209 ? T202 : 23'h0;
  assign T202 = T203[5'h16:1'h0];
  assign T203 = T207 >> T204;
  assign T204 = 5'h2 - T205;
  assign T205 = T206[3'h4:1'h0];
  assign T206 = in_in1[5'h1f:5'h17];
  assign T207 = {1'h1, T208};
  assign T208 = in_in1[5'h16:1'h0];
  assign T209 = T215 | T210;
  assign T210 = T213 & T211;
  assign T211 = T212 < 7'h2;
  assign T212 = T206[3'h6:1'h0];
  assign T213 = T214 == 2'h1;
  assign T214 = T206[4'h8:3'h7];
  assign T215 = T216 == 3'h1;
  assign T216 = T206[4'h8:3'h6];
  assign T217 = T222 | T218;
  assign T218 = T220 & T219;
  assign T219 = T206[3'h6:3'h6];
  assign T220 = T221 == 2'h3;
  assign T221 = T206[4'h8:3'h7];
  assign T222 = T225 | T223;
  assign T223 = T224 == 2'h2;
  assign T224 = T206[4'h8:3'h7];
  assign T225 = T227 & T226;
  assign T226 = T211 ^ 1'h1;
  assign T227 = T228 == 2'h1;
  assign T228 = T206[4'h8:3'h7];
  assign T229 = T222 ? T232 : T230;
  assign T230 = 8'h0 - T231;
  assign T231 = {7'h0, T220};
  assign T232 = T233 - 8'h81;
  assign T233 = T206[3'h7:1'h0];
  assign T234 = in_in1[6'h20:6'h20];
  assign T235 = 32'h0 - T236;
  assign T236 = {31'h0, T237};
  assign T237 = unrec_s[5'h1f:5'h1f];
  assign T238 = io_in_valid ? io_in_bits_single : in_single;
  assign T239 = {54'h0, classify_out};
  assign classify_out = in_single ? classify_s : classify_d;
  assign classify_d = {T270, T240};
  assign T240 = {T265, T241};
  assign T241 = {T260, T242};
  assign T242 = {T252, T243};
  assign T243 = T245 & T244;
  assign T244 = in_in1[7'h40:7'h40];
  assign T245 = T249 & T246;
  assign T246 = T247 ^ 1'h1;
  assign T247 = T248[4'h9:4'h9];
  assign T248 = in_in1[6'h3f:6'h34];
  assign T249 = T250 == 2'h3;
  assign T250 = T251[2'h2:1'h1];
  assign T251 = T248[4'hb:4'h9];
  assign T252 = T253 & T244;
  assign T253 = T255 | T254;
  assign T254 = T250 == 2'h2;
  assign T255 = T259 & T256;
  assign T256 = T257 ^ 1'h1;
  assign T257 = T258 < 10'h2;
  assign T258 = T248[4'h9:1'h0];
  assign T259 = T250 == 2'h1;
  assign T260 = T261 & T244;
  assign T261 = T264 | T262;
  assign T262 = T263 & T257;
  assign T263 = T250 == 2'h1;
  assign T264 = T251 == 3'h1;
  assign T265 = {T268, T266};
  assign T266 = T267 & T244;
  assign T267 = T251 == 3'h0;
  assign T268 = T267 & T269;
  assign T269 = T244 ^ 1'h1;
  assign T270 = {T279, T271};
  assign T271 = {T277, T272};
  assign T272 = {T275, T273};
  assign T273 = T261 & T274;
  assign T274 = T244 ^ 1'h1;
  assign T275 = T253 & T276;
  assign T276 = T244 ^ 1'h1;
  assign T277 = T245 & T278;
  assign T278 = T244 ^ 1'h1;
  assign T279 = {T285, T280};
  assign T280 = T284 & T281;
  assign T281 = T282 ^ 1'h1;
  assign T282 = T283[6'h33:6'h33];
  assign T283 = in_in1[6'h33:1'h0];
  assign T284 = T251 == 3'h7;
  assign T285 = T284 & T286;
  assign T286 = T283[6'h33:6'h33];
  assign classify_s = {T317, T287};
  assign T287 = {T312, T288};
  assign T288 = {T307, T289};
  assign T289 = {T299, T290};
  assign T290 = T292 & T291;
  assign T291 = in_in1[6'h20:6'h20];
  assign T292 = T296 & T293;
  assign T293 = T294 ^ 1'h1;
  assign T294 = T295[3'h6:3'h6];
  assign T295 = in_in1[5'h1f:5'h17];
  assign T296 = T297 == 2'h3;
  assign T297 = T298[2'h2:1'h1];
  assign T298 = T295[4'h8:3'h6];
  assign T299 = T300 & T291;
  assign T300 = T302 | T301;
  assign T301 = T297 == 2'h2;
  assign T302 = T306 & T303;
  assign T303 = T304 ^ 1'h1;
  assign T304 = T305 < 7'h2;
  assign T305 = T295[3'h6:1'h0];
  assign T306 = T297 == 2'h1;
  assign T307 = T308 & T291;
  assign T308 = T311 | T309;
  assign T309 = T310 & T304;
  assign T310 = T297 == 2'h1;
  assign T311 = T298 == 3'h1;
  assign T312 = {T315, T313};
  assign T313 = T314 & T291;
  assign T314 = T298 == 3'h0;
  assign T315 = T314 & T316;
  assign T316 = T291 ^ 1'h1;
  assign T317 = {T326, T318};
  assign T318 = {T324, T319};
  assign T319 = {T322, T320};
  assign T320 = T308 & T321;
  assign T321 = T291 ^ 1'h1;
  assign T322 = T300 & T323;
  assign T323 = T291 ^ 1'h1;
  assign T324 = T292 & T325;
  assign T325 = T291 ^ 1'h1;
  assign T326 = {T332, T327};
  assign T327 = T331 & T328;
  assign T328 = T329 ^ 1'h1;
  assign T329 = T330[5'h16:5'h16];
  assign T330 = in_in1[5'h16:1'h0];
  assign T331 = T298 == 3'h7;
  assign T332 = T331 & T333;
  assign T333 = T330[5'h16:5'h16];
  assign T334 = in_rm[1'h0:1'h0];
  assign T335 = {63'h0, T336};
  assign T336 = T337 != 3'h0;
  assign T337 = T340 & T338;
  assign T338 = {1'h0, T339};
  assign T339 = {dcmp_io_a_lt_b, dcmp_io_a_eq_b};
  assign T340 = ~ in_rm;
  assign T341 = T371 ? T345 : T342;
  assign T342 = {T369, T343};
  assign T343 = T344;
  assign T344 = T345[5'h1f:1'h0];
  assign T345 = T72 ? T352 : T346;
  assign T346 = T347;
  assign T347 = T351 ? T350 : T348;
  assign T348 = T109 ? T349 : T84;
  assign T349 = ~ T84;
  assign T350 = T348 + 64'h1;
  assign T351 = T94 ^ T109;
  assign T352 = T367 ? 64'h8000000000000000 : T353;
  assign T353 = T365 ? 64'hffffffff80000000 : T354;
  assign T354 = T362 ? 64'h7fffffffffffffff : T355;
  assign T355 = {T360, T356};
  assign T356 = T357 ? 32'h7fffffff : 32'hffffffff;
  assign T357 = T359 & T358;
  assign T358 = T109 ^ 1'h1;
  assign T359 = T139 == 2'h1;
  assign T360 = T361 ? 32'hffffffff : 32'h0;
  assign T361 = T356[5'h1f:5'h1f];
  assign T362 = T364 & T363;
  assign T363 = T109 ^ 1'h1;
  assign T364 = T139 == 2'h3;
  assign T365 = T366 & T109;
  assign T366 = T139 == 2'h1;
  assign T367 = T368 & T109;
  assign T368 = T139 == 2'h3;
  assign T369 = T370 ? 32'hffffffff : 32'h0;
  assign T370 = T343[5'h1f:5'h1f];
  assign T371 = in_typ[1'h1:1'h1];
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_lt = dcmp_io_a_lt_b;
  assign io_out_valid = valid;
  recodedFloatNCompare dcmp(
       .io_a( in_in1 ),
       .io_b( in_in2 ),
       .io_a_eq_b( dcmp_io_a_eq_b ),
       .io_a_lt_b( dcmp_io_a_lt_b ),
       .io_a_eq_b_invalid( dcmp_io_a_eq_b_invalid ),
       .io_a_lt_b_invalid( dcmp_io_a_lt_b_invalid )
  );

  always @(posedge clk) begin
    if(T25) begin
      in_in2 <= T2;
    end else if(io_in_valid) begin
      in_in2 <= io_in_bits_in2;
    end
    if(T25) begin
      in_in1 <= T34;
    end else if(io_in_valid) begin
      in_in1 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      in_rm <= io_in_bits_rm;
    end
    if(io_in_valid) begin
      in_cmd <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      in_typ <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      in_single <= io_in_bits_single;
    end
    valid <= io_in_valid;
  end
endmodule

module IntToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc
);

  reg [4:0] R0;
  wire[4:0] T1;
  reg [4:0] R2;
  wire[4:0] T3;
  wire[4:0] mux_exc;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[1:0] T7;
  wire T8;
  wire[1:0] T9;
  wire[2:0] T10;
  wire T11;
  wire[38:0] T12;
  wire[126:0] T13;
  wire[5:0] T14;
  wire[5:0] T15;
  wire[5:0] T16;
  wire[5:0] T17;
  wire[5:0] T18;
  wire[5:0] T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire[5:0] T22;
  wire[5:0] T23;
  wire[5:0] T24;
  wire[5:0] T25;
  wire[5:0] T26;
  wire[5:0] T27;
  wire[5:0] T28;
  wire[5:0] T29;
  wire[5:0] T30;
  wire[5:0] T31;
  wire[5:0] T32;
  wire[5:0] T33;
  wire[5:0] T34;
  wire[5:0] T35;
  wire[5:0] T36;
  wire[5:0] T37;
  wire[5:0] T38;
  wire[5:0] T39;
  wire[5:0] T40;
  wire[5:0] T41;
  wire[5:0] T42;
  wire[5:0] T43;
  wire[5:0] T44;
  wire[5:0] T45;
  wire[5:0] T46;
  wire[4:0] T47;
  wire[4:0] T48;
  wire[4:0] T49;
  wire[4:0] T50;
  wire[4:0] T51;
  wire[4:0] T52;
  wire[4:0] T53;
  wire[4:0] T54;
  wire[4:0] T55;
  wire[4:0] T56;
  wire[4:0] T57;
  wire[4:0] T58;
  wire[4:0] T59;
  wire[4:0] T60;
  wire[4:0] T61;
  wire[4:0] T62;
  wire[3:0] T63;
  wire[3:0] T64;
  wire[3:0] T65;
  wire[3:0] T66;
  wire[3:0] T67;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[2:0] T71;
  wire[2:0] T72;
  wire[2:0] T73;
  wire[2:0] T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire T77;
  wire[63:0] T78;
  wire[63:0] T79;
  wire[63:0] T80;
  wire[31:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  reg [64:0] R84;
  wire[64:0] T85;
  wire[63:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  reg [1:0] R92;
  wire[1:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire[1:0] T161;
  wire T162;
  reg  R163;
  wire T164;
  wire T165;
  wire[4:0] T166;
  reg [4:0] R167;
  wire[4:0] T168;
  wire[4:0] T169;
  wire[1:0] T170;
  wire T171;
  wire[1:0] T172;
  wire[2:0] T173;
  wire T174;
  wire[9:0] T175;
  wire[126:0] T176;
  wire[5:0] T177;
  wire[5:0] T178;
  wire[5:0] T179;
  wire[5:0] T180;
  wire[5:0] T181;
  wire[5:0] T182;
  wire[5:0] T183;
  wire[5:0] T184;
  wire[5:0] T185;
  wire[5:0] T186;
  wire[5:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[5:0] T190;
  wire[5:0] T191;
  wire[5:0] T192;
  wire[5:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire[5:0] T196;
  wire[5:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[5:0] T200;
  wire[5:0] T201;
  wire[5:0] T202;
  wire[5:0] T203;
  wire[5:0] T204;
  wire[5:0] T205;
  wire[5:0] T206;
  wire[5:0] T207;
  wire[5:0] T208;
  wire[5:0] T209;
  wire[4:0] T210;
  wire[4:0] T211;
  wire[4:0] T212;
  wire[4:0] T213;
  wire[4:0] T214;
  wire[4:0] T215;
  wire[4:0] T216;
  wire[4:0] T217;
  wire[4:0] T218;
  wire[4:0] T219;
  wire[4:0] T220;
  wire[4:0] T221;
  wire[4:0] T222;
  wire[4:0] T223;
  wire[4:0] T224;
  wire[4:0] T225;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[3:0] T230;
  wire[3:0] T231;
  wire[3:0] T232;
  wire[3:0] T233;
  wire[2:0] T234;
  wire[2:0] T235;
  wire[2:0] T236;
  wire[2:0] T237;
  wire[1:0] T238;
  wire[1:0] T239;
  wire T240;
  wire[63:0] T241;
  wire[63:0] T242;
  wire[63:0] T243;
  wire[31:0] T244;
  wire[63:0] T245;
  wire[63:0] T246;
  wire[63:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire[1:0] T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire T321;
  wire T322;
  reg  R323;
  wire T324;
  reg  R325;
  wire T326;
  reg [64:0] R327;
  wire[64:0] T328;
  reg [64:0] R329;
  wire[64:0] T330;
  wire[64:0] mux_data;
  wire[64:0] T331;
  wire[64:0] T332;
  wire[64:0] T333;
  wire[64:0] T334;
  wire[63:0] T335;
  wire[51:0] T336;
  wire[51:0] T337;
  wire[51:0] T338;
  wire[126:0] T339;
  wire[5:0] T340;
  wire[5:0] T341;
  wire[5:0] T342;
  wire[5:0] T343;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[5:0] T349;
  wire[5:0] T350;
  wire[5:0] T351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[5:0] T357;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[5:0] T365;
  wire[5:0] T366;
  wire[5:0] T367;
  wire[5:0] T368;
  wire[5:0] T369;
  wire[5:0] T370;
  wire[5:0] T371;
  wire[5:0] T372;
  wire[4:0] T373;
  wire[4:0] T374;
  wire[4:0] T375;
  wire[4:0] T376;
  wire[4:0] T377;
  wire[4:0] T378;
  wire[4:0] T379;
  wire[4:0] T380;
  wire[4:0] T381;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire[4:0] T385;
  wire[4:0] T386;
  wire[4:0] T387;
  wire[4:0] T388;
  wire[3:0] T389;
  wire[3:0] T390;
  wire[3:0] T391;
  wire[3:0] T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[2:0] T397;
  wire[2:0] T398;
  wire[2:0] T399;
  wire[2:0] T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire T403;
  wire[63:0] T404;
  wire[63:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire[10:0] T469;
  wire[11:0] T470;
  wire[11:0] T471;
  wire[9:0] T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire[1:0] T477;
  wire[11:0] T478;
  wire[11:0] T479;
  wire[10:0] T480;
  wire[10:0] T481;
  wire[10:0] T482;
  wire[1:0] T483;
  wire T484;
  wire T485;
  wire T486;
  wire[11:0] T487;
  wire[11:0] T488;
  wire[11:0] T489;
  wire[11:0] T490;
  wire[5:0] T491;
  wire T492;
  wire[64:0] T493;
  wire[32:0] T494;
  wire[31:0] T495;
  wire[22:0] T496;
  wire[22:0] T497;
  wire[22:0] T498;
  wire[62:0] T499;
  wire[4:0] T500;
  wire[4:0] T501;
  wire[4:0] T502;
  wire[4:0] T503;
  wire[4:0] T504;
  wire[4:0] T505;
  wire[4:0] T506;
  wire[4:0] T507;
  wire[4:0] T508;
  wire[4:0] T509;
  wire[4:0] T510;
  wire[4:0] T511;
  wire[4:0] T512;
  wire[4:0] T513;
  wire[4:0] T514;
  wire[4:0] T515;
  wire[4:0] T516;
  wire[3:0] T517;
  wire[3:0] T518;
  wire[3:0] T519;
  wire[3:0] T520;
  wire[3:0] T521;
  wire[3:0] T522;
  wire[3:0] T523;
  wire[3:0] T524;
  wire[2:0] T525;
  wire[2:0] T526;
  wire[2:0] T527;
  wire[2:0] T528;
  wire[1:0] T529;
  wire[1:0] T530;
  wire T531;
  wire[31:0] T532;
  wire[31:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire[7:0] T565;
  wire[8:0] T566;
  wire[8:0] T567;
  wire[6:0] T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire[1:0] T573;
  wire[8:0] T574;
  wire[8:0] T575;
  wire[7:0] T576;
  wire[7:0] T577;
  wire[7:0] T578;
  wire[1:0] T579;
  wire T580;
  wire T581;
  wire T582;
  wire[8:0] T583;
  wire[8:0] T584;
  wire[8:0] T585;
  wire[8:0] T586;
  wire[4:0] T587;
  wire T588;
  wire[64:0] T589;
  wire[32:0] T590;
  wire[31:0] T591;
  wire[22:0] T592;
  wire[24:0] T593;
  wire[24:0] T594;
  wire[23:0] T595;
  wire[24:0] T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  reg [2:0] R603;
  wire[2:0] T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire T610;
  wire[1:0] T611;
  wire T612;
  wire[8:0] T613;
  wire[7:0] T614;
  wire[7:0] T615;
  wire[7:0] T616;
  wire T617;
  wire[7:0] T618;
  wire[6:0] T619;
  wire[5:0] T620;
  wire T621;
  wire[64:0] T622;
  wire[63:0] T623;
  wire[51:0] T624;
  wire[53:0] T625;
  wire[53:0] T626;
  wire[52:0] T627;
  wire[53:0] T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire[1:0] T639;
  wire T640;
  wire[1:0] T641;
  wire T642;
  wire[11:0] T643;
  wire[10:0] T644;
  wire[10:0] T645;
  wire[10:0] T646;
  wire T647;
  wire[10:0] T648;
  wire[9:0] T649;
  wire[5:0] T650;
  wire T651;
  reg  R652;
  wire T653;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R2 = {1{$random}};
    R84 = {3{$random}};
    R92 = {1{$random}};
    R163 = {1{$random}};
    R167 = {1{$random}};
    R323 = {1{$random}};
    R325 = {1{$random}};
    R327 = {3{$random}};
    R329 = {3{$random}};
    R603 = {1{$random}};
    R652 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R325 ? R2 : R0;
  assign T3 = R323 ? mux_exc : R2;
  assign mux_exc = T4;
  assign T4 = T321 ? T169 : T5;
  assign T5 = T162 ? T6 : 5'h0;
  assign T6 = {3'h0, T7};
  assign T7 = {1'h0, T8};
  assign T8 = T9 != 2'h0;
  assign T9 = T10[1'h1:1'h0];
  assign T10 = {T161, T11};
  assign T11 = T12 != 39'h0;
  assign T12 = T13[6'h26:1'h0];
  assign T13 = T79 << T14;
  assign T14 = ~ T15;
  assign T15 = T160 ? 6'h3f : T16;
  assign T16 = T159 ? 6'h3e : T17;
  assign T17 = T158 ? 6'h3d : T18;
  assign T18 = T157 ? 6'h3c : T19;
  assign T19 = T156 ? 6'h3b : T20;
  assign T20 = T155 ? 6'h3a : T21;
  assign T21 = T154 ? 6'h39 : T22;
  assign T22 = T153 ? 6'h38 : T23;
  assign T23 = T152 ? 6'h37 : T24;
  assign T24 = T151 ? 6'h36 : T25;
  assign T25 = T150 ? 6'h35 : T26;
  assign T26 = T149 ? 6'h34 : T27;
  assign T27 = T148 ? 6'h33 : T28;
  assign T28 = T147 ? 6'h32 : T29;
  assign T29 = T146 ? 6'h31 : T30;
  assign T30 = T145 ? 6'h30 : T31;
  assign T31 = T144 ? 6'h2f : T32;
  assign T32 = T143 ? 6'h2e : T33;
  assign T33 = T142 ? 6'h2d : T34;
  assign T34 = T141 ? 6'h2c : T35;
  assign T35 = T140 ? 6'h2b : T36;
  assign T36 = T139 ? 6'h2a : T37;
  assign T37 = T138 ? 6'h29 : T38;
  assign T38 = T137 ? 6'h28 : T39;
  assign T39 = T136 ? 6'h27 : T40;
  assign T40 = T135 ? 6'h26 : T41;
  assign T41 = T134 ? 6'h25 : T42;
  assign T42 = T133 ? 6'h24 : T43;
  assign T43 = T132 ? 6'h23 : T44;
  assign T44 = T131 ? 6'h22 : T45;
  assign T45 = T130 ? 6'h21 : T46;
  assign T46 = T129 ? 6'h20 : T47;
  assign T47 = T128 ? 5'h1f : T48;
  assign T48 = T127 ? 5'h1e : T49;
  assign T49 = T126 ? 5'h1d : T50;
  assign T50 = T125 ? 5'h1c : T51;
  assign T51 = T124 ? 5'h1b : T52;
  assign T52 = T123 ? 5'h1a : T53;
  assign T53 = T122 ? 5'h19 : T54;
  assign T54 = T121 ? 5'h18 : T55;
  assign T55 = T120 ? 5'h17 : T56;
  assign T56 = T119 ? 5'h16 : T57;
  assign T57 = T118 ? 5'h15 : T58;
  assign T58 = T117 ? 5'h14 : T59;
  assign T59 = T116 ? 5'h13 : T60;
  assign T60 = T115 ? 5'h12 : T61;
  assign T61 = T114 ? 5'h11 : T62;
  assign T62 = T113 ? 5'h10 : T63;
  assign T63 = T112 ? 4'hf : T64;
  assign T64 = T111 ? 4'he : T65;
  assign T65 = T110 ? 4'hd : T66;
  assign T66 = T109 ? 4'hc : T67;
  assign T67 = T108 ? 4'hb : T68;
  assign T68 = T107 ? 4'ha : T69;
  assign T69 = T106 ? 4'h9 : T70;
  assign T70 = T105 ? 4'h8 : T71;
  assign T71 = T104 ? 3'h7 : T72;
  assign T72 = T103 ? 3'h6 : T73;
  assign T73 = T102 ? 3'h5 : T74;
  assign T74 = T101 ? 3'h4 : T75;
  assign T75 = T100 ? 2'h3 : T76;
  assign T76 = T99 ? 2'h2 : T77;
  assign T77 = T78[1'h1:1'h1];
  assign T78 = T79[6'h3f:1'h0];
  assign T79 = T96 ? T82 : T80;
  assign T80 = {32'h0, T81};
  assign T81 = T82[5'h1f:1'h0];
  assign T82 = T87 ? T86 : T83;
  assign T83 = R84[6'h3f:1'h0];
  assign T85 = io_in_valid ? io_in_bits_in1 : R84;
  assign T86 = 64'h0 - T83;
  assign T87 = T95 ? T94 : T88;
  assign T88 = T90 ? T89 : 1'h0;
  assign T89 = T83[6'h3f:6'h3f];
  assign T90 = T91 == 2'h3;
  assign T91 = R92 ^ 2'h1;
  assign T93 = io_in_valid ? io_in_bits_typ : R92;
  assign T94 = T83[5'h1f:5'h1f];
  assign T95 = T91 == 2'h1;
  assign T96 = T98 | T97;
  assign T97 = T91 == 2'h2;
  assign T98 = T91 == 2'h3;
  assign T99 = T78[2'h2:2'h2];
  assign T100 = T78[2'h3:2'h3];
  assign T101 = T78[3'h4:3'h4];
  assign T102 = T78[3'h5:3'h5];
  assign T103 = T78[3'h6:3'h6];
  assign T104 = T78[3'h7:3'h7];
  assign T105 = T78[4'h8:4'h8];
  assign T106 = T78[4'h9:4'h9];
  assign T107 = T78[4'ha:4'ha];
  assign T108 = T78[4'hb:4'hb];
  assign T109 = T78[4'hc:4'hc];
  assign T110 = T78[4'hd:4'hd];
  assign T111 = T78[4'he:4'he];
  assign T112 = T78[4'hf:4'hf];
  assign T113 = T78[5'h10:5'h10];
  assign T114 = T78[5'h11:5'h11];
  assign T115 = T78[5'h12:5'h12];
  assign T116 = T78[5'h13:5'h13];
  assign T117 = T78[5'h14:5'h14];
  assign T118 = T78[5'h15:5'h15];
  assign T119 = T78[5'h16:5'h16];
  assign T120 = T78[5'h17:5'h17];
  assign T121 = T78[5'h18:5'h18];
  assign T122 = T78[5'h19:5'h19];
  assign T123 = T78[5'h1a:5'h1a];
  assign T124 = T78[5'h1b:5'h1b];
  assign T125 = T78[5'h1c:5'h1c];
  assign T126 = T78[5'h1d:5'h1d];
  assign T127 = T78[5'h1e:5'h1e];
  assign T128 = T78[5'h1f:5'h1f];
  assign T129 = T78[6'h20:6'h20];
  assign T130 = T78[6'h21:6'h21];
  assign T131 = T78[6'h22:6'h22];
  assign T132 = T78[6'h23:6'h23];
  assign T133 = T78[6'h24:6'h24];
  assign T134 = T78[6'h25:6'h25];
  assign T135 = T78[6'h26:6'h26];
  assign T136 = T78[6'h27:6'h27];
  assign T137 = T78[6'h28:6'h28];
  assign T138 = T78[6'h29:6'h29];
  assign T139 = T78[6'h2a:6'h2a];
  assign T140 = T78[6'h2b:6'h2b];
  assign T141 = T78[6'h2c:6'h2c];
  assign T142 = T78[6'h2d:6'h2d];
  assign T143 = T78[6'h2e:6'h2e];
  assign T144 = T78[6'h2f:6'h2f];
  assign T145 = T78[6'h30:6'h30];
  assign T146 = T78[6'h31:6'h31];
  assign T147 = T78[6'h32:6'h32];
  assign T148 = T78[6'h33:6'h33];
  assign T149 = T78[6'h34:6'h34];
  assign T150 = T78[6'h35:6'h35];
  assign T151 = T78[6'h36:6'h36];
  assign T152 = T78[6'h37:6'h37];
  assign T153 = T78[6'h38:6'h38];
  assign T154 = T78[6'h39:6'h39];
  assign T155 = T78[6'h3a:6'h3a];
  assign T156 = T78[6'h3b:6'h3b];
  assign T157 = T78[6'h3c:6'h3c];
  assign T158 = T78[6'h3d:6'h3d];
  assign T159 = T78[6'h3e:6'h3e];
  assign T160 = T78[6'h3f:6'h3f];
  assign T161 = T13[6'h28:6'h27];
  assign T162 = T165 & R163;
  assign T164 = io_in_valid ? io_in_bits_single : R163;
  assign T165 = T166 == 5'h0;
  assign T166 = R167 & 5'h4;
  assign T168 = io_in_valid ? io_in_bits_cmd : R167;
  assign T169 = {3'h0, T170};
  assign T170 = {1'h0, T171};
  assign T171 = T172 != 2'h0;
  assign T172 = T173[1'h1:1'h0];
  assign T173 = {T320, T174};
  assign T174 = T175 != 10'h0;
  assign T175 = T176[4'h9:1'h0];
  assign T176 = T242 << T177;
  assign T177 = ~ T178;
  assign T178 = T319 ? 6'h3f : T179;
  assign T179 = T318 ? 6'h3e : T180;
  assign T180 = T317 ? 6'h3d : T181;
  assign T181 = T316 ? 6'h3c : T182;
  assign T182 = T315 ? 6'h3b : T183;
  assign T183 = T314 ? 6'h3a : T184;
  assign T184 = T313 ? 6'h39 : T185;
  assign T185 = T312 ? 6'h38 : T186;
  assign T186 = T311 ? 6'h37 : T187;
  assign T187 = T310 ? 6'h36 : T188;
  assign T188 = T309 ? 6'h35 : T189;
  assign T189 = T308 ? 6'h34 : T190;
  assign T190 = T307 ? 6'h33 : T191;
  assign T191 = T306 ? 6'h32 : T192;
  assign T192 = T305 ? 6'h31 : T193;
  assign T193 = T304 ? 6'h30 : T194;
  assign T194 = T303 ? 6'h2f : T195;
  assign T195 = T302 ? 6'h2e : T196;
  assign T196 = T301 ? 6'h2d : T197;
  assign T197 = T300 ? 6'h2c : T198;
  assign T198 = T299 ? 6'h2b : T199;
  assign T199 = T298 ? 6'h2a : T200;
  assign T200 = T297 ? 6'h29 : T201;
  assign T201 = T296 ? 6'h28 : T202;
  assign T202 = T295 ? 6'h27 : T203;
  assign T203 = T294 ? 6'h26 : T204;
  assign T204 = T293 ? 6'h25 : T205;
  assign T205 = T292 ? 6'h24 : T206;
  assign T206 = T291 ? 6'h23 : T207;
  assign T207 = T290 ? 6'h22 : T208;
  assign T208 = T289 ? 6'h21 : T209;
  assign T209 = T288 ? 6'h20 : T210;
  assign T210 = T287 ? 5'h1f : T211;
  assign T211 = T286 ? 5'h1e : T212;
  assign T212 = T285 ? 5'h1d : T213;
  assign T213 = T284 ? 5'h1c : T214;
  assign T214 = T283 ? 5'h1b : T215;
  assign T215 = T282 ? 5'h1a : T216;
  assign T216 = T281 ? 5'h19 : T217;
  assign T217 = T280 ? 5'h18 : T218;
  assign T218 = T279 ? 5'h17 : T219;
  assign T219 = T278 ? 5'h16 : T220;
  assign T220 = T277 ? 5'h15 : T221;
  assign T221 = T276 ? 5'h14 : T222;
  assign T222 = T275 ? 5'h13 : T223;
  assign T223 = T274 ? 5'h12 : T224;
  assign T224 = T273 ? 5'h11 : T225;
  assign T225 = T272 ? 5'h10 : T226;
  assign T226 = T271 ? 4'hf : T227;
  assign T227 = T270 ? 4'he : T228;
  assign T228 = T269 ? 4'hd : T229;
  assign T229 = T268 ? 4'hc : T230;
  assign T230 = T267 ? 4'hb : T231;
  assign T231 = T266 ? 4'ha : T232;
  assign T232 = T265 ? 4'h9 : T233;
  assign T233 = T264 ? 4'h8 : T234;
  assign T234 = T263 ? 3'h7 : T235;
  assign T235 = T262 ? 3'h6 : T236;
  assign T236 = T261 ? 3'h5 : T237;
  assign T237 = T260 ? 3'h4 : T238;
  assign T238 = T259 ? 2'h3 : T239;
  assign T239 = T258 ? 2'h2 : T240;
  assign T240 = T241[1'h1:1'h1];
  assign T241 = T242[6'h3f:1'h0];
  assign T242 = T255 ? T245 : T243;
  assign T243 = {32'h0, T244};
  assign T244 = T245[5'h1f:1'h0];
  assign T245 = T248 ? T247 : T246;
  assign T246 = R84[6'h3f:1'h0];
  assign T247 = 64'h0 - T246;
  assign T248 = T254 ? T253 : T249;
  assign T249 = T251 ? T250 : 1'h0;
  assign T250 = T246[6'h3f:6'h3f];
  assign T251 = T252 == 2'h3;
  assign T252 = R92 ^ 2'h1;
  assign T253 = T246[5'h1f:5'h1f];
  assign T254 = T252 == 2'h1;
  assign T255 = T257 | T256;
  assign T256 = T252 == 2'h2;
  assign T257 = T252 == 2'h3;
  assign T258 = T241[2'h2:2'h2];
  assign T259 = T241[2'h3:2'h3];
  assign T260 = T241[3'h4:3'h4];
  assign T261 = T241[3'h5:3'h5];
  assign T262 = T241[3'h6:3'h6];
  assign T263 = T241[3'h7:3'h7];
  assign T264 = T241[4'h8:4'h8];
  assign T265 = T241[4'h9:4'h9];
  assign T266 = T241[4'ha:4'ha];
  assign T267 = T241[4'hb:4'hb];
  assign T268 = T241[4'hc:4'hc];
  assign T269 = T241[4'hd:4'hd];
  assign T270 = T241[4'he:4'he];
  assign T271 = T241[4'hf:4'hf];
  assign T272 = T241[5'h10:5'h10];
  assign T273 = T241[5'h11:5'h11];
  assign T274 = T241[5'h12:5'h12];
  assign T275 = T241[5'h13:5'h13];
  assign T276 = T241[5'h14:5'h14];
  assign T277 = T241[5'h15:5'h15];
  assign T278 = T241[5'h16:5'h16];
  assign T279 = T241[5'h17:5'h17];
  assign T280 = T241[5'h18:5'h18];
  assign T281 = T241[5'h19:5'h19];
  assign T282 = T241[5'h1a:5'h1a];
  assign T283 = T241[5'h1b:5'h1b];
  assign T284 = T241[5'h1c:5'h1c];
  assign T285 = T241[5'h1d:5'h1d];
  assign T286 = T241[5'h1e:5'h1e];
  assign T287 = T241[5'h1f:5'h1f];
  assign T288 = T241[6'h20:6'h20];
  assign T289 = T241[6'h21:6'h21];
  assign T290 = T241[6'h22:6'h22];
  assign T291 = T241[6'h23:6'h23];
  assign T292 = T241[6'h24:6'h24];
  assign T293 = T241[6'h25:6'h25];
  assign T294 = T241[6'h26:6'h26];
  assign T295 = T241[6'h27:6'h27];
  assign T296 = T241[6'h28:6'h28];
  assign T297 = T241[6'h29:6'h29];
  assign T298 = T241[6'h2a:6'h2a];
  assign T299 = T241[6'h2b:6'h2b];
  assign T300 = T241[6'h2c:6'h2c];
  assign T301 = T241[6'h2d:6'h2d];
  assign T302 = T241[6'h2e:6'h2e];
  assign T303 = T241[6'h2f:6'h2f];
  assign T304 = T241[6'h30:6'h30];
  assign T305 = T241[6'h31:6'h31];
  assign T306 = T241[6'h32:6'h32];
  assign T307 = T241[6'h33:6'h33];
  assign T308 = T241[6'h34:6'h34];
  assign T309 = T241[6'h35:6'h35];
  assign T310 = T241[6'h36:6'h36];
  assign T311 = T241[6'h37:6'h37];
  assign T312 = T241[6'h38:6'h38];
  assign T313 = T241[6'h39:6'h39];
  assign T314 = T241[6'h3a:6'h3a];
  assign T315 = T241[6'h3b:6'h3b];
  assign T316 = T241[6'h3c:6'h3c];
  assign T317 = T241[6'h3d:6'h3d];
  assign T318 = T241[6'h3e:6'h3e];
  assign T319 = T241[6'h3f:6'h3f];
  assign T320 = T176[4'hb:4'ha];
  assign T321 = T165 & T322;
  assign T322 = R163 ^ 1'h1;
  assign T324 = reset ? 1'h0 : io_in_valid;
  assign T326 = reset ? 1'h0 : R323;
  assign io_out_bits_data = R327;
  assign T328 = R325 ? R329 : R327;
  assign T330 = R323 ? mux_data : R329;
  assign mux_data = T331;
  assign T331 = T321 ? T622 : T332;
  assign T332 = T162 ? T589 : T333;
  assign T333 = R163 ? T493 : T334;
  assign T334 = {T492, T335};
  assign T335 = {T470, T336};
  assign T336 = T468 ? T338 : T337;
  assign T337 = R84[6'h33:1'h0];
  assign T338 = T339[6'h3e:4'hb];
  assign T339 = T405 << T340;
  assign T340 = ~ T341;
  assign T341 = T467 ? 6'h3f : T342;
  assign T342 = T466 ? 6'h3e : T343;
  assign T343 = T465 ? 6'h3d : T344;
  assign T344 = T464 ? 6'h3c : T345;
  assign T345 = T463 ? 6'h3b : T346;
  assign T346 = T462 ? 6'h3a : T347;
  assign T347 = T461 ? 6'h39 : T348;
  assign T348 = T460 ? 6'h38 : T349;
  assign T349 = T459 ? 6'h37 : T350;
  assign T350 = T458 ? 6'h36 : T351;
  assign T351 = T457 ? 6'h35 : T352;
  assign T352 = T456 ? 6'h34 : T353;
  assign T353 = T455 ? 6'h33 : T354;
  assign T354 = T454 ? 6'h32 : T355;
  assign T355 = T453 ? 6'h31 : T356;
  assign T356 = T452 ? 6'h30 : T357;
  assign T357 = T451 ? 6'h2f : T358;
  assign T358 = T450 ? 6'h2e : T359;
  assign T359 = T449 ? 6'h2d : T360;
  assign T360 = T448 ? 6'h2c : T361;
  assign T361 = T447 ? 6'h2b : T362;
  assign T362 = T446 ? 6'h2a : T363;
  assign T363 = T445 ? 6'h29 : T364;
  assign T364 = T444 ? 6'h28 : T365;
  assign T365 = T443 ? 6'h27 : T366;
  assign T366 = T442 ? 6'h26 : T367;
  assign T367 = T441 ? 6'h25 : T368;
  assign T368 = T440 ? 6'h24 : T369;
  assign T369 = T439 ? 6'h23 : T370;
  assign T370 = T438 ? 6'h22 : T371;
  assign T371 = T437 ? 6'h21 : T372;
  assign T372 = T436 ? 6'h20 : T373;
  assign T373 = T435 ? 5'h1f : T374;
  assign T374 = T434 ? 5'h1e : T375;
  assign T375 = T433 ? 5'h1d : T376;
  assign T376 = T432 ? 5'h1c : T377;
  assign T377 = T431 ? 5'h1b : T378;
  assign T378 = T430 ? 5'h1a : T379;
  assign T379 = T429 ? 5'h19 : T380;
  assign T380 = T428 ? 5'h18 : T381;
  assign T381 = T427 ? 5'h17 : T382;
  assign T382 = T426 ? 5'h16 : T383;
  assign T383 = T425 ? 5'h15 : T384;
  assign T384 = T424 ? 5'h14 : T385;
  assign T385 = T423 ? 5'h13 : T386;
  assign T386 = T422 ? 5'h12 : T387;
  assign T387 = T421 ? 5'h11 : T388;
  assign T388 = T420 ? 5'h10 : T389;
  assign T389 = T419 ? 4'hf : T390;
  assign T390 = T418 ? 4'he : T391;
  assign T391 = T417 ? 4'hd : T392;
  assign T392 = T416 ? 4'hc : T393;
  assign T393 = T415 ? 4'hb : T394;
  assign T394 = T414 ? 4'ha : T395;
  assign T395 = T413 ? 4'h9 : T396;
  assign T396 = T412 ? 4'h8 : T397;
  assign T397 = T411 ? 3'h7 : T398;
  assign T398 = T410 ? 3'h6 : T399;
  assign T399 = T409 ? 3'h5 : T400;
  assign T400 = T408 ? 3'h4 : T401;
  assign T401 = T407 ? 2'h3 : T402;
  assign T402 = T406 ? 2'h2 : T403;
  assign T403 = T404[1'h1:1'h1];
  assign T404 = T405[6'h3f:1'h0];
  assign T405 = T337 << 4'hc;
  assign T406 = T404[2'h2:2'h2];
  assign T407 = T404[2'h3:2'h3];
  assign T408 = T404[3'h4:3'h4];
  assign T409 = T404[3'h5:3'h5];
  assign T410 = T404[3'h6:3'h6];
  assign T411 = T404[3'h7:3'h7];
  assign T412 = T404[4'h8:4'h8];
  assign T413 = T404[4'h9:4'h9];
  assign T414 = T404[4'ha:4'ha];
  assign T415 = T404[4'hb:4'hb];
  assign T416 = T404[4'hc:4'hc];
  assign T417 = T404[4'hd:4'hd];
  assign T418 = T404[4'he:4'he];
  assign T419 = T404[4'hf:4'hf];
  assign T420 = T404[5'h10:5'h10];
  assign T421 = T404[5'h11:5'h11];
  assign T422 = T404[5'h12:5'h12];
  assign T423 = T404[5'h13:5'h13];
  assign T424 = T404[5'h14:5'h14];
  assign T425 = T404[5'h15:5'h15];
  assign T426 = T404[5'h16:5'h16];
  assign T427 = T404[5'h17:5'h17];
  assign T428 = T404[5'h18:5'h18];
  assign T429 = T404[5'h19:5'h19];
  assign T430 = T404[5'h1a:5'h1a];
  assign T431 = T404[5'h1b:5'h1b];
  assign T432 = T404[5'h1c:5'h1c];
  assign T433 = T404[5'h1d:5'h1d];
  assign T434 = T404[5'h1e:5'h1e];
  assign T435 = T404[5'h1f:5'h1f];
  assign T436 = T404[6'h20:6'h20];
  assign T437 = T404[6'h21:6'h21];
  assign T438 = T404[6'h22:6'h22];
  assign T439 = T404[6'h23:6'h23];
  assign T440 = T404[6'h24:6'h24];
  assign T441 = T404[6'h25:6'h25];
  assign T442 = T404[6'h26:6'h26];
  assign T443 = T404[6'h27:6'h27];
  assign T444 = T404[6'h28:6'h28];
  assign T445 = T404[6'h29:6'h29];
  assign T446 = T404[6'h2a:6'h2a];
  assign T447 = T404[6'h2b:6'h2b];
  assign T448 = T404[6'h2c:6'h2c];
  assign T449 = T404[6'h2d:6'h2d];
  assign T450 = T404[6'h2e:6'h2e];
  assign T451 = T404[6'h2f:6'h2f];
  assign T452 = T404[6'h30:6'h30];
  assign T453 = T404[6'h31:6'h31];
  assign T454 = T404[6'h32:6'h32];
  assign T455 = T404[6'h33:6'h33];
  assign T456 = T404[6'h34:6'h34];
  assign T457 = T404[6'h35:6'h35];
  assign T458 = T404[6'h36:6'h36];
  assign T459 = T404[6'h37:6'h37];
  assign T460 = T404[6'h38:6'h38];
  assign T461 = T404[6'h39:6'h39];
  assign T462 = T404[6'h3a:6'h3a];
  assign T463 = T404[6'h3b:6'h3b];
  assign T464 = T404[6'h3c:6'h3c];
  assign T465 = T404[6'h3d:6'h3d];
  assign T466 = T404[6'h3e:6'h3e];
  assign T467 = T404[6'h3f:6'h3f];
  assign T468 = T469 == 11'h0;
  assign T469 = R84[6'h3e:6'h34];
  assign T470 = T478 | T471;
  assign T471 = {2'h0, T472};
  assign T472 = T473 << 4'h9;
  assign T473 = T476 & T474;
  assign T474 = T475 ^ 1'h1;
  assign T475 = T337 == 52'h0;
  assign T476 = T477 == 2'h3;
  assign T477 = T478[4'hb:4'ha];
  assign T478 = T487 + T479;
  assign T479 = {1'h0, T480};
  assign T480 = T486 ? 11'h0 : T481;
  assign T481 = 11'h400 | T482;
  assign T482 = {9'h0, T483};
  assign T483 = T484 ? 2'h2 : 2'h1;
  assign T484 = T468 & T485;
  assign T485 = T475 ^ 1'h1;
  assign T486 = T468 & T475;
  assign T487 = T468 ? T489 : T488;
  assign T488 = {1'h0, T469};
  assign T489 = T475 ? 12'h0 : T490;
  assign T490 = {6'h3f, T491};
  assign T491 = ~ T340;
  assign T492 = R84[6'h3f:6'h3f];
  assign T493 = {32'hffffffff, T494};
  assign T494 = {T588, T495};
  assign T495 = {T566, T496};
  assign T496 = T564 ? T498 : T497;
  assign T497 = R84[5'h16:1'h0];
  assign T498 = T499[5'h1e:4'h8];
  assign T499 = T533 << T500;
  assign T500 = ~ T501;
  assign T501 = T563 ? 5'h1f : T502;
  assign T502 = T562 ? 5'h1e : T503;
  assign T503 = T561 ? 5'h1d : T504;
  assign T504 = T560 ? 5'h1c : T505;
  assign T505 = T559 ? 5'h1b : T506;
  assign T506 = T558 ? 5'h1a : T507;
  assign T507 = T557 ? 5'h19 : T508;
  assign T508 = T556 ? 5'h18 : T509;
  assign T509 = T555 ? 5'h17 : T510;
  assign T510 = T554 ? 5'h16 : T511;
  assign T511 = T553 ? 5'h15 : T512;
  assign T512 = T552 ? 5'h14 : T513;
  assign T513 = T551 ? 5'h13 : T514;
  assign T514 = T550 ? 5'h12 : T515;
  assign T515 = T549 ? 5'h11 : T516;
  assign T516 = T548 ? 5'h10 : T517;
  assign T517 = T547 ? 4'hf : T518;
  assign T518 = T546 ? 4'he : T519;
  assign T519 = T545 ? 4'hd : T520;
  assign T520 = T544 ? 4'hc : T521;
  assign T521 = T543 ? 4'hb : T522;
  assign T522 = T542 ? 4'ha : T523;
  assign T523 = T541 ? 4'h9 : T524;
  assign T524 = T540 ? 4'h8 : T525;
  assign T525 = T539 ? 3'h7 : T526;
  assign T526 = T538 ? 3'h6 : T527;
  assign T527 = T537 ? 3'h5 : T528;
  assign T528 = T536 ? 3'h4 : T529;
  assign T529 = T535 ? 2'h3 : T530;
  assign T530 = T534 ? 2'h2 : T531;
  assign T531 = T532[1'h1:1'h1];
  assign T532 = T533[5'h1f:1'h0];
  assign T533 = T497 << 4'h9;
  assign T534 = T532[2'h2:2'h2];
  assign T535 = T532[2'h3:2'h3];
  assign T536 = T532[3'h4:3'h4];
  assign T537 = T532[3'h5:3'h5];
  assign T538 = T532[3'h6:3'h6];
  assign T539 = T532[3'h7:3'h7];
  assign T540 = T532[4'h8:4'h8];
  assign T541 = T532[4'h9:4'h9];
  assign T542 = T532[4'ha:4'ha];
  assign T543 = T532[4'hb:4'hb];
  assign T544 = T532[4'hc:4'hc];
  assign T545 = T532[4'hd:4'hd];
  assign T546 = T532[4'he:4'he];
  assign T547 = T532[4'hf:4'hf];
  assign T548 = T532[5'h10:5'h10];
  assign T549 = T532[5'h11:5'h11];
  assign T550 = T532[5'h12:5'h12];
  assign T551 = T532[5'h13:5'h13];
  assign T552 = T532[5'h14:5'h14];
  assign T553 = T532[5'h15:5'h15];
  assign T554 = T532[5'h16:5'h16];
  assign T555 = T532[5'h17:5'h17];
  assign T556 = T532[5'h18:5'h18];
  assign T557 = T532[5'h19:5'h19];
  assign T558 = T532[5'h1a:5'h1a];
  assign T559 = T532[5'h1b:5'h1b];
  assign T560 = T532[5'h1c:5'h1c];
  assign T561 = T532[5'h1d:5'h1d];
  assign T562 = T532[5'h1e:5'h1e];
  assign T563 = T532[5'h1f:5'h1f];
  assign T564 = T565 == 8'h0;
  assign T565 = R84[5'h1e:5'h17];
  assign T566 = T574 | T567;
  assign T567 = {2'h0, T568};
  assign T568 = T569 << 3'h6;
  assign T569 = T572 & T570;
  assign T570 = T571 ^ 1'h1;
  assign T571 = T497 == 23'h0;
  assign T572 = T573 == 2'h3;
  assign T573 = T574[4'h8:3'h7];
  assign T574 = T583 + T575;
  assign T575 = {1'h0, T576};
  assign T576 = T582 ? 8'h0 : T577;
  assign T577 = 8'h80 | T578;
  assign T578 = {6'h0, T579};
  assign T579 = T580 ? 2'h2 : 2'h1;
  assign T580 = T564 & T581;
  assign T581 = T571 ^ 1'h1;
  assign T582 = T564 & T571;
  assign T583 = T564 ? T585 : T584;
  assign T584 = {1'h0, T565};
  assign T585 = T571 ? 9'h0 : T586;
  assign T586 = {4'hf, T587};
  assign T587 = ~ T500;
  assign T588 = R84[5'h1f:5'h1f];
  assign T589 = {32'hffffffff, T590};
  assign T590 = {T87, T591};
  assign T591 = {T613, T592};
  assign T592 = T593[5'h16:1'h0];
  assign T593 = T597 ? T596 : T594;
  assign T594 = {1'h0, T595};
  assign T595 = T13[6'h3f:6'h28];
  assign T596 = T594 + 25'h1;
  assign T597 = T612 ? T607 : T598;
  assign T598 = T606 ? T605 : T599;
  assign T599 = T602 ? T600 : 1'h0;
  assign T600 = T601 & T8;
  assign T601 = T87 ^ 1'h1;
  assign T602 = R603 == 3'h3;
  assign T604 = io_in_valid ? io_in_bits_rm : R603;
  assign T605 = T87 & T8;
  assign T606 = R603 == 3'h2;
  assign T607 = T610 | T608;
  assign T608 = T609 == 2'h3;
  assign T609 = T10[1'h1:1'h0];
  assign T610 = T611 == 2'h3;
  assign T611 = T10[2'h2:1'h1];
  assign T612 = R603 == 3'h0;
  assign T613 = {T621, T614};
  assign T614 = T615[3'h7:1'h0];
  assign T615 = T618 + T616;
  assign T616 = {7'h0, T617};
  assign T617 = T593[5'h18:5'h18];
  assign T618 = {1'h0, T619};
  assign T619 = {1'h0, T620};
  assign T620 = ~ T14;
  assign T621 = T13[6'h3f:6'h3f];
  assign T622 = {T248, T623};
  assign T623 = {T643, T624};
  assign T624 = T625[6'h33:1'h0];
  assign T625 = T629 ? T628 : T626;
  assign T626 = {1'h0, T627};
  assign T627 = T176[6'h3f:4'hb];
  assign T628 = T626 + 54'h1;
  assign T629 = T642 ? T637 : T630;
  assign T630 = T636 ? T635 : T631;
  assign T631 = T634 ? T632 : 1'h0;
  assign T632 = T633 & T171;
  assign T633 = T248 ^ 1'h1;
  assign T634 = R603 == 3'h3;
  assign T635 = T248 & T171;
  assign T636 = R603 == 3'h2;
  assign T637 = T640 | T638;
  assign T638 = T639 == 2'h3;
  assign T639 = T173[1'h1:1'h0];
  assign T640 = T641 == 2'h3;
  assign T641 = T173[2'h2:1'h1];
  assign T642 = R603 == 3'h0;
  assign T643 = {T651, T644};
  assign T644 = T645[4'ha:1'h0];
  assign T645 = T648 + T646;
  assign T646 = {10'h0, T647};
  assign T647 = T625[6'h35:6'h35];
  assign T648 = {1'h0, T649};
  assign T649 = {4'h0, T650};
  assign T650 = ~ T177;
  assign T651 = T176[6'h3f:6'h3f];
  assign io_out_valid = R652;
  assign T653 = reset ? 1'h0 : R325;

  always @(posedge clk) begin
    if(R325) begin
      R0 <= R2;
    end
    if(R323) begin
      R2 <= mux_exc;
    end
    if(io_in_valid) begin
      R84 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R92 <= io_in_bits_typ;
    end
    if(io_in_valid) begin
      R163 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R167 <= io_in_bits_cmd;
    end
    if(reset) begin
      R323 <= 1'h0;
    end else begin
      R323 <= io_in_valid;
    end
    if(reset) begin
      R325 <= 1'h0;
    end else begin
      R325 <= R323;
    end
    if(R325) begin
      R327 <= R329;
    end
    if(R323) begin
      R329 <= mux_data;
    end
    if(io_in_valid) begin
      R603 <= io_in_bits_rm;
    end
    if(reset) begin
      R652 <= 1'h0;
    end else begin
      R652 <= R325;
    end
  end
endmodule

module FPToFP(input clk, input reset,
    input  io_in_valid,
    input [4:0] io_in_bits_cmd,
    input  io_in_bits_ldst,
    input  io_in_bits_wen,
    input  io_in_bits_ren1,
    input  io_in_bits_ren2,
    input  io_in_bits_ren3,
    input  io_in_bits_swap23,
    input  io_in_bits_single,
    input  io_in_bits_fromint,
    input  io_in_bits_toint,
    input  io_in_bits_fastpipe,
    input  io_in_bits_fma,
    input  io_in_bits_round,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output[64:0] io_out_bits_data,
    output[4:0] io_out_bits_exc,
    input  io_lt
);

  reg [4:0] R0;
  wire[4:0] T1;
  wire[4:0] mux_exc;
  wire[4:0] T2;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] minmax_exc;
  wire T5;
  wire issnan2;
  wire T6;
  wire T7;
  wire T8;
  reg [64:0] R9;
  wire[64:0] T10;
  wire T11;
  reg  R12;
  wire T13;
  wire isnan2;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire issnan1;
  wire T18;
  wire T19;
  wire T20;
  reg [64:0] R21;
  wire[64:0] T22;
  wire T23;
  wire isnan1;
  wire T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire[4:0] T29;
  reg [4:0] R30;
  wire[4:0] T31;
  wire[4:0] T32;
  wire[2:0] T33;
  wire[1:0] T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  wire[2:0] T41;
  wire T42;
  wire T43;
  wire T44;
  wire[11:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire[1:0] T53;
  wire[2:0] T54;
  wire T55;
  wire T56;
  wire[27:0] T57;
  wire[51:0] T58;
  wire T59;
  wire[23:0] T60;
  wire[48:0] T61;
  wire[4:0] T62;
  wire[11:0] T63;
  wire[11:0] T64;
  wire T65;
  wire T66;
  wire T67;
  wire[48:0] T68;
  wire[47:0] T69;
  wire[23:0] T70;
  wire[1:0] T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire[24:0] T77;
  wire[24:0] T78;
  wire[24:0] T79;
  wire[24:0] T80;
  wire[55:0] T81;
  wire[4:0] T82;
  wire[24:0] T83;
  wire[22:0] T84;
  wire[24:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  reg [2:0] R93;
  wire[2:0] T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire[1:0] T99;
  wire T100;
  wire[1:0] T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire[4:0] T111;
  wire[4:0] T112;
  wire T113;
  wire T114;
  wire T115;
  wire[22:0] T116;
  wire T117;
  wire[2:0] T118;
  wire T119;
  wire T120;
  reg  R121;
  wire T122;
  reg [64:0] R123;
  wire[64:0] T124;
  wire[64:0] mux_data;
  wire[64:0] T125;
  wire[64:0] T126;
  wire[64:0] T127;
  wire[64:0] fsgnj;
  wire[32:0] T128;
  wire[31:0] T129;
  wire sign_s;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire[31:0] T139;
  wire[30:0] T140;
  wire sign_d;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire isLHS;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire[64:0] T156;
  wire[32:0] T157;
  wire[31:0] T158;
  wire[22:0] T159;
  wire[22:0] T160;
  wire[22:0] T161;
  wire[22:0] T162;
  wire[22:0] T163;
  wire[22:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire[22:0] T174;
  wire[22:0] T175;
  wire[8:0] T176;
  wire[8:0] T177;
  wire[8:0] T178;
  wire[8:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire[8:0] T182;
  wire T183;
  wire[8:0] T184;
  wire[6:0] T185;
  wire[8:0] T186;
  wire[8:0] T187;
  wire[64:0] T188;
  wire[63:0] T189;
  wire[51:0] T190;
  wire[51:0] T191;
  wire[51:0] T192;
  wire[51:0] T193;
  wire[11:0] T194;
  wire[11:0] T195;
  wire[11:0] T196;
  wire[11:0] T197;
  wire T198;
  wire[11:0] T199;
  wire[7:0] T200;
  wire T201;
  wire[11:0] T202;
  wire[10:0] T203;
  wire T204;
  wire[11:0] T205;
  wire T206;
  wire T207;
  reg  R208;
  wire T209;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R9 = {3{$random}};
    R12 = {1{$random}};
    R21 = {3{$random}};
    R30 = {1{$random}};
    R93 = {1{$random}};
    R121 = {1{$random}};
    R123 = {3{$random}};
    R208 = {1{$random}};
  end
`endif

  assign io_out_bits_exc = R0;
  assign T1 = R121 ? mux_exc : R0;
  assign mux_exc = T2;
  assign T2 = T119 ? T112 : T3;
  assign T3 = T109 ? T32 : T4;
  assign T4 = T28 ? 5'h0 : minmax_exc;
  assign minmax_exc = {T5, 4'h0};
  assign T5 = issnan1 | issnan2;
  assign issnan2 = isnan2 & T6;
  assign T6 = ~ T7;
  assign T7 = R12 ? T11 : T8;
  assign T8 = R9[6'h33:6'h33];
  assign T10 = io_in_valid ? io_in_bits_in2 : R9;
  assign T11 = R9[5'h16:5'h16];
  assign T13 = io_in_valid ? io_in_bits_single : R12;
  assign isnan2 = R12 ? T16 : T14;
  assign T14 = T15 == 3'h7;
  assign T15 = R9[6'h3f:6'h3d];
  assign T16 = T17 == 3'h7;
  assign T17 = R9[5'h1f:5'h1d];
  assign issnan1 = isnan1 & T18;
  assign T18 = ~ T19;
  assign T19 = R12 ? T23 : T20;
  assign T20 = R21[6'h33:6'h33];
  assign T22 = io_in_valid ? io_in_bits_in1 : R21;
  assign T23 = R21[5'h16:5'h16];
  assign isnan1 = R12 ? T26 : T24;
  assign T24 = T25 == 3'h7;
  assign T25 = R21[6'h3f:6'h3d];
  assign T26 = T27 == 3'h7;
  assign T27 = R21[5'h1f:5'h1d];
  assign T28 = T29 == 5'h4;
  assign T29 = R30 & 5'h5;
  assign T31 = io_in_valid ? io_in_bits_cmd : R30;
  assign T32 = {T104, T33};
  assign T33 = {T74, T34};
  assign T34 = {T72, T35};
  assign T35 = T46 | T36;
  assign T36 = T44 & T37;
  assign T37 = T38 ^ 1'h1;
  assign T38 = T42 | T39;
  assign T39 = T40 == 2'h3;
  assign T40 = T41[2'h2:1'h1];
  assign T41 = R21[6'h3f:6'h3d];
  assign T42 = T43 ^ 1'h1;
  assign T43 = T41 != 3'h0;
  assign T44 = T45 < 12'h76a;
  assign T45 = R21[6'h3f:6'h34];
  assign T46 = T50 | T47;
  assign T47 = T49 & T48;
  assign T48 = T38 ^ 1'h1;
  assign T49 = 12'h87f < T45;
  assign T50 = T52 & T51;
  assign T51 = T38 ^ 1'h1;
  assign T52 = T53 != 2'h0;
  assign T53 = T54[1'h1:1'h0];
  assign T54 = {T71, T55};
  assign T55 = T59 | T56;
  assign T56 = T57 != 28'h0;
  assign T57 = T58[5'h1b:1'h0];
  assign T58 = R21[6'h33:1'h0];
  assign T59 = T60 != 24'h0;
  assign T60 = T61[5'h17:1'h0];
  assign T61 = T68 >> T62;
  assign T62 = T63[3'h4:1'h0];
  assign T63 = T65 ? T64 : 12'h0;
  assign T64 = 12'h782 - T45;
  assign T65 = T67 & T66;
  assign T66 = T45 <= 12'h781;
  assign T67 = 12'h76a <= T45;
  assign T68 = {1'h1, T69};
  assign T69 = {T70, 24'h0};
  assign T70 = T58[6'h33:5'h1c];
  assign T71 = T61[5'h19:5'h18];
  assign T72 = T36 | T73;
  assign T73 = T65 & T50;
  assign T74 = T47 | T75;
  assign T75 = T103 & T76;
  assign T76 = T77[5'h18:5'h18];
  assign T77 = T86 ? T85 : T78;
  assign T78 = T83 | T79;
  assign T79 = ~ T80;
  assign T80 = T81[5'h18:1'h0];
  assign T81 = 25'h1ffffff << T82;
  assign T82 = T62;
  assign T83 = {2'h1, T84};
  assign T84 = T58[6'h33:5'h1d];
  assign T85 = T78 + 25'h1;
  assign T86 = T102 ? T97 : T87;
  assign T87 = T96 ? T95 : T88;
  assign T88 = T92 ? T89 : 1'h0;
  assign T89 = T90 & T50;
  assign T90 = T91 ^ 1'h1;
  assign T91 = R21[7'h40:7'h40];
  assign T92 = R93 == 3'h3;
  assign T94 = io_in_valid ? io_in_bits_rm : R93;
  assign T95 = T91 & T50;
  assign T96 = R93 == 3'h2;
  assign T97 = T100 | T98;
  assign T98 = T99 == 2'h3;
  assign T99 = T54[2'h2:1'h1];
  assign T100 = T101 == 2'h3;
  assign T101 = T54[1'h1:1'h0];
  assign T102 = R93 == 3'h0;
  assign T103 = T45 == 12'h87f;
  assign T104 = {T105, 1'h0};
  assign T105 = T108 & T106;
  assign T106 = T107 ^ 1'h1;
  assign T107 = T58[6'h33:6'h33];
  assign T108 = T41 == 3'h7;
  assign T109 = T110 & R12;
  assign T110 = T111 == 5'h0;
  assign T111 = R30 & 5'h4;
  assign T112 = T113 << 3'h4;
  assign T113 = T117 & T114;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116[5'h16:5'h16];
  assign T116 = R21[5'h16:1'h0];
  assign T117 = T118 == 3'h7;
  assign T118 = R21[5'h1f:5'h1d];
  assign T119 = T110 & T120;
  assign T120 = R12 ^ 1'h1;
  assign T122 = reset ? 1'h0 : io_in_valid;
  assign io_out_bits_data = R123;
  assign T124 = R121 ? mux_data : R123;
  assign mux_data = T125;
  assign T125 = T119 ? T188 : T126;
  assign T126 = T109 ? T156 : T127;
  assign T127 = T151 ? fsgnj : R9;
  assign fsgnj = {T139, T128};
  assign T128 = {sign_s, T129};
  assign T129 = R21[5'h1f:1'h0];
  assign sign_s = T133 ^ T130;
  assign T130 = T132 & T131;
  assign T131 = R9[6'h20:6'h20];
  assign T132 = R12 & T28;
  assign T133 = T136 ? T135 : T134;
  assign T134 = R93[1'h0:1'h0];
  assign T135 = R21[6'h20:6'h20];
  assign T136 = T138 | T137;
  assign T137 = T132 ^ 1'h1;
  assign T138 = R93[1'h1:1'h1];
  assign T139 = {sign_d, T140};
  assign T140 = R21[6'h3f:6'h21];
  assign sign_d = T145 ^ T141;
  assign T141 = T143 & T142;
  assign T142 = R9[7'h40:7'h40];
  assign T143 = T144 & T28;
  assign T144 = R12 ^ 1'h1;
  assign T145 = T148 ? T147 : T146;
  assign T146 = R93[1'h0:1'h0];
  assign T147 = R21[7'h40:7'h40];
  assign T148 = T150 | T149;
  assign T149 = T143 ^ 1'h1;
  assign T150 = R93[1'h1:1'h1];
  assign T151 = T28 | isLHS;
  assign isLHS = isnan2 | T152;
  assign T152 = T154 & T153;
  assign T153 = isnan1 ^ 1'h1;
  assign T154 = T155 != io_lt;
  assign T155 = R93[1'h0:1'h0];
  assign T156 = {32'hffffffff, T157};
  assign T157 = {T91, T158};
  assign T158 = {T176, T159};
  assign T159 = T38 ? T174 : T160;
  assign T160 = T47 ? T163 : T161;
  assign T161 = T36 ? 23'h0 : T162;
  assign T162 = T77[5'h16:1'h0];
  assign T163 = 23'h0 - T164;
  assign T164 = {22'h0, T165};
  assign T165 = T166 ^ 1'h1;
  assign T166 = T168 | T167;
  assign T167 = R93 == 3'h0;
  assign T168 = T172 | T169;
  assign T169 = T171 & T170;
  assign T170 = T91 ^ 1'h1;
  assign T171 = R93 == 3'h3;
  assign T172 = T173 & T91;
  assign T173 = R93 == 3'h2;
  assign T174 = 23'h0 - T175;
  assign T175 = {22'h0, T108};
  assign T176 = T38 ? T187 : T177;
  assign T177 = T47 ? T186 : T178;
  assign T178 = T36 ? T184 : T179;
  assign T179 = T183 ? T182 : T180;
  assign T180 = T181 + 9'h100;
  assign T181 = T45[4'h8:1'h0];
  assign T182 = T180 + 9'h1;
  assign T183 = T77[5'h18:5'h18];
  assign T184 = {2'h0, T185};
  assign T185 = T168 ? 7'h6b : 7'h0;
  assign T186 = T166 ? 9'h180 : 9'h17f;
  assign T187 = T41 << 3'h6;
  assign T188 = {T207, T189};
  assign T189 = {T194, T190};
  assign T190 = T192 | T191;
  assign T191 = T116 << 5'h1d;
  assign T192 = 52'h0 - T193;
  assign T193 = {51'h0, T117};
  assign T194 = T206 ? T205 : T195;
  assign T195 = T204 ? T202 : T196;
  assign T196 = T201 ? T199 : T197;
  assign T197 = T198 ? 12'hc00 : 12'he00;
  assign T198 = T118 < 3'h7;
  assign T199 = {4'h8, T200};
  assign T200 = R21[5'h1e:5'h17];
  assign T201 = T118 < 3'h6;
  assign T202 = {1'h0, T203};
  assign T203 = {3'h7, T200};
  assign T204 = T118 < 3'h4;
  assign T205 = {4'h0, T200};
  assign T206 = T118 < 3'h1;
  assign T207 = R21[6'h20:6'h20];
  assign io_out_valid = R208;
  assign T209 = reset ? 1'h0 : R121;

  always @(posedge clk) begin
    if(R121) begin
      R0 <= mux_exc;
    end
    if(io_in_valid) begin
      R9 <= io_in_bits_in2;
    end
    if(io_in_valid) begin
      R12 <= io_in_bits_single;
    end
    if(io_in_valid) begin
      R21 <= io_in_bits_in1;
    end
    if(io_in_valid) begin
      R30 <= io_in_bits_cmd;
    end
    if(io_in_valid) begin
      R93 <= io_in_bits_rm;
    end
    if(reset) begin
      R121 <= 1'h0;
    end else begin
      R121 <= io_in_valid;
    end
    if(R121) begin
      R123 <= mux_data;
    end
    if(reset) begin
      R208 <= 1'h0;
    end else begin
      R208 <= R121;
    end
  end
endmodule

module FPU(input clk, input reset,
    input  io_ctrl_valid,
    output io_ctrl_fcsr_rdy,
    output io_ctrl_nack_mem,
    output io_ctrl_illegal_rm,
    input  io_ctrl_killx,
    input  io_ctrl_killm,
    output[4:0] io_ctrl_dec_cmd,
    output io_ctrl_dec_ldst,
    output io_ctrl_dec_wen,
    output io_ctrl_dec_ren1,
    output io_ctrl_dec_ren2,
    output io_ctrl_dec_ren3,
    output io_ctrl_dec_swap23,
    output io_ctrl_dec_single,
    output io_ctrl_dec_fromint,
    output io_ctrl_dec_toint,
    output io_ctrl_dec_fastpipe,
    output io_ctrl_dec_fma,
    output io_ctrl_dec_round,
    output io_ctrl_sboard_set,
    output io_ctrl_sboard_clr,
    output[4:0] io_ctrl_sboard_clra,
    input [31:0] io_dpath_inst,
    input [63:0] io_dpath_fromint_data,
    input [2:0] io_dpath_fcsr_rm,
    output io_dpath_fcsr_flags_valid,
    output[4:0] io_dpath_fcsr_flags_bits,
    output[63:0] io_dpath_store_data,
    output[63:0] io_dpath_toint_data,
    input  io_dpath_dmem_resp_val,
    input [2:0] io_dpath_dmem_resp_type,
    input [4:0] io_dpath_dmem_resp_tag,
    input [63:0] io_dpath_dmem_resp_data
);

  wire fpiu_io_out_bits_lt;
  wire[64:0] req_in3;
  wire[64:0] T0;
  reg [64:0] regfile [31:0];
  wire[64:0] T1;
  wire[64:0] T2;
  wire[96:0] T3;
  wire[96:0] T4;
  wire[64:0] T5;
  wire[64:0] fpmu_io_out_bits_data;
  wire[64:0] ifpu_io_out_bits_data;
  wire T6;
  wire[1:0] T7;
  wire[1:0] wsrc;
  reg [6:0] winfo_0;
  wire[6:0] T8;
  wire[6:0] T9;
  reg [6:0] winfo_1;
  wire[6:0] T10;
  wire[6:0] mem_winfo;
  wire[4:0] T11;
  reg [31:0] mem_reg_inst;
  wire[31:0] T12;
  reg [31:0] ex_reg_inst;
  wire[31:0] T13;
  reg  ex_reg_valid;
  wire T14;
  wire[1:0] T15;
  wire[1:0] T16;
  wire T17;
  wire T18;
  reg  mem_ctrl_single;
  wire T19;
  reg  ex_ctrl_single;
  wire T20;
  wire fp_decoder_io_sigs_single;
  reg  mem_ctrl_fma;
  wire T21;
  reg  ex_ctrl_fma;
  wire T22;
  wire fp_decoder_io_sigs_fma;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire[1:0] T26;
  wire T27;
  reg  mem_ctrl_fromint;
  wire T28;
  reg  ex_ctrl_fromint;
  wire T29;
  wire fp_decoder_io_sigs_fromint;
  wire T30;
  wire T31;
  wire T32;
  wire[1:0] memLatencyMask;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  reg  mem_ctrl_fastpipe;
  wire T42;
  reg  ex_ctrl_fastpipe;
  wire T43;
  wire fp_decoder_io_sigs_fastpipe;
  wire T44;
  reg  write_port_busy;
  wire T45;
  wire T46;
  wire T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire[3:0] T50;
  wire T51;
  wire T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire[2:0] T55;
  wire T56;
  wire[3:0] T57;
  wire[3:0] T58;
  wire[3:0] T59;
  wire[2:0] T60;
  wire[3:0] T61;
  reg [1:0] wen;
  wire[1:0] T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire killm;
  wire mem_wen;
  wire T71;
  wire T72;
  reg  mem_reg_valid;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire[2:0] T78;
  wire[2:0] T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire[2:0] T87;
  wire[2:0] T88;
  wire[2:0] T89;
  wire[1:0] T90;
  wire[2:0] T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire[96:0] T97;
  wire[96:0] T98;
  wire[64:0] sfma_io_out_bits_data;
  wire[96:0] T99;
  wire[64:0] dfma_io_out_bits_data;
  wire T100;
  wire T101;
  wire T102;
  wire[4:0] T103;
  wire[4:0] waddr;
  wire[4:0] T104;
  wire[64:0] T105;
  wire[64:0] load_wb_data_recoded;
  wire[64:0] rec_d;
  wire[63:0] T106;
  wire[51:0] T107;
  wire[51:0] T108;
  reg [63:0] load_wb_data;
  wire[63:0] T109;
  wire[51:0] T110;
  wire[126:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] T114;
  wire[5:0] T115;
  wire[5:0] T116;
  wire[5:0] T117;
  wire[5:0] T118;
  wire[5:0] T119;
  wire[5:0] T120;
  wire[5:0] T121;
  wire[5:0] T122;
  wire[5:0] T123;
  wire[5:0] T124;
  wire[5:0] T125;
  wire[5:0] T126;
  wire[5:0] T127;
  wire[5:0] T128;
  wire[5:0] T129;
  wire[5:0] T130;
  wire[5:0] T131;
  wire[5:0] T132;
  wire[5:0] T133;
  wire[5:0] T134;
  wire[5:0] T135;
  wire[5:0] T136;
  wire[5:0] T137;
  wire[5:0] T138;
  wire[5:0] T139;
  wire[5:0] T140;
  wire[5:0] T141;
  wire[5:0] T142;
  wire[5:0] T143;
  wire[5:0] T144;
  wire[4:0] T145;
  wire[4:0] T146;
  wire[4:0] T147;
  wire[4:0] T148;
  wire[4:0] T149;
  wire[4:0] T150;
  wire[4:0] T151;
  wire[4:0] T152;
  wire[4:0] T153;
  wire[4:0] T154;
  wire[4:0] T155;
  wire[4:0] T156;
  wire[4:0] T157;
  wire[4:0] T158;
  wire[4:0] T159;
  wire[4:0] T160;
  wire[3:0] T161;
  wire[3:0] T162;
  wire[3:0] T163;
  wire[3:0] T164;
  wire[3:0] T165;
  wire[3:0] T166;
  wire[3:0] T167;
  wire[3:0] T168;
  wire[2:0] T169;
  wire[2:0] T170;
  wire[2:0] T171;
  wire[2:0] T172;
  wire[1:0] T173;
  wire[1:0] T174;
  wire T175;
  wire[63:0] T176;
  wire[63:0] T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire[10:0] T241;
  wire[11:0] T242;
  wire[11:0] T243;
  wire[9:0] T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[11:0] T250;
  wire[11:0] T251;
  wire[10:0] T252;
  wire[10:0] T253;
  wire[10:0] T254;
  wire[1:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[11:0] T259;
  wire[11:0] T260;
  wire[11:0] T261;
  wire[11:0] T262;
  wire[5:0] T263;
  wire T264;
  wire[64:0] T265;
  wire[32:0] rec_s;
  wire[31:0] T266;
  wire[22:0] T267;
  wire[22:0] T268;
  wire[22:0] T269;
  wire[62:0] T270;
  wire[4:0] T271;
  wire[4:0] T272;
  wire[4:0] T273;
  wire[4:0] T274;
  wire[4:0] T275;
  wire[4:0] T276;
  wire[4:0] T277;
  wire[4:0] T278;
  wire[4:0] T279;
  wire[4:0] T280;
  wire[4:0] T281;
  wire[4:0] T282;
  wire[4:0] T283;
  wire[4:0] T284;
  wire[4:0] T285;
  wire[4:0] T286;
  wire[4:0] T287;
  wire[3:0] T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[3:0] T294;
  wire[3:0] T295;
  wire[2:0] T296;
  wire[2:0] T297;
  wire[2:0] T298;
  wire[2:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire[7:0] T336;
  wire[8:0] T337;
  wire[8:0] T338;
  wire[6:0] T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[1:0] T344;
  wire[8:0] T345;
  wire[8:0] T346;
  wire[7:0] T347;
  wire[7:0] T348;
  wire[7:0] T349;
  wire[1:0] T350;
  wire T351;
  wire T352;
  wire T353;
  wire[8:0] T354;
  wire[8:0] T355;
  wire[8:0] T356;
  wire[8:0] T357;
  wire[4:0] T358;
  wire T359;
  reg  load_wb_single;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  reg  load_wb;
  reg [4:0] load_wb_tag;
  wire[4:0] T364;
  reg [4:0] ex_ra3;
  wire[4:0] T365;
  wire[4:0] T366;
  wire[4:0] T367;
  wire T368;
  wire fp_decoder_io_sigs_ren3;
  wire[4:0] T369;
  wire T370;
  wire T371;
  wire fp_decoder_io_sigs_swap23;
  wire T372;
  wire fp_decoder_io_sigs_ldst;
  wire T373;
  wire fp_decoder_io_sigs_ren2;
  wire[64:0] req_in2;
  wire[64:0] T374;
  reg [4:0] ex_ra2;
  wire[4:0] T375;
  wire[4:0] T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire[64:0] req_in1;
  wire[64:0] T381;
  reg [4:0] ex_ra1;
  wire[4:0] T382;
  wire[4:0] T383;
  wire[4:0] T384;
  wire T385;
  wire fp_decoder_io_sigs_ren1;
  wire[4:0] T386;
  wire T387;
  wire[1:0] req_typ;
  wire[1:0] T388;
  wire[2:0] req_rm;
  wire[2:0] ex_rm;
  wire[2:0] T389;
  wire T390;
  wire[2:0] T391;
  wire req_round;
  reg  ex_ctrl_round;
  wire T392;
  wire fp_decoder_io_sigs_round;
  wire req_fma;
  wire req_fastpipe;
  wire req_toint;
  reg  ex_ctrl_toint;
  wire T393;
  wire fp_decoder_io_sigs_toint;
  wire req_fromint;
  wire req_single;
  wire req_swap23;
  reg  ex_ctrl_swap23;
  wire T394;
  wire req_ren3;
  reg  ex_ctrl_ren3;
  wire T395;
  wire req_ren2;
  reg  ex_ctrl_ren2;
  wire T396;
  wire req_ren1;
  reg  ex_ctrl_ren1;
  wire T397;
  wire req_wen;
  reg  ex_ctrl_wen;
  wire T398;
  wire fp_decoder_io_sigs_wen;
  wire req_ldst;
  reg  ex_ctrl_ldst;
  wire T399;
  wire[4:0] req_cmd;
  reg [4:0] ex_ctrl_cmd;
  wire[4:0] T400;
  wire[4:0] fp_decoder_io_sigs_cmd;
  wire T401;
  wire[64:0] T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire[4:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire[63:0] fpiu_io_out_bits_toint;
  wire[63:0] fpiu_io_out_bits_store;
  wire[4:0] T413;
  wire[4:0] T414;
  wire[4:0] T415;
  wire[4:0] T416;
  wire[4:0] fpmu_io_out_bits_exc;
  wire[4:0] ifpu_io_out_bits_exc;
  wire T417;
  wire[1:0] T418;
  wire[4:0] T419;
  wire[4:0] sfma_io_out_bits_exc;
  wire[4:0] dfma_io_out_bits_exc;
  wire T420;
  wire T421;
  wire T422;
  wire[4:0] T423;
  reg [4:0] wb_toint_exc;
  wire[4:0] T424;
  wire[4:0] fpiu_io_out_bits_exc;
  reg  mem_ctrl_toint;
  wire T425;
  wire wb_toint_valid;
  reg  wb_ctrl_toint;
  wire T426;
  reg  wb_reg_valid;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  reg  R433;
  wire T434;
  wire T435;
  wire T436;
  wire fp_inflight;
  wire T437;
  wire T438;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      regfile[initvar] = {3{$random}};
    winfo_0 = {1{$random}};
    winfo_1 = {1{$random}};
    mem_reg_inst = {1{$random}};
    ex_reg_inst = {1{$random}};
    ex_reg_valid = {1{$random}};
    mem_ctrl_single = {1{$random}};
    ex_ctrl_single = {1{$random}};
    mem_ctrl_fma = {1{$random}};
    ex_ctrl_fma = {1{$random}};
    mem_ctrl_fromint = {1{$random}};
    ex_ctrl_fromint = {1{$random}};
    mem_ctrl_fastpipe = {1{$random}};
    ex_ctrl_fastpipe = {1{$random}};
    write_port_busy = {1{$random}};
    wen = {1{$random}};
    mem_reg_valid = {1{$random}};
    load_wb_data = {2{$random}};
    load_wb_single = {1{$random}};
    load_wb = {1{$random}};
    load_wb_tag = {1{$random}};
    ex_ra3 = {1{$random}};
    ex_ra2 = {1{$random}};
    ex_ra1 = {1{$random}};
    ex_ctrl_round = {1{$random}};
    ex_ctrl_toint = {1{$random}};
    ex_ctrl_swap23 = {1{$random}};
    ex_ctrl_ren3 = {1{$random}};
    ex_ctrl_ren2 = {1{$random}};
    ex_ctrl_ren1 = {1{$random}};
    ex_ctrl_wen = {1{$random}};
    ex_ctrl_ldst = {1{$random}};
    ex_ctrl_cmd = {1{$random}};
    wb_toint_exc = {1{$random}};
    mem_ctrl_toint = {1{$random}};
    wb_ctrl_toint = {1{$random}};
    wb_reg_valid = {1{$random}};
    R433 = {1{$random}};
  end
`endif

  assign req_in3 = T0;
  assign T0 = regfile[ex_ra3];
  assign T2 = T3[7'h40:1'h0];
  assign T3 = T101 ? T97 : T4;
  assign T4 = {32'h0, T5};
  assign T5 = T6 ? ifpu_io_out_bits_data : fpmu_io_out_bits_data;
  assign T6 = T7[1'h0:1'h0];
  assign T7 = wsrc;
  assign wsrc = winfo_0 >> 3'h5;
  assign T8 = T93 ? mem_winfo : T9;
  assign T9 = T92 ? winfo_1 : winfo_0;
  assign T10 = T30 ? mem_winfo : winfo_1;
  assign mem_winfo = {T15, T11};
  assign T11 = mem_reg_inst[4'hb:3'h7];
  assign T12 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T13 = io_ctrl_valid ? io_dpath_inst : ex_reg_inst;
  assign T14 = reset ? 1'h0 : io_ctrl_valid;
  assign T15 = T23 | T16;
  assign T16 = T17 ? 2'h3 : 2'h0;
  assign T17 = mem_ctrl_fma & T18;
  assign T18 = mem_ctrl_single ^ 1'h1;
  assign T19 = ex_reg_valid ? ex_ctrl_single : mem_ctrl_single;
  assign T20 = io_ctrl_valid ? fp_decoder_io_sigs_single : ex_ctrl_single;
  assign T21 = ex_reg_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign T22 = io_ctrl_valid ? fp_decoder_io_sigs_fma : ex_ctrl_fma;
  assign T23 = T26 | T24;
  assign T24 = T25 ? 2'h2 : 2'h0;
  assign T25 = mem_ctrl_fma & mem_ctrl_single;
  assign T26 = {1'h0, T27};
  assign T27 = 1'h0 | mem_ctrl_fromint;
  assign T28 = ex_reg_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign T29 = io_ctrl_valid ? fp_decoder_io_sigs_fromint : ex_ctrl_fromint;
  assign T30 = mem_wen & T31;
  assign T31 = T44 & T32;
  assign T32 = memLatencyMask[1'h1:1'h1];
  assign memLatencyMask = T36 | T33;
  assign T33 = T34 ? 2'h2 : 2'h0;
  assign T34 = mem_ctrl_fma & T35;
  assign T35 = mem_ctrl_single ^ 1'h1;
  assign T36 = T39 | T37;
  assign T37 = {1'h0, T38};
  assign T38 = mem_ctrl_fma & mem_ctrl_single;
  assign T39 = T41 | T40;
  assign T40 = mem_ctrl_fromint ? 2'h2 : 2'h0;
  assign T41 = {1'h0, mem_ctrl_fastpipe};
  assign T42 = ex_reg_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign T43 = io_ctrl_valid ? fp_decoder_io_sigs_fastpipe : ex_ctrl_fastpipe;
  assign T44 = write_port_busy ^ 1'h1;
  assign T45 = ex_reg_valid ? T46 : write_port_busy;
  assign T46 = T76 | T47;
  assign T47 = T48 != 4'h0;
  assign T48 = T61 & T49;
  assign T49 = T53 | T50;
  assign T50 = T51 ? 4'h8 : 4'h0;
  assign T51 = ex_ctrl_fma & T52;
  assign T52 = ex_ctrl_single ^ 1'h1;
  assign T53 = T57 | T54;
  assign T54 = {1'h0, T55};
  assign T55 = T56 ? 3'h4 : 3'h0;
  assign T56 = ex_ctrl_fma & ex_ctrl_single;
  assign T57 = T59 | T58;
  assign T58 = ex_ctrl_fromint ? 4'h8 : 4'h0;
  assign T59 = {1'h0, T60};
  assign T60 = ex_ctrl_fastpipe ? 3'h4 : 3'h0;
  assign T61 = {2'h0, wen};
  assign T62 = reset ? 2'h0 : T63;
  assign T63 = T69 ? T66 : T64;
  assign T64 = {1'h0, T65};
  assign T65 = wen >> 1'h1;
  assign T66 = T67 | memLatencyMask;
  assign T67 = {1'h0, T68};
  assign T68 = wen >> 1'h1;
  assign T69 = mem_wen & T70;
  assign T70 = killm ^ 1'h1;
  assign killm = io_ctrl_killm | io_ctrl_nack_mem;
  assign mem_wen = mem_reg_valid & T71;
  assign T71 = T72 | mem_ctrl_fromint;
  assign T72 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T73 = reset ? 1'h0 : T74;
  assign T74 = ex_reg_valid & T75;
  assign T75 = io_ctrl_killx ^ 1'h1;
  assign T76 = mem_wen & T77;
  assign T77 = T78 != 3'h0;
  assign T78 = T91 & T79;
  assign T79 = T83 | T80;
  assign T80 = T81 ? 3'h4 : 3'h0;
  assign T81 = ex_ctrl_fma & T82;
  assign T82 = ex_ctrl_single ^ 1'h1;
  assign T83 = T87 | T84;
  assign T84 = {1'h0, T85};
  assign T85 = T86 ? 2'h2 : 2'h0;
  assign T86 = ex_ctrl_fma & ex_ctrl_single;
  assign T87 = T89 | T88;
  assign T88 = ex_ctrl_fromint ? 3'h4 : 3'h0;
  assign T89 = {1'h0, T90};
  assign T90 = ex_ctrl_fastpipe ? 2'h2 : 2'h0;
  assign T91 = {1'h0, memLatencyMask};
  assign T92 = wen[1'h1:1'h1];
  assign T93 = mem_wen & T94;
  assign T94 = T96 & T95;
  assign T95 = memLatencyMask[1'h0:1'h0];
  assign T96 = write_port_busy ^ 1'h1;
  assign T97 = T100 ? T99 : T98;
  assign T98 = {32'hffffffff, sfma_io_out_bits_data};
  assign T99 = {32'h0, dfma_io_out_bits_data};
  assign T100 = T7[1'h0:1'h0];
  assign T101 = T7[1'h1:1'h1];
  assign T102 = wen[1'h0:1'h0];
  assign T103 = waddr[3'h4:1'h0];
  assign waddr = T104;
  assign T104 = winfo_0[3'h4:1'h0];
  assign load_wb_data_recoded = load_wb_single ? T265 : rec_d;
  assign rec_d = {T264, T106};
  assign T106 = {T242, T107};
  assign T107 = T240 ? T110 : T108;
  assign T108 = load_wb_data[6'h33:1'h0];
  assign T109 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_data : load_wb_data;
  assign T110 = T111[6'h3e:4'hb];
  assign T111 = T177 << T112;
  assign T112 = ~ T113;
  assign T113 = T239 ? 6'h3f : T114;
  assign T114 = T238 ? 6'h3e : T115;
  assign T115 = T237 ? 6'h3d : T116;
  assign T116 = T236 ? 6'h3c : T117;
  assign T117 = T235 ? 6'h3b : T118;
  assign T118 = T234 ? 6'h3a : T119;
  assign T119 = T233 ? 6'h39 : T120;
  assign T120 = T232 ? 6'h38 : T121;
  assign T121 = T231 ? 6'h37 : T122;
  assign T122 = T230 ? 6'h36 : T123;
  assign T123 = T229 ? 6'h35 : T124;
  assign T124 = T228 ? 6'h34 : T125;
  assign T125 = T227 ? 6'h33 : T126;
  assign T126 = T226 ? 6'h32 : T127;
  assign T127 = T225 ? 6'h31 : T128;
  assign T128 = T224 ? 6'h30 : T129;
  assign T129 = T223 ? 6'h2f : T130;
  assign T130 = T222 ? 6'h2e : T131;
  assign T131 = T221 ? 6'h2d : T132;
  assign T132 = T220 ? 6'h2c : T133;
  assign T133 = T219 ? 6'h2b : T134;
  assign T134 = T218 ? 6'h2a : T135;
  assign T135 = T217 ? 6'h29 : T136;
  assign T136 = T216 ? 6'h28 : T137;
  assign T137 = T215 ? 6'h27 : T138;
  assign T138 = T214 ? 6'h26 : T139;
  assign T139 = T213 ? 6'h25 : T140;
  assign T140 = T212 ? 6'h24 : T141;
  assign T141 = T211 ? 6'h23 : T142;
  assign T142 = T210 ? 6'h22 : T143;
  assign T143 = T209 ? 6'h21 : T144;
  assign T144 = T208 ? 6'h20 : T145;
  assign T145 = T207 ? 5'h1f : T146;
  assign T146 = T206 ? 5'h1e : T147;
  assign T147 = T205 ? 5'h1d : T148;
  assign T148 = T204 ? 5'h1c : T149;
  assign T149 = T203 ? 5'h1b : T150;
  assign T150 = T202 ? 5'h1a : T151;
  assign T151 = T201 ? 5'h19 : T152;
  assign T152 = T200 ? 5'h18 : T153;
  assign T153 = T199 ? 5'h17 : T154;
  assign T154 = T198 ? 5'h16 : T155;
  assign T155 = T197 ? 5'h15 : T156;
  assign T156 = T196 ? 5'h14 : T157;
  assign T157 = T195 ? 5'h13 : T158;
  assign T158 = T194 ? 5'h12 : T159;
  assign T159 = T193 ? 5'h11 : T160;
  assign T160 = T192 ? 5'h10 : T161;
  assign T161 = T191 ? 4'hf : T162;
  assign T162 = T190 ? 4'he : T163;
  assign T163 = T189 ? 4'hd : T164;
  assign T164 = T188 ? 4'hc : T165;
  assign T165 = T187 ? 4'hb : T166;
  assign T166 = T186 ? 4'ha : T167;
  assign T167 = T185 ? 4'h9 : T168;
  assign T168 = T184 ? 4'h8 : T169;
  assign T169 = T183 ? 3'h7 : T170;
  assign T170 = T182 ? 3'h6 : T171;
  assign T171 = T181 ? 3'h5 : T172;
  assign T172 = T180 ? 3'h4 : T173;
  assign T173 = T179 ? 2'h3 : T174;
  assign T174 = T178 ? 2'h2 : T175;
  assign T175 = T176[1'h1:1'h1];
  assign T176 = T177[6'h3f:1'h0];
  assign T177 = T108 << 4'hc;
  assign T178 = T176[2'h2:2'h2];
  assign T179 = T176[2'h3:2'h3];
  assign T180 = T176[3'h4:3'h4];
  assign T181 = T176[3'h5:3'h5];
  assign T182 = T176[3'h6:3'h6];
  assign T183 = T176[3'h7:3'h7];
  assign T184 = T176[4'h8:4'h8];
  assign T185 = T176[4'h9:4'h9];
  assign T186 = T176[4'ha:4'ha];
  assign T187 = T176[4'hb:4'hb];
  assign T188 = T176[4'hc:4'hc];
  assign T189 = T176[4'hd:4'hd];
  assign T190 = T176[4'he:4'he];
  assign T191 = T176[4'hf:4'hf];
  assign T192 = T176[5'h10:5'h10];
  assign T193 = T176[5'h11:5'h11];
  assign T194 = T176[5'h12:5'h12];
  assign T195 = T176[5'h13:5'h13];
  assign T196 = T176[5'h14:5'h14];
  assign T197 = T176[5'h15:5'h15];
  assign T198 = T176[5'h16:5'h16];
  assign T199 = T176[5'h17:5'h17];
  assign T200 = T176[5'h18:5'h18];
  assign T201 = T176[5'h19:5'h19];
  assign T202 = T176[5'h1a:5'h1a];
  assign T203 = T176[5'h1b:5'h1b];
  assign T204 = T176[5'h1c:5'h1c];
  assign T205 = T176[5'h1d:5'h1d];
  assign T206 = T176[5'h1e:5'h1e];
  assign T207 = T176[5'h1f:5'h1f];
  assign T208 = T176[6'h20:6'h20];
  assign T209 = T176[6'h21:6'h21];
  assign T210 = T176[6'h22:6'h22];
  assign T211 = T176[6'h23:6'h23];
  assign T212 = T176[6'h24:6'h24];
  assign T213 = T176[6'h25:6'h25];
  assign T214 = T176[6'h26:6'h26];
  assign T215 = T176[6'h27:6'h27];
  assign T216 = T176[6'h28:6'h28];
  assign T217 = T176[6'h29:6'h29];
  assign T218 = T176[6'h2a:6'h2a];
  assign T219 = T176[6'h2b:6'h2b];
  assign T220 = T176[6'h2c:6'h2c];
  assign T221 = T176[6'h2d:6'h2d];
  assign T222 = T176[6'h2e:6'h2e];
  assign T223 = T176[6'h2f:6'h2f];
  assign T224 = T176[6'h30:6'h30];
  assign T225 = T176[6'h31:6'h31];
  assign T226 = T176[6'h32:6'h32];
  assign T227 = T176[6'h33:6'h33];
  assign T228 = T176[6'h34:6'h34];
  assign T229 = T176[6'h35:6'h35];
  assign T230 = T176[6'h36:6'h36];
  assign T231 = T176[6'h37:6'h37];
  assign T232 = T176[6'h38:6'h38];
  assign T233 = T176[6'h39:6'h39];
  assign T234 = T176[6'h3a:6'h3a];
  assign T235 = T176[6'h3b:6'h3b];
  assign T236 = T176[6'h3c:6'h3c];
  assign T237 = T176[6'h3d:6'h3d];
  assign T238 = T176[6'h3e:6'h3e];
  assign T239 = T176[6'h3f:6'h3f];
  assign T240 = T241 == 11'h0;
  assign T241 = load_wb_data[6'h3e:6'h34];
  assign T242 = T250 | T243;
  assign T243 = {2'h0, T244};
  assign T244 = T245 << 4'h9;
  assign T245 = T248 & T246;
  assign T246 = T247 ^ 1'h1;
  assign T247 = T108 == 52'h0;
  assign T248 = T249 == 2'h3;
  assign T249 = T250[4'hb:4'ha];
  assign T250 = T259 + T251;
  assign T251 = {1'h0, T252};
  assign T252 = T258 ? 11'h0 : T253;
  assign T253 = 11'h400 | T254;
  assign T254 = {9'h0, T255};
  assign T255 = T256 ? 2'h2 : 2'h1;
  assign T256 = T240 & T257;
  assign T257 = T247 ^ 1'h1;
  assign T258 = T240 & T247;
  assign T259 = T240 ? T261 : T260;
  assign T260 = {1'h0, T241};
  assign T261 = T247 ? 12'h0 : T262;
  assign T262 = {6'h3f, T263};
  assign T263 = ~ T112;
  assign T264 = load_wb_data[6'h3f:6'h3f];
  assign T265 = {32'hffffffff, rec_s};
  assign rec_s = {T359, T266};
  assign T266 = {T337, T267};
  assign T267 = T335 ? T269 : T268;
  assign T268 = load_wb_data[5'h16:1'h0];
  assign T269 = T270[5'h1e:4'h8];
  assign T270 = T304 << T271;
  assign T271 = ~ T272;
  assign T272 = T334 ? 5'h1f : T273;
  assign T273 = T333 ? 5'h1e : T274;
  assign T274 = T332 ? 5'h1d : T275;
  assign T275 = T331 ? 5'h1c : T276;
  assign T276 = T330 ? 5'h1b : T277;
  assign T277 = T329 ? 5'h1a : T278;
  assign T278 = T328 ? 5'h19 : T279;
  assign T279 = T327 ? 5'h18 : T280;
  assign T280 = T326 ? 5'h17 : T281;
  assign T281 = T325 ? 5'h16 : T282;
  assign T282 = T324 ? 5'h15 : T283;
  assign T283 = T323 ? 5'h14 : T284;
  assign T284 = T322 ? 5'h13 : T285;
  assign T285 = T321 ? 5'h12 : T286;
  assign T286 = T320 ? 5'h11 : T287;
  assign T287 = T319 ? 5'h10 : T288;
  assign T288 = T318 ? 4'hf : T289;
  assign T289 = T317 ? 4'he : T290;
  assign T290 = T316 ? 4'hd : T291;
  assign T291 = T315 ? 4'hc : T292;
  assign T292 = T314 ? 4'hb : T293;
  assign T293 = T313 ? 4'ha : T294;
  assign T294 = T312 ? 4'h9 : T295;
  assign T295 = T311 ? 4'h8 : T296;
  assign T296 = T310 ? 3'h7 : T297;
  assign T297 = T309 ? 3'h6 : T298;
  assign T298 = T308 ? 3'h5 : T299;
  assign T299 = T307 ? 3'h4 : T300;
  assign T300 = T306 ? 2'h3 : T301;
  assign T301 = T305 ? 2'h2 : T302;
  assign T302 = T303[1'h1:1'h1];
  assign T303 = T304[5'h1f:1'h0];
  assign T304 = T268 << 4'h9;
  assign T305 = T303[2'h2:2'h2];
  assign T306 = T303[2'h3:2'h3];
  assign T307 = T303[3'h4:3'h4];
  assign T308 = T303[3'h5:3'h5];
  assign T309 = T303[3'h6:3'h6];
  assign T310 = T303[3'h7:3'h7];
  assign T311 = T303[4'h8:4'h8];
  assign T312 = T303[4'h9:4'h9];
  assign T313 = T303[4'ha:4'ha];
  assign T314 = T303[4'hb:4'hb];
  assign T315 = T303[4'hc:4'hc];
  assign T316 = T303[4'hd:4'hd];
  assign T317 = T303[4'he:4'he];
  assign T318 = T303[4'hf:4'hf];
  assign T319 = T303[5'h10:5'h10];
  assign T320 = T303[5'h11:5'h11];
  assign T321 = T303[5'h12:5'h12];
  assign T322 = T303[5'h13:5'h13];
  assign T323 = T303[5'h14:5'h14];
  assign T324 = T303[5'h15:5'h15];
  assign T325 = T303[5'h16:5'h16];
  assign T326 = T303[5'h17:5'h17];
  assign T327 = T303[5'h18:5'h18];
  assign T328 = T303[5'h19:5'h19];
  assign T329 = T303[5'h1a:5'h1a];
  assign T330 = T303[5'h1b:5'h1b];
  assign T331 = T303[5'h1c:5'h1c];
  assign T332 = T303[5'h1d:5'h1d];
  assign T333 = T303[5'h1e:5'h1e];
  assign T334 = T303[5'h1f:5'h1f];
  assign T335 = T336 == 8'h0;
  assign T336 = load_wb_data[5'h1e:5'h17];
  assign T337 = T345 | T338;
  assign T338 = {2'h0, T339};
  assign T339 = T340 << 3'h6;
  assign T340 = T343 & T341;
  assign T341 = T342 ^ 1'h1;
  assign T342 = T268 == 23'h0;
  assign T343 = T344 == 2'h3;
  assign T344 = T345[4'h8:3'h7];
  assign T345 = T354 + T346;
  assign T346 = {1'h0, T347};
  assign T347 = T353 ? 8'h0 : T348;
  assign T348 = 8'h80 | T349;
  assign T349 = {6'h0, T350};
  assign T350 = T351 ? 2'h2 : 2'h1;
  assign T351 = T335 & T352;
  assign T352 = T342 ^ 1'h1;
  assign T353 = T335 & T342;
  assign T354 = T335 ? T356 : T355;
  assign T355 = {1'h0, T336};
  assign T356 = T342 ? 9'h0 : T357;
  assign T357 = {4'hf, T358};
  assign T358 = ~ T271;
  assign T359 = load_wb_data[5'h1f:5'h1f];
  assign T360 = io_dpath_dmem_resp_val ? T361 : load_wb_single;
  assign T361 = T363 | T362;
  assign T362 = io_dpath_dmem_resp_type == 3'h6;
  assign T363 = io_dpath_dmem_resp_type == 3'h2;
  assign T364 = io_dpath_dmem_resp_val ? io_dpath_dmem_resp_tag : load_wb_tag;
  assign T365 = T370 ? T369 : T366;
  assign T366 = T368 ? T367 : ex_ra3;
  assign T367 = io_dpath_inst[5'h1f:5'h1b];
  assign T368 = io_ctrl_valid & fp_decoder_io_sigs_ren3;
  assign T369 = io_dpath_inst[5'h18:5'h14];
  assign T370 = T373 & T371;
  assign T371 = T372 & fp_decoder_io_sigs_swap23;
  assign T372 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign T373 = io_ctrl_valid & fp_decoder_io_sigs_ren2;
  assign req_in2 = T374;
  assign T374 = regfile[ex_ra2];
  assign T375 = T377 ? T376 : ex_ra2;
  assign T376 = io_dpath_inst[5'h18:5'h14];
  assign T377 = T373 & T378;
  assign T378 = T380 & T379;
  assign T379 = fp_decoder_io_sigs_swap23 ^ 1'h1;
  assign T380 = fp_decoder_io_sigs_ldst ^ 1'h1;
  assign req_in1 = T381;
  assign T381 = regfile[ex_ra1];
  assign T382 = T387 ? T386 : T383;
  assign T383 = T385 ? T384 : ex_ra1;
  assign T384 = io_dpath_inst[5'h13:4'hf];
  assign T385 = io_ctrl_valid & fp_decoder_io_sigs_ren1;
  assign T386 = io_dpath_inst[5'h18:5'h14];
  assign T387 = T373 & fp_decoder_io_sigs_ldst;
  assign req_typ = T388;
  assign T388 = ex_reg_inst[5'h15:5'h14];
  assign req_rm = ex_rm;
  assign ex_rm = T390 ? io_dpath_fcsr_rm : T389;
  assign T389 = ex_reg_inst[4'he:4'hc];
  assign T390 = T391 == 3'h7;
  assign T391 = ex_reg_inst[4'he:4'hc];
  assign req_round = ex_ctrl_round;
  assign T392 = io_ctrl_valid ? fp_decoder_io_sigs_round : ex_ctrl_round;
  assign req_fma = ex_ctrl_fma;
  assign req_fastpipe = ex_ctrl_fastpipe;
  assign req_toint = ex_ctrl_toint;
  assign T393 = io_ctrl_valid ? fp_decoder_io_sigs_toint : ex_ctrl_toint;
  assign req_fromint = ex_ctrl_fromint;
  assign req_single = ex_ctrl_single;
  assign req_swap23 = ex_ctrl_swap23;
  assign T394 = io_ctrl_valid ? fp_decoder_io_sigs_swap23 : ex_ctrl_swap23;
  assign req_ren3 = ex_ctrl_ren3;
  assign T395 = io_ctrl_valid ? fp_decoder_io_sigs_ren3 : ex_ctrl_ren3;
  assign req_ren2 = ex_ctrl_ren2;
  assign T396 = io_ctrl_valid ? fp_decoder_io_sigs_ren2 : ex_ctrl_ren2;
  assign req_ren1 = ex_ctrl_ren1;
  assign T397 = io_ctrl_valid ? fp_decoder_io_sigs_ren1 : ex_ctrl_ren1;
  assign req_wen = ex_ctrl_wen;
  assign T398 = io_ctrl_valid ? fp_decoder_io_sigs_wen : ex_ctrl_wen;
  assign req_ldst = ex_ctrl_ldst;
  assign T399 = io_ctrl_valid ? fp_decoder_io_sigs_ldst : ex_ctrl_ldst;
  assign req_cmd = ex_ctrl_cmd;
  assign T400 = io_ctrl_valid ? fp_decoder_io_sigs_cmd : ex_ctrl_cmd;
  assign T401 = ex_reg_valid & ex_ctrl_fastpipe;
  assign T402 = {1'h0, io_dpath_fromint_data};
  assign T403 = ex_reg_valid & ex_ctrl_fromint;
  assign T404 = ex_reg_valid & T405;
  assign T405 = ex_ctrl_toint | T406;
  assign T406 = T407 == 5'h5;
  assign T407 = ex_ctrl_cmd & 5'hd;
  assign T408 = T410 & T409;
  assign T409 = ex_ctrl_single ^ 1'h1;
  assign T410 = ex_reg_valid & ex_ctrl_fma;
  assign T411 = T412 & ex_ctrl_single;
  assign T412 = ex_reg_valid & ex_ctrl_fma;
  assign io_dpath_toint_data = fpiu_io_out_bits_toint;
  assign io_dpath_store_data = fpiu_io_out_bits_store;
  assign io_dpath_fcsr_flags_bits = T413;
  assign T413 = T423 | T414;
  assign T414 = T422 ? T415 : 5'h0;
  assign T415 = T421 ? T419 : T416;
  assign T416 = T417 ? ifpu_io_out_bits_exc : fpmu_io_out_bits_exc;
  assign T417 = T418[1'h0:1'h0];
  assign T418 = wsrc;
  assign T419 = T420 ? dfma_io_out_bits_exc : sfma_io_out_bits_exc;
  assign T420 = T418[1'h0:1'h0];
  assign T421 = T418[1'h1:1'h1];
  assign T422 = wen[1'h0:1'h0];
  assign T423 = wb_toint_valid ? wb_toint_exc : 5'h0;
  assign T424 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T425 = ex_reg_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign T426 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign T427 = reset ? 1'h0 : T428;
  assign T428 = mem_reg_valid & T429;
  assign T429 = killm ^ 1'h1;
  assign io_dpath_fcsr_flags_valid = T430;
  assign T430 = wb_toint_valid | T431;
  assign T431 = wen[1'h0:1'h0];
  assign io_ctrl_sboard_clra = waddr;
  assign io_ctrl_sboard_clr = 1'h0;
  assign io_ctrl_sboard_set = T432;
  assign T432 = wb_reg_valid & R433;
  assign io_ctrl_dec_round = fp_decoder_io_sigs_round;
  assign io_ctrl_dec_fma = fp_decoder_io_sigs_fma;
  assign io_ctrl_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_ctrl_dec_toint = fp_decoder_io_sigs_toint;
  assign io_ctrl_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_ctrl_dec_single = fp_decoder_io_sigs_single;
  assign io_ctrl_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_ctrl_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_ctrl_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_ctrl_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_ctrl_dec_wen = fp_decoder_io_sigs_wen;
  assign io_ctrl_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_ctrl_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_ctrl_illegal_rm = T434;
  assign T434 = T435 & ex_ctrl_round;
  assign T435 = ex_rm[2'h2:2'h2];
  assign io_ctrl_nack_mem = write_port_busy;
  assign io_ctrl_fcsr_rdy = T436;
  assign T436 = fp_inflight ^ 1'h1;
  assign fp_inflight = T438 | T437;
  assign T437 = wen != 2'h0;
  assign T438 = wb_reg_valid & wb_ctrl_toint;
  FPUDecoder fp_decoder(
       .io_inst( io_dpath_inst ),
       .io_sigs_cmd( fp_decoder_io_sigs_cmd ),
       .io_sigs_ldst( fp_decoder_io_sigs_ldst ),
       .io_sigs_wen( fp_decoder_io_sigs_wen ),
       .io_sigs_ren1( fp_decoder_io_sigs_ren1 ),
       .io_sigs_ren2( fp_decoder_io_sigs_ren2 ),
       .io_sigs_ren3( fp_decoder_io_sigs_ren3 ),
       .io_sigs_swap23( fp_decoder_io_sigs_swap23 ),
       .io_sigs_single( fp_decoder_io_sigs_single ),
       .io_sigs_fromint( fp_decoder_io_sigs_fromint ),
       .io_sigs_toint( fp_decoder_io_sigs_toint ),
       .io_sigs_fastpipe( fp_decoder_io_sigs_fastpipe ),
       .io_sigs_fma( fp_decoder_io_sigs_fma ),
       .io_sigs_round( fp_decoder_io_sigs_round )
  );
  FPUFMAPipe_0 sfma(.clk(clk), .reset(reset),
       .io_in_valid( T411 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( sfma_io_out_bits_data ),
       .io_out_bits_exc( sfma_io_out_bits_exc )
  );
  FPUFMAPipe_1 dfma(.clk(clk), .reset(reset),
       .io_in_valid( T408 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( dfma_io_out_bits_data ),
       .io_out_bits_exc( dfma_io_out_bits_exc )
  );
  FPToInt fpiu(.clk(clk),
       .io_in_valid( T404 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_lt( fpiu_io_out_bits_lt ),
       .io_out_bits_store( fpiu_io_out_bits_store ),
       .io_out_bits_toint( fpiu_io_out_bits_toint ),
       .io_out_bits_exc( fpiu_io_out_bits_exc )
  );
  IntToFP ifpu(.clk(clk), .reset(reset),
       .io_in_valid( T403 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( T402 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( ifpu_io_out_bits_data ),
       .io_out_bits_exc( ifpu_io_out_bits_exc )
  );
  FPToFP fpmu(.clk(clk), .reset(reset),
       .io_in_valid( T401 ),
       .io_in_bits_cmd( req_cmd ),
       .io_in_bits_ldst( req_ldst ),
       .io_in_bits_wen( req_wen ),
       .io_in_bits_ren1( req_ren1 ),
       .io_in_bits_ren2( req_ren2 ),
       .io_in_bits_ren3( req_ren3 ),
       .io_in_bits_swap23( req_swap23 ),
       .io_in_bits_single( req_single ),
       .io_in_bits_fromint( req_fromint ),
       .io_in_bits_toint( req_toint ),
       .io_in_bits_fastpipe( req_fastpipe ),
       .io_in_bits_fma( req_fma ),
       .io_in_bits_round( req_round ),
       .io_in_bits_rm( req_rm ),
       .io_in_bits_typ( req_typ ),
       .io_in_bits_in1( req_in1 ),
       .io_in_bits_in2( req_in2 ),
       .io_in_bits_in3( req_in3 ),
       //.io_out_valid(  )
       .io_out_bits_data( fpmu_io_out_bits_data ),
       .io_out_bits_exc( fpmu_io_out_bits_exc ),
       .io_lt( fpiu_io_out_bits_lt )
  );

  always @(posedge clk) begin
    if (T102)
      regfile[T103] <= T2;
    if(T93) begin
      winfo_0 <= mem_winfo;
    end else if(T92) begin
      winfo_0 <= winfo_1;
    end
    if(T30) begin
      winfo_1 <= mem_winfo;
    end
    if(ex_reg_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if(io_ctrl_valid) begin
      ex_reg_inst <= io_dpath_inst;
    end
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_ctrl_valid;
    end
    if(ex_reg_valid) begin
      mem_ctrl_single <= ex_ctrl_single;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_single <= fp_decoder_io_sigs_single;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fma <= ex_ctrl_fma;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fma <= fp_decoder_io_sigs_fma;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fromint <= ex_ctrl_fromint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fromint <= fp_decoder_io_sigs_fromint;
    end
    if(ex_reg_valid) begin
      mem_ctrl_fastpipe <= ex_ctrl_fastpipe;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_fastpipe <= fp_decoder_io_sigs_fastpipe;
    end
    if(ex_reg_valid) begin
      write_port_busy <= T46;
    end
    if(reset) begin
      wen <= 2'h0;
    end else if(T69) begin
      wen <= T66;
    end else begin
      wen <= T64;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T74;
    end
    if (load_wb)
      regfile[load_wb_tag] <= load_wb_data_recoded;
    if(io_dpath_dmem_resp_val) begin
      load_wb_data <= io_dpath_dmem_resp_data;
    end
    if(io_dpath_dmem_resp_val) begin
      load_wb_single <= T361;
    end
    load_wb <= io_dpath_dmem_resp_val;
    if(io_dpath_dmem_resp_val) begin
      load_wb_tag <= io_dpath_dmem_resp_tag;
    end
    if(T370) begin
      ex_ra3 <= T369;
    end else if(T368) begin
      ex_ra3 <= T367;
    end
    if(T377) begin
      ex_ra2 <= T376;
    end
    if(T387) begin
      ex_ra1 <= T386;
    end else if(T385) begin
      ex_ra1 <= T384;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_round <= fp_decoder_io_sigs_round;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_toint <= fp_decoder_io_sigs_toint;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_swap23 <= fp_decoder_io_sigs_swap23;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren3 <= fp_decoder_io_sigs_ren3;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren2 <= fp_decoder_io_sigs_ren2;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ren1 <= fp_decoder_io_sigs_ren1;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_wen <= fp_decoder_io_sigs_wen;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_ldst <= fp_decoder_io_sigs_ldst;
    end
    if(io_ctrl_valid) begin
      ex_ctrl_cmd <= fp_decoder_io_sigs_cmd;
    end
    if(mem_ctrl_toint) begin
      wb_toint_exc <= fpiu_io_out_bits_exc;
    end
    if(ex_reg_valid) begin
      mem_ctrl_toint <= ex_ctrl_toint;
    end
    if(mem_reg_valid) begin
      wb_ctrl_toint <= mem_ctrl_toint;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T428;
    end
    R433 <= 1'h0;
  end
endmodule

module Core(input clk, input reset,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr,
    output io_imem_req_valid,
    output[43:0] io_imem_req_bits_pc,
    output io_imem_resp_ready,
    input  io_imem_resp_valid,
    input [43:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input  io_imem_resp_bits_xcpt_ma,
    input  io_imem_resp_bits_xcpt_if,
    input  io_imem_btb_resp_valid,
    input  io_imem_btb_resp_bits_taken,
    input [42:0] io_imem_btb_resp_bits_target,
    input [2:0] io_imem_btb_resp_bits_entry,
    input [3:0] io_imem_btb_resp_bits_bht_index,
    input [1:0] io_imem_btb_resp_bits_bht_value,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output[42:0] io_imem_btb_update_bits_prediction_bits_target,
    output[2:0] io_imem_btb_update_bits_prediction_bits_entry,
    output[3:0] io_imem_btb_update_bits_prediction_bits_bht_index,
    output[1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output[42:0] io_imem_btb_update_bits_pc,
    output[42:0] io_imem_btb_update_bits_target,
    output[42:0] io_imem_btb_update_bits_returnAddr,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isCall,
    output io_imem_btb_update_bits_isReturn,
    output io_imem_btb_update_bits_incorrectTarget,
    //output io_imem_ptw_req_ready
    input  io_imem_ptw_req_valid,
    input [29:0] io_imem_ptw_req_bits,
    //output io_imem_ptw_resp_valid
    //output io_imem_ptw_resp_bits_error
    //output[18:0] io_imem_ptw_resp_bits_ppn
    //output[5:0] io_imem_ptw_resp_bits_perm
    //output[7:0] io_imem_ptw_status_ip
    //output[7:0] io_imem_ptw_status_im
    //output[6:0] io_imem_ptw_status_zero
    //output io_imem_ptw_status_er
    //output io_imem_ptw_status_vm
    //output io_imem_ptw_status_s64
    //output io_imem_ptw_status_u64
    //output io_imem_ptw_status_ef
    //output io_imem_ptw_status_pei
    //output io_imem_ptw_status_ei
    //output io_imem_ptw_status_ps
    //output io_imem_ptw_status_s
    //output io_imem_ptw_invalidate
    //output io_imem_ptw_sret
    output io_imem_invalidate,
    input  io_dmem_req_ready,
    output io_dmem_req_valid,
    output io_dmem_req_bits_kill,
    output[2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output[43:0] io_dmem_req_bits_addr,
    output[63:0] io_dmem_req_bits_data,
    output[7:0] io_dmem_req_bits_tag,
    output[4:0] io_dmem_req_bits_cmd,
    input  io_dmem_resp_valid,
    input  io_dmem_resp_bits_nack,
    input  io_dmem_resp_bits_replay,
    input [2:0] io_dmem_resp_bits_typ,
    input  io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data,
    input [63:0] io_dmem_resp_bits_data_subword,
    input [7:0] io_dmem_resp_bits_tag,
    input [3:0] io_dmem_resp_bits_cmd,
    input [43:0] io_dmem_resp_bits_addr,
    input [63:0] io_dmem_resp_bits_store_data,
    input  io_dmem_replay_next_valid,
    input [7:0] io_dmem_replay_next_bits,
    input  io_dmem_xcpt_ma_ld,
    input  io_dmem_xcpt_ma_st,
    input  io_dmem_xcpt_pf_ld,
    input  io_dmem_xcpt_pf_st,
    //output io_dmem_ptw_req_ready
    input  io_dmem_ptw_req_valid,
    input [29:0] io_dmem_ptw_req_bits,
    //output io_dmem_ptw_resp_valid
    //output io_dmem_ptw_resp_bits_error
    //output[18:0] io_dmem_ptw_resp_bits_ppn
    //output[5:0] io_dmem_ptw_resp_bits_perm
    //output[7:0] io_dmem_ptw_status_ip
    //output[7:0] io_dmem_ptw_status_im
    //output[6:0] io_dmem_ptw_status_zero
    //output io_dmem_ptw_status_er
    //output io_dmem_ptw_status_vm
    //output io_dmem_ptw_status_s64
    //output io_dmem_ptw_status_u64
    //output io_dmem_ptw_status_ef
    //output io_dmem_ptw_status_pei
    //output io_dmem_ptw_status_ei
    //output io_dmem_ptw_status_ps
    //output io_dmem_ptw_status_s
    //output io_dmem_ptw_invalidate
    //output io_dmem_ptw_sret
    input  io_dmem_ordered,
    output[31:0] io_ptw_ptbr,
    output io_ptw_invalidate,
    output io_ptw_sret,
    output[7:0] io_ptw_status_ip,
    output[7:0] io_ptw_status_im,
    output[6:0] io_ptw_status_zero,
    output io_ptw_status_er,
    output io_ptw_status_vm,
    output io_ptw_status_s64,
    output io_ptw_status_u64,
    output io_ptw_status_ef,
    output io_ptw_status_pei,
    output io_ptw_status_ei,
    output io_ptw_status_ps,
    output io_ptw_status_s,
    input  io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output[6:0] io_rocc_cmd_bits_inst_funct,
    output[4:0] io_rocc_cmd_bits_inst_rs2,
    output[4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output[4:0] io_rocc_cmd_bits_inst_rd,
    output[6:0] io_rocc_cmd_bits_inst_opcode,
    output[63:0] io_rocc_cmd_bits_rs1,
    output[63:0] io_rocc_cmd_bits_rs2,
    //output io_rocc_resp_ready
    input  io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    //output io_rocc_mem_req_ready
    input  io_rocc_mem_req_valid,
    input  io_rocc_mem_req_bits_kill,
    input [2:0] io_rocc_mem_req_bits_typ,
    input  io_rocc_mem_req_bits_phys,
    input [43:0] io_rocc_mem_req_bits_addr,
    input [63:0] io_rocc_mem_req_bits_data,
    input [7:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    //output io_rocc_mem_resp_valid
    //output io_rocc_mem_resp_bits_nack
    //output io_rocc_mem_resp_bits_replay
    //output[2:0] io_rocc_mem_resp_bits_typ
    //output io_rocc_mem_resp_bits_has_data
    //output[63:0] io_rocc_mem_resp_bits_data
    //output[63:0] io_rocc_mem_resp_bits_data_subword
    //output[7:0] io_rocc_mem_resp_bits_tag
    //output[3:0] io_rocc_mem_resp_bits_cmd
    //output[43:0] io_rocc_mem_resp_bits_addr
    //output[63:0] io_rocc_mem_resp_bits_store_data
    //output io_rocc_mem_replay_next_valid
    //output[7:0] io_rocc_mem_replay_next_bits
    //output io_rocc_mem_xcpt_ma_ld
    //output io_rocc_mem_xcpt_ma_st
    //output io_rocc_mem_xcpt_pf_ld
    //output io_rocc_mem_xcpt_pf_st
    input  io_rocc_mem_ptw_req_ready,
    //output io_rocc_mem_ptw_req_valid
    //output[29:0] io_rocc_mem_ptw_req_bits
    input  io_rocc_mem_ptw_resp_valid,
    input  io_rocc_mem_ptw_resp_bits_error,
    input [18:0] io_rocc_mem_ptw_resp_bits_ppn,
    input [5:0] io_rocc_mem_ptw_resp_bits_perm,
    input [7:0] io_rocc_mem_ptw_status_ip,
    input [7:0] io_rocc_mem_ptw_status_im,
    input [6:0] io_rocc_mem_ptw_status_zero,
    input  io_rocc_mem_ptw_status_er,
    input  io_rocc_mem_ptw_status_vm,
    input  io_rocc_mem_ptw_status_s64,
    input  io_rocc_mem_ptw_status_u64,
    input  io_rocc_mem_ptw_status_ef,
    input  io_rocc_mem_ptw_status_pei,
    input  io_rocc_mem_ptw_status_ei,
    input  io_rocc_mem_ptw_status_ps,
    input  io_rocc_mem_ptw_status_s,
    input  io_rocc_mem_ptw_invalidate,
    input  io_rocc_mem_ptw_sret,
    //output io_rocc_mem_ordered
    input  io_rocc_busy,
    output io_rocc_s,
    input  io_rocc_interrupt,
    //output io_rocc_imem_acquire_ready
    input  io_rocc_imem_acquire_valid,
    input [1:0] io_rocc_imem_acquire_bits_header_src,
    input [1:0] io_rocc_imem_acquire_bits_header_dst,
    input [25:0] io_rocc_imem_acquire_bits_payload_addr,
    input [1:0] io_rocc_imem_acquire_bits_payload_client_xact_id,
    input [511:0] io_rocc_imem_acquire_bits_payload_data,
    input [2:0] io_rocc_imem_acquire_bits_payload_a_type,
    input [5:0] io_rocc_imem_acquire_bits_payload_write_mask,
    input [2:0] io_rocc_imem_acquire_bits_payload_subword_addr,
    input [3:0] io_rocc_imem_acquire_bits_payload_atomic_opcode,
    input  io_rocc_imem_grant_ready,
    //output io_rocc_imem_grant_valid
    //output[1:0] io_rocc_imem_grant_bits_header_src
    //output[1:0] io_rocc_imem_grant_bits_header_dst
    //output[511:0] io_rocc_imem_grant_bits_payload_data
    //output[1:0] io_rocc_imem_grant_bits_payload_client_xact_id
    //output[2:0] io_rocc_imem_grant_bits_payload_master_xact_id
    //output[3:0] io_rocc_imem_grant_bits_payload_g_type
    //output io_rocc_imem_finish_ready
    input  io_rocc_imem_finish_valid,
    input [1:0] io_rocc_imem_finish_bits_header_src,
    input [1:0] io_rocc_imem_finish_bits_header_dst,
    input [2:0] io_rocc_imem_finish_bits_payload_master_xact_id,
    //output io_rocc_iptw_req_ready
    input  io_rocc_iptw_req_valid,
    input [29:0] io_rocc_iptw_req_bits,
    //output io_rocc_iptw_resp_valid
    //output io_rocc_iptw_resp_bits_error
    //output[18:0] io_rocc_iptw_resp_bits_ppn
    //output[5:0] io_rocc_iptw_resp_bits_perm
    //output[7:0] io_rocc_iptw_status_ip
    //output[7:0] io_rocc_iptw_status_im
    //output[6:0] io_rocc_iptw_status_zero
    //output io_rocc_iptw_status_er
    //output io_rocc_iptw_status_vm
    //output io_rocc_iptw_status_s64
    //output io_rocc_iptw_status_u64
    //output io_rocc_iptw_status_ef
    //output io_rocc_iptw_status_pei
    //output io_rocc_iptw_status_ei
    //output io_rocc_iptw_status_ps
    //output io_rocc_iptw_status_s
    //output io_rocc_iptw_invalidate
    //output io_rocc_iptw_sret
    //output io_rocc_dptw_req_ready
    input  io_rocc_dptw_req_valid,
    input [29:0] io_rocc_dptw_req_bits,
    //output io_rocc_dptw_resp_valid
    //output io_rocc_dptw_resp_bits_error
    //output[18:0] io_rocc_dptw_resp_bits_ppn
    //output[5:0] io_rocc_dptw_resp_bits_perm
    //output[7:0] io_rocc_dptw_status_ip
    //output[7:0] io_rocc_dptw_status_im
    //output[6:0] io_rocc_dptw_status_zero
    //output io_rocc_dptw_status_er
    //output io_rocc_dptw_status_vm
    //output io_rocc_dptw_status_s64
    //output io_rocc_dptw_status_u64
    //output io_rocc_dptw_status_ef
    //output io_rocc_dptw_status_pei
    //output io_rocc_dptw_status_ei
    //output io_rocc_dptw_status_ps
    //output io_rocc_dptw_status_s
    //output io_rocc_dptw_invalidate
    //output io_rocc_dptw_sret
    //output io_rocc_pptw_req_ready
    input  io_rocc_pptw_req_valid,
    input [29:0] io_rocc_pptw_req_bits,
    //output io_rocc_pptw_resp_valid
    //output io_rocc_pptw_resp_bits_error
    //output[18:0] io_rocc_pptw_resp_bits_ppn
    //output[5:0] io_rocc_pptw_resp_bits_perm
    //output[7:0] io_rocc_pptw_status_ip
    //output[7:0] io_rocc_pptw_status_im
    //output[6:0] io_rocc_pptw_status_zero
    //output io_rocc_pptw_status_er
    //output io_rocc_pptw_status_vm
    //output io_rocc_pptw_status_s64
    //output io_rocc_pptw_status_u64
    //output io_rocc_pptw_status_ef
    //output io_rocc_pptw_status_pei
    //output io_rocc_pptw_status_ei
    //output io_rocc_pptw_status_ps
    //output io_rocc_pptw_status_s
    //output io_rocc_pptw_invalidate
    //output io_rocc_pptw_sret
    output io_rocc_exception
);

  wire[63:0] dpath_io_fpu_dmem_resp_data;
  wire[4:0] dpath_io_fpu_dmem_resp_tag;
  wire[2:0] dpath_io_fpu_dmem_resp_type;
  wire dpath_io_fpu_dmem_resp_val;
  wire[2:0] dpath_io_fpu_fcsr_rm;
  wire[63:0] dpath_io_fpu_fromint_data;
  wire[31:0] dpath_io_fpu_inst;
  wire ctrl_io_fpu_killm;
  wire ctrl_io_fpu_killx;
  wire ctrl_io_fpu_valid;
  wire[63:0] FPU_io_dpath_toint_data;
  wire[63:0] FPU_io_dpath_store_data;
  wire[4:0] FPU_io_dpath_fcsr_flags_bits;
  wire FPU_io_dpath_fcsr_flags_valid;
  wire ctrl_io_dpath_badvaddr_wen;
  wire[63:0] ctrl_io_dpath_cause;
  wire ctrl_io_dpath_exception;
  wire ctrl_io_dpath_retire;
  wire ctrl_io_dpath_ll_ready;
  wire[1:0] ctrl_io_dpath_bypass_src_0;
  wire[1:0] ctrl_io_dpath_bypass_src_1;
  wire ctrl_io_dpath_bypass_0;
  wire ctrl_io_dpath_bypass_1;
  wire ctrl_io_dpath_mem_rocc_val;
  wire ctrl_io_dpath_ex_rocc_val;
  wire ctrl_io_dpath_ex_rs2_val;
  wire[2:0] ctrl_io_dpath_ex_mem_type;
  wire ctrl_io_dpath_wb_wen;
  wire ctrl_io_dpath_mem_wen;
  wire ctrl_io_dpath_mem_branch;
  wire ctrl_io_dpath_mem_jalr;
  wire ctrl_io_dpath_ex_valid;
  wire ctrl_io_dpath_ex_wen;
  wire ctrl_io_dpath_mem_fp_val;
  wire ctrl_io_dpath_ex_fp_val;
  wire ctrl_io_dpath_wb_load;
  wire ctrl_io_dpath_mem_load;
  wire ctrl_io_dpath_sret;
  wire[2:0] ctrl_io_dpath_csr;
  wire ctrl_io_dpath_div_mul_kill;
  wire ctrl_io_dpath_div_mul_val;
  wire[3:0] ctrl_io_dpath_fn_alu;
  wire ctrl_io_dpath_fn_dw;
  wire[2:0] ctrl_io_dpath_sel_imm;
  wire[1:0] ctrl_io_dpath_sel_alu1;
  wire[2:0] ctrl_io_dpath_sel_alu2;
  wire ctrl_io_dpath_ren_0;
  wire ctrl_io_dpath_ren_1;
  wire ctrl_io_dpath_killd;
  wire[2:0] ctrl_io_dpath_sel_pc;
  wire[4:0] FPU_io_ctrl_sboard_clra;
  wire FPU_io_ctrl_sboard_clr;
  wire FPU_io_ctrl_sboard_set;
  wire FPU_io_ctrl_dec_round;
  wire FPU_io_ctrl_dec_fma;
  wire FPU_io_ctrl_dec_fastpipe;
  wire FPU_io_ctrl_dec_toint;
  wire FPU_io_ctrl_dec_fromint;
  wire FPU_io_ctrl_dec_single;
  wire FPU_io_ctrl_dec_swap23;
  wire FPU_io_ctrl_dec_ren3;
  wire FPU_io_ctrl_dec_ren2;
  wire FPU_io_ctrl_dec_ren1;
  wire FPU_io_ctrl_dec_wen;
  wire FPU_io_ctrl_dec_ldst;
  wire[4:0] FPU_io_ctrl_dec_cmd;
  wire FPU_io_ctrl_illegal_rm;
  wire FPU_io_ctrl_nack_mem;
  wire FPU_io_ctrl_fcsr_rdy;
  wire dpath_io_ctrl_csr_replay;
  wire[4:0] dpath_io_ctrl_fp_sboard_clra;
  wire dpath_io_ctrl_fp_sboard_clr;
  wire dpath_io_ctrl_status_s;
  wire dpath_io_ctrl_status_ps;
  wire dpath_io_ctrl_status_ei;
  wire dpath_io_ctrl_status_pei;
  wire dpath_io_ctrl_status_ef;
  wire dpath_io_ctrl_status_u64;
  wire dpath_io_ctrl_status_s64;
  wire dpath_io_ctrl_status_vm;
  wire dpath_io_ctrl_status_er;
  wire[6:0] dpath_io_ctrl_status_zero;
  wire[7:0] dpath_io_ctrl_status_im;
  wire[7:0] dpath_io_ctrl_status_ip;
  wire[4:0] dpath_io_ctrl_wb_waddr;
  wire[4:0] dpath_io_ctrl_mem_waddr;
  wire dpath_io_ctrl_mem_rs1_ra;
  wire[4:0] dpath_io_ctrl_ex_waddr;
  wire[4:0] dpath_io_ctrl_ll_waddr;
  wire dpath_io_ctrl_ll_wen;
  wire dpath_io_ctrl_div_mul_rdy;
  wire dpath_io_ctrl_mem_misprediction;
  wire dpath_io_ctrl_mem_br_taken;
  wire[31:0] dpath_io_ctrl_inst;
  wire ctrl_io_rocc_exception;
  wire ctrl_io_rocc_s;
  wire[63:0] dpath_io_rocc_cmd_bits_rs2;
  wire[63:0] dpath_io_rocc_cmd_bits_rs1;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_opcode;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rd;
  wire dpath_io_rocc_cmd_bits_inst_xs2;
  wire dpath_io_rocc_cmd_bits_inst_xs1;
  wire dpath_io_rocc_cmd_bits_inst_xd;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs1;
  wire[4:0] dpath_io_rocc_cmd_bits_inst_rs2;
  wire[6:0] dpath_io_rocc_cmd_bits_inst_funct;
  wire ctrl_io_rocc_cmd_valid;
  wire dpath_io_ptw_status_s;
  wire dpath_io_ptw_status_ps;
  wire dpath_io_ptw_status_ei;
  wire dpath_io_ptw_status_pei;
  wire dpath_io_ptw_status_ef;
  wire dpath_io_ptw_status_u64;
  wire dpath_io_ptw_status_s64;
  wire dpath_io_ptw_status_vm;
  wire dpath_io_ptw_status_er;
  wire[6:0] dpath_io_ptw_status_zero;
  wire[7:0] dpath_io_ptw_status_im;
  wire[7:0] dpath_io_ptw_status_ip;
  wire dpath_io_ptw_sret;
  wire dpath_io_ptw_invalidate;
  wire[31:0] dpath_io_ptw_ptbr;
  wire[4:0] ctrl_io_dmem_req_bits_cmd;
  wire[7:0] dpath_io_dmem_req_bits_tag;
  wire[63:0] dpath_io_dmem_req_bits_data;
  wire[43:0] dpath_io_dmem_req_bits_addr;
  wire ctrl_io_dmem_req_bits_phys;
  wire[2:0] ctrl_io_dmem_req_bits_typ;
  wire ctrl_io_dmem_req_bits_kill;
  wire ctrl_io_dmem_req_valid;
  wire ctrl_io_imem_invalidate;
  wire ctrl_io_imem_btb_update_bits_incorrectTarget;
  wire ctrl_io_imem_btb_update_bits_isReturn;
  wire ctrl_io_imem_btb_update_bits_isCall;
  wire ctrl_io_imem_btb_update_bits_isJump;
  wire ctrl_io_imem_btb_update_bits_taken;
  wire[42:0] dpath_io_imem_btb_update_bits_returnAddr;
  wire[42:0] dpath_io_imem_btb_update_bits_target;
  wire[42:0] dpath_io_imem_btb_update_bits_pc;
  wire[1:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[3:0] ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[2:0] ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  wire[42:0] ctrl_io_imem_btb_update_bits_prediction_bits_target;
  wire ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  wire ctrl_io_imem_btb_update_bits_prediction_valid;
  wire ctrl_io_imem_btb_update_valid;
  wire ctrl_io_imem_resp_ready;
  wire[43:0] dpath_io_imem_req_bits_pc;
  wire ctrl_io_imem_req_valid;
  wire dpath_io_host_debug_stats_pcr;
  wire dpath_io_host_ipi_rep_ready;
  wire dpath_io_host_ipi_req_bits;
  wire dpath_io_host_ipi_req_valid;
  wire[63:0] dpath_io_host_pcr_rep_bits;
  wire dpath_io_host_pcr_rep_valid;
  wire dpath_io_host_pcr_req_ready;


  assign io_rocc_exception = ctrl_io_rocc_exception;
  assign io_rocc_s = ctrl_io_rocc_s;
  assign io_rocc_cmd_bits_rs2 = dpath_io_rocc_cmd_bits_rs2;
  assign io_rocc_cmd_bits_rs1 = dpath_io_rocc_cmd_bits_rs1;
  assign io_rocc_cmd_bits_inst_opcode = dpath_io_rocc_cmd_bits_inst_opcode;
  assign io_rocc_cmd_bits_inst_rd = dpath_io_rocc_cmd_bits_inst_rd;
  assign io_rocc_cmd_bits_inst_xs2 = dpath_io_rocc_cmd_bits_inst_xs2;
  assign io_rocc_cmd_bits_inst_xs1 = dpath_io_rocc_cmd_bits_inst_xs1;
  assign io_rocc_cmd_bits_inst_xd = dpath_io_rocc_cmd_bits_inst_xd;
  assign io_rocc_cmd_bits_inst_rs1 = dpath_io_rocc_cmd_bits_inst_rs1;
  assign io_rocc_cmd_bits_inst_rs2 = dpath_io_rocc_cmd_bits_inst_rs2;
  assign io_rocc_cmd_bits_inst_funct = dpath_io_rocc_cmd_bits_inst_funct;
  assign io_rocc_cmd_valid = ctrl_io_rocc_cmd_valid;
  assign io_ptw_status_s = dpath_io_ptw_status_s;
  assign io_ptw_status_ps = dpath_io_ptw_status_ps;
  assign io_ptw_status_ei = dpath_io_ptw_status_ei;
  assign io_ptw_status_pei = dpath_io_ptw_status_pei;
  assign io_ptw_status_ef = dpath_io_ptw_status_ef;
  assign io_ptw_status_u64 = dpath_io_ptw_status_u64;
  assign io_ptw_status_s64 = dpath_io_ptw_status_s64;
  assign io_ptw_status_vm = dpath_io_ptw_status_vm;
  assign io_ptw_status_er = dpath_io_ptw_status_er;
  assign io_ptw_status_zero = dpath_io_ptw_status_zero;
  assign io_ptw_status_im = dpath_io_ptw_status_im;
  assign io_ptw_status_ip = dpath_io_ptw_status_ip;
  assign io_ptw_sret = dpath_io_ptw_sret;
  assign io_ptw_invalidate = dpath_io_ptw_invalidate;
  assign io_ptw_ptbr = dpath_io_ptw_ptbr;
  assign io_dmem_req_bits_cmd = ctrl_io_dmem_req_bits_cmd;
  assign io_dmem_req_bits_tag = dpath_io_dmem_req_bits_tag;
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data;
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr;
  assign io_dmem_req_bits_phys = ctrl_io_dmem_req_bits_phys;
  assign io_dmem_req_bits_typ = ctrl_io_dmem_req_bits_typ;
  assign io_dmem_req_bits_kill = ctrl_io_dmem_req_bits_kill;
  assign io_dmem_req_valid = ctrl_io_dmem_req_valid;
  assign io_imem_invalidate = ctrl_io_imem_invalidate;
  assign io_imem_btb_update_bits_incorrectTarget = ctrl_io_imem_btb_update_bits_incorrectTarget;
  assign io_imem_btb_update_bits_isReturn = ctrl_io_imem_btb_update_bits_isReturn;
  assign io_imem_btb_update_bits_isCall = ctrl_io_imem_btb_update_bits_isCall;
  assign io_imem_btb_update_bits_isJump = ctrl_io_imem_btb_update_bits_isJump;
  assign io_imem_btb_update_bits_taken = ctrl_io_imem_btb_update_bits_taken;
  assign io_imem_btb_update_bits_returnAddr = dpath_io_imem_btb_update_bits_returnAddr;
  assign io_imem_btb_update_bits_target = dpath_io_imem_btb_update_bits_target;
  assign io_imem_btb_update_bits_pc = dpath_io_imem_btb_update_bits_pc;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = ctrl_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_btb_update_bits_prediction_bits_bht_index = ctrl_io_imem_btb_update_bits_prediction_bits_bht_index;
  assign io_imem_btb_update_bits_prediction_bits_entry = ctrl_io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_btb_update_bits_prediction_bits_target = ctrl_io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_btb_update_bits_prediction_bits_taken = ctrl_io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_btb_update_bits_prediction_valid = ctrl_io_imem_btb_update_bits_prediction_valid;
  assign io_imem_btb_update_valid = ctrl_io_imem_btb_update_valid;
  assign io_imem_resp_ready = ctrl_io_imem_resp_ready;
  assign io_imem_req_bits_pc = dpath_io_imem_req_bits_pc;
  assign io_imem_req_valid = ctrl_io_imem_req_valid;
  assign io_host_debug_stats_pcr = dpath_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = dpath_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = dpath_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = dpath_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = dpath_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = dpath_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = dpath_io_host_pcr_req_ready;
  Control ctrl(.clk(clk), .reset(reset),
       .io_dpath_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_dpath_killd( ctrl_io_dpath_killd ),
       .io_dpath_ren_1( ctrl_io_dpath_ren_1 ),
       .io_dpath_ren_0( ctrl_io_dpath_ren_0 ),
       .io_dpath_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_dpath_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_dpath_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_dpath_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_dpath_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_dpath_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_dpath_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_dpath_div_val(  )
       //.io_dpath_div_kill(  )
       .io_dpath_csr( ctrl_io_dpath_csr ),
       .io_dpath_sret( ctrl_io_dpath_sret ),
       .io_dpath_mem_load( ctrl_io_dpath_mem_load ),
       .io_dpath_wb_load( ctrl_io_dpath_wb_load ),
       .io_dpath_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_dpath_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_dpath_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_dpath_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_dpath_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_dpath_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_dpath_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_dpath_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_dpath_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_dpath_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_dpath_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_dpath_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_dpath_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_dpath_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_dpath_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_dpath_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_dpath_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_dpath_retire( ctrl_io_dpath_retire ),
       .io_dpath_exception( ctrl_io_dpath_exception ),
       .io_dpath_cause( ctrl_io_dpath_cause ),
       .io_dpath_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_dpath_inst( dpath_io_ctrl_inst ),
       //.io_dpath_jalr_eq(  )
       .io_dpath_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_dpath_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_dpath_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_dpath_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_dpath_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_dpath_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_dpath_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_dpath_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_dpath_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_dpath_status_ip( dpath_io_ctrl_status_ip ),
       .io_dpath_status_im( dpath_io_ctrl_status_im ),
       .io_dpath_status_zero( dpath_io_ctrl_status_zero ),
       .io_dpath_status_er( dpath_io_ctrl_status_er ),
       .io_dpath_status_vm( dpath_io_ctrl_status_vm ),
       .io_dpath_status_s64( dpath_io_ctrl_status_s64 ),
       .io_dpath_status_u64( dpath_io_ctrl_status_u64 ),
       .io_dpath_status_ef( dpath_io_ctrl_status_ef ),
       .io_dpath_status_pei( dpath_io_ctrl_status_pei ),
       .io_dpath_status_ei( dpath_io_ctrl_status_ei ),
       .io_dpath_status_ps( dpath_io_ctrl_status_ps ),
       .io_dpath_status_s( dpath_io_ctrl_status_s ),
       .io_dpath_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_dpath_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_dpath_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_imem_req_valid( ctrl_io_imem_req_valid ),
       //.io_imem_req_bits_pc(  )
       .io_imem_resp_ready( ctrl_io_imem_resp_ready ),
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( ctrl_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( ctrl_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( ctrl_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( ctrl_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( ctrl_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( ctrl_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( ctrl_io_imem_btb_update_bits_prediction_bits_bht_value ),
       //.io_imem_btb_update_bits_pc(  )
       //.io_imem_btb_update_bits_target(  )
       //.io_imem_btb_update_bits_returnAddr(  )
       .io_imem_btb_update_bits_taken( ctrl_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( ctrl_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( ctrl_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( ctrl_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( ctrl_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( ctrl_io_imem_invalidate ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       .io_dmem_req_valid( ctrl_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( ctrl_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( ctrl_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( ctrl_io_dmem_req_bits_phys ),
       //.io_dmem_req_bits_addr(  )
       //.io_dmem_req_bits_data(  )
       //.io_dmem_req_bits_tag(  )
       .io_dmem_req_bits_cmd( ctrl_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_fpu_valid( ctrl_io_fpu_valid ),
       .io_fpu_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_fpu_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_fpu_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_fpu_killx( ctrl_io_fpu_killx ),
       .io_fpu_killm( ctrl_io_fpu_killm ),
       .io_fpu_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_fpu_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_fpu_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_fpu_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_fpu_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_fpu_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_fpu_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_fpu_dec_single( FPU_io_ctrl_dec_single ),
       .io_fpu_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_fpu_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_fpu_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_fpu_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_fpu_dec_round( FPU_io_ctrl_dec_round ),
       .io_fpu_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_fpu_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_fpu_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       .io_rocc_cmd_valid( ctrl_io_rocc_cmd_valid ),
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       .io_rocc_s( ctrl_io_rocc_s ),
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits ),
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       .io_rocc_exception( ctrl_io_rocc_exception )
  );
  Datapath dpath(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( dpath_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( dpath_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( dpath_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( dpath_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( dpath_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( dpath_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( dpath_io_host_debug_stats_pcr ),
       .io_ctrl_sel_pc( ctrl_io_dpath_sel_pc ),
       .io_ctrl_killd( ctrl_io_dpath_killd ),
       .io_ctrl_ren_1( ctrl_io_dpath_ren_1 ),
       .io_ctrl_ren_0( ctrl_io_dpath_ren_0 ),
       .io_ctrl_sel_alu2( ctrl_io_dpath_sel_alu2 ),
       .io_ctrl_sel_alu1( ctrl_io_dpath_sel_alu1 ),
       .io_ctrl_sel_imm( ctrl_io_dpath_sel_imm ),
       .io_ctrl_fn_dw( ctrl_io_dpath_fn_dw ),
       .io_ctrl_fn_alu( ctrl_io_dpath_fn_alu ),
       .io_ctrl_div_mul_val( ctrl_io_dpath_div_mul_val ),
       .io_ctrl_div_mul_kill( ctrl_io_dpath_div_mul_kill ),
       //.io_ctrl_div_val(  )
       //.io_ctrl_div_kill(  )
       .io_ctrl_csr( ctrl_io_dpath_csr ),
       .io_ctrl_sret( ctrl_io_dpath_sret ),
       .io_ctrl_mem_load( ctrl_io_dpath_mem_load ),
       .io_ctrl_wb_load( ctrl_io_dpath_wb_load ),
       .io_ctrl_ex_fp_val( ctrl_io_dpath_ex_fp_val ),
       .io_ctrl_mem_fp_val( ctrl_io_dpath_mem_fp_val ),
       .io_ctrl_ex_wen( ctrl_io_dpath_ex_wen ),
       .io_ctrl_ex_valid( ctrl_io_dpath_ex_valid ),
       .io_ctrl_mem_jalr( ctrl_io_dpath_mem_jalr ),
       .io_ctrl_mem_branch( ctrl_io_dpath_mem_branch ),
       .io_ctrl_mem_wen( ctrl_io_dpath_mem_wen ),
       .io_ctrl_wb_wen( ctrl_io_dpath_wb_wen ),
       .io_ctrl_ex_mem_type( ctrl_io_dpath_ex_mem_type ),
       .io_ctrl_ex_rs2_val( ctrl_io_dpath_ex_rs2_val ),
       .io_ctrl_ex_rocc_val( ctrl_io_dpath_ex_rocc_val ),
       .io_ctrl_mem_rocc_val( ctrl_io_dpath_mem_rocc_val ),
       .io_ctrl_bypass_1( ctrl_io_dpath_bypass_1 ),
       .io_ctrl_bypass_0( ctrl_io_dpath_bypass_0 ),
       .io_ctrl_bypass_src_1( ctrl_io_dpath_bypass_src_1 ),
       .io_ctrl_bypass_src_0( ctrl_io_dpath_bypass_src_0 ),
       .io_ctrl_ll_ready( ctrl_io_dpath_ll_ready ),
       .io_ctrl_retire( ctrl_io_dpath_retire ),
       .io_ctrl_exception( ctrl_io_dpath_exception ),
       .io_ctrl_cause( ctrl_io_dpath_cause ),
       .io_ctrl_badvaddr_wen( ctrl_io_dpath_badvaddr_wen ),
       .io_ctrl_inst( dpath_io_ctrl_inst ),
       //.io_ctrl_jalr_eq(  )
       .io_ctrl_mem_br_taken( dpath_io_ctrl_mem_br_taken ),
       .io_ctrl_mem_misprediction( dpath_io_ctrl_mem_misprediction ),
       .io_ctrl_div_mul_rdy( dpath_io_ctrl_div_mul_rdy ),
       .io_ctrl_ll_wen( dpath_io_ctrl_ll_wen ),
       .io_ctrl_ll_waddr( dpath_io_ctrl_ll_waddr ),
       .io_ctrl_ex_waddr( dpath_io_ctrl_ex_waddr ),
       .io_ctrl_mem_rs1_ra( dpath_io_ctrl_mem_rs1_ra ),
       .io_ctrl_mem_waddr( dpath_io_ctrl_mem_waddr ),
       .io_ctrl_wb_waddr( dpath_io_ctrl_wb_waddr ),
       .io_ctrl_status_ip( dpath_io_ctrl_status_ip ),
       .io_ctrl_status_im( dpath_io_ctrl_status_im ),
       .io_ctrl_status_zero( dpath_io_ctrl_status_zero ),
       .io_ctrl_status_er( dpath_io_ctrl_status_er ),
       .io_ctrl_status_vm( dpath_io_ctrl_status_vm ),
       .io_ctrl_status_s64( dpath_io_ctrl_status_s64 ),
       .io_ctrl_status_u64( dpath_io_ctrl_status_u64 ),
       .io_ctrl_status_ef( dpath_io_ctrl_status_ef ),
       .io_ctrl_status_pei( dpath_io_ctrl_status_pei ),
       .io_ctrl_status_ei( dpath_io_ctrl_status_ei ),
       .io_ctrl_status_ps( dpath_io_ctrl_status_ps ),
       .io_ctrl_status_s( dpath_io_ctrl_status_s ),
       .io_ctrl_fp_sboard_clr( dpath_io_ctrl_fp_sboard_clr ),
       .io_ctrl_fp_sboard_clra( dpath_io_ctrl_fp_sboard_clra ),
       .io_ctrl_csr_replay( dpath_io_ctrl_csr_replay ),
       .io_dmem_req_ready( io_dmem_req_ready ),
       //.io_dmem_req_valid(  )
       //.io_dmem_req_bits_kill(  )
       //.io_dmem_req_bits_typ(  )
       //.io_dmem_req_bits_phys(  )
       .io_dmem_req_bits_addr( dpath_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( dpath_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( dpath_io_dmem_req_bits_tag ),
       //.io_dmem_req_bits_cmd(  )
       .io_dmem_resp_valid( io_dmem_resp_valid ),
       .io_dmem_resp_bits_nack( io_dmem_resp_bits_nack ),
       .io_dmem_resp_bits_replay( io_dmem_resp_bits_replay ),
       .io_dmem_resp_bits_typ( io_dmem_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( io_dmem_resp_bits_has_data ),
       .io_dmem_resp_bits_data( io_dmem_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( io_dmem_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( io_dmem_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( io_dmem_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( io_dmem_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( io_dmem_resp_bits_store_data ),
       .io_dmem_replay_next_valid( io_dmem_replay_next_valid ),
       .io_dmem_replay_next_bits( io_dmem_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( io_dmem_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( io_dmem_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( io_dmem_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( io_dmem_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       .io_dmem_ptw_req_valid( io_dmem_ptw_req_valid ),
       .io_dmem_ptw_req_bits( io_dmem_ptw_req_bits ),
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( io_dmem_ordered ),
       .io_ptw_ptbr( dpath_io_ptw_ptbr ),
       .io_ptw_invalidate( dpath_io_ptw_invalidate ),
       .io_ptw_sret( dpath_io_ptw_sret ),
       .io_ptw_status_ip( dpath_io_ptw_status_ip ),
       .io_ptw_status_im( dpath_io_ptw_status_im ),
       .io_ptw_status_zero( dpath_io_ptw_status_zero ),
       .io_ptw_status_er( dpath_io_ptw_status_er ),
       .io_ptw_status_vm( dpath_io_ptw_status_vm ),
       .io_ptw_status_s64( dpath_io_ptw_status_s64 ),
       .io_ptw_status_u64( dpath_io_ptw_status_u64 ),
       .io_ptw_status_ef( dpath_io_ptw_status_ef ),
       .io_ptw_status_pei( dpath_io_ptw_status_pei ),
       .io_ptw_status_ei( dpath_io_ptw_status_ei ),
       .io_ptw_status_ps( dpath_io_ptw_status_ps ),
       .io_ptw_status_s( dpath_io_ptw_status_s ),
       //.io_imem_req_valid(  )
       .io_imem_req_bits_pc( dpath_io_imem_req_bits_pc ),
       //.io_imem_resp_ready(  )
       .io_imem_resp_valid( io_imem_resp_valid ),
       .io_imem_resp_bits_pc( io_imem_resp_bits_pc ),
       .io_imem_resp_bits_data( io_imem_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( io_imem_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( io_imem_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( io_imem_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( io_imem_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( io_imem_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( io_imem_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( io_imem_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( io_imem_btb_resp_bits_bht_value ),
       //.io_imem_btb_update_valid(  )
       //.io_imem_btb_update_bits_prediction_valid(  )
       //.io_imem_btb_update_bits_prediction_bits_taken(  )
       //.io_imem_btb_update_bits_prediction_bits_target(  )
       //.io_imem_btb_update_bits_prediction_bits_entry(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_index(  )
       //.io_imem_btb_update_bits_prediction_bits_bht_value(  )
       .io_imem_btb_update_bits_pc( dpath_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( dpath_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( dpath_io_imem_btb_update_bits_returnAddr ),
       //.io_imem_btb_update_bits_taken(  )
       //.io_imem_btb_update_bits_isJump(  )
       //.io_imem_btb_update_bits_isCall(  )
       //.io_imem_btb_update_bits_isReturn(  )
       //.io_imem_btb_update_bits_incorrectTarget(  )
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( io_imem_ptw_req_valid ),
       .io_imem_ptw_req_bits( io_imem_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       //.io_imem_invalidate(  )
       .io_fpu_inst( dpath_io_fpu_inst ),
       .io_fpu_fromint_data( dpath_io_fpu_fromint_data ),
       .io_fpu_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_fpu_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_fpu_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_fpu_store_data( FPU_io_dpath_store_data ),
       .io_fpu_toint_data( FPU_io_dpath_toint_data ),
       .io_fpu_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_fpu_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_fpu_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_fpu_dmem_resp_data( dpath_io_fpu_dmem_resp_data ),
       .io_rocc_cmd_ready( io_rocc_cmd_ready ),
       //.io_rocc_cmd_valid(  )
       .io_rocc_cmd_bits_inst_funct( dpath_io_rocc_cmd_bits_inst_funct ),
       .io_rocc_cmd_bits_inst_rs2( dpath_io_rocc_cmd_bits_inst_rs2 ),
       .io_rocc_cmd_bits_inst_rs1( dpath_io_rocc_cmd_bits_inst_rs1 ),
       .io_rocc_cmd_bits_inst_xd( dpath_io_rocc_cmd_bits_inst_xd ),
       .io_rocc_cmd_bits_inst_xs1( dpath_io_rocc_cmd_bits_inst_xs1 ),
       .io_rocc_cmd_bits_inst_xs2( dpath_io_rocc_cmd_bits_inst_xs2 ),
       .io_rocc_cmd_bits_inst_rd( dpath_io_rocc_cmd_bits_inst_rd ),
       .io_rocc_cmd_bits_inst_opcode( dpath_io_rocc_cmd_bits_inst_opcode ),
       .io_rocc_cmd_bits_rs1( dpath_io_rocc_cmd_bits_rs1 ),
       .io_rocc_cmd_bits_rs2( dpath_io_rocc_cmd_bits_rs2 ),
       //.io_rocc_resp_ready(  )
       .io_rocc_resp_valid( io_rocc_resp_valid ),
       .io_rocc_resp_bits_rd( io_rocc_resp_bits_rd ),
       .io_rocc_resp_bits_data( io_rocc_resp_bits_data ),
       //.io_rocc_mem_req_ready(  )
       .io_rocc_mem_req_valid( io_rocc_mem_req_valid ),
       .io_rocc_mem_req_bits_kill( io_rocc_mem_req_bits_kill ),
       .io_rocc_mem_req_bits_typ( io_rocc_mem_req_bits_typ ),
       .io_rocc_mem_req_bits_phys( io_rocc_mem_req_bits_phys ),
       .io_rocc_mem_req_bits_addr( io_rocc_mem_req_bits_addr ),
       .io_rocc_mem_req_bits_data( io_rocc_mem_req_bits_data ),
       .io_rocc_mem_req_bits_tag( io_rocc_mem_req_bits_tag ),
       .io_rocc_mem_req_bits_cmd( io_rocc_mem_req_bits_cmd ),
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       .io_rocc_mem_ptw_req_ready( io_rocc_mem_ptw_req_ready ),
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       .io_rocc_mem_ptw_resp_valid( io_rocc_mem_ptw_resp_valid ),
       .io_rocc_mem_ptw_resp_bits_error( io_rocc_mem_ptw_resp_bits_error ),
       .io_rocc_mem_ptw_resp_bits_ppn( io_rocc_mem_ptw_resp_bits_ppn ),
       .io_rocc_mem_ptw_resp_bits_perm( io_rocc_mem_ptw_resp_bits_perm ),
       .io_rocc_mem_ptw_status_ip( io_rocc_mem_ptw_status_ip ),
       .io_rocc_mem_ptw_status_im( io_rocc_mem_ptw_status_im ),
       .io_rocc_mem_ptw_status_zero( io_rocc_mem_ptw_status_zero ),
       .io_rocc_mem_ptw_status_er( io_rocc_mem_ptw_status_er ),
       .io_rocc_mem_ptw_status_vm( io_rocc_mem_ptw_status_vm ),
       .io_rocc_mem_ptw_status_s64( io_rocc_mem_ptw_status_s64 ),
       .io_rocc_mem_ptw_status_u64( io_rocc_mem_ptw_status_u64 ),
       .io_rocc_mem_ptw_status_ef( io_rocc_mem_ptw_status_ef ),
       .io_rocc_mem_ptw_status_pei( io_rocc_mem_ptw_status_pei ),
       .io_rocc_mem_ptw_status_ei( io_rocc_mem_ptw_status_ei ),
       .io_rocc_mem_ptw_status_ps( io_rocc_mem_ptw_status_ps ),
       .io_rocc_mem_ptw_status_s( io_rocc_mem_ptw_status_s ),
       .io_rocc_mem_ptw_invalidate( io_rocc_mem_ptw_invalidate ),
       .io_rocc_mem_ptw_sret( io_rocc_mem_ptw_sret ),
       //.io_rocc_mem_ordered(  )
       .io_rocc_busy( io_rocc_busy ),
       //.io_rocc_s(  )
       .io_rocc_interrupt( io_rocc_interrupt ),
       //.io_rocc_imem_acquire_ready(  )
       .io_rocc_imem_acquire_valid( io_rocc_imem_acquire_valid ),
       .io_rocc_imem_acquire_bits_header_src( io_rocc_imem_acquire_bits_header_src ),
       .io_rocc_imem_acquire_bits_header_dst( io_rocc_imem_acquire_bits_header_dst ),
       .io_rocc_imem_acquire_bits_payload_addr( io_rocc_imem_acquire_bits_payload_addr ),
       .io_rocc_imem_acquire_bits_payload_client_xact_id( io_rocc_imem_acquire_bits_payload_client_xact_id ),
       .io_rocc_imem_acquire_bits_payload_data( io_rocc_imem_acquire_bits_payload_data ),
       .io_rocc_imem_acquire_bits_payload_a_type( io_rocc_imem_acquire_bits_payload_a_type ),
       .io_rocc_imem_acquire_bits_payload_write_mask( io_rocc_imem_acquire_bits_payload_write_mask ),
       .io_rocc_imem_acquire_bits_payload_subword_addr( io_rocc_imem_acquire_bits_payload_subword_addr ),
       .io_rocc_imem_acquire_bits_payload_atomic_opcode( io_rocc_imem_acquire_bits_payload_atomic_opcode ),
       .io_rocc_imem_grant_ready( io_rocc_imem_grant_ready ),
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       .io_rocc_imem_finish_valid( io_rocc_imem_finish_valid ),
       .io_rocc_imem_finish_bits_header_src( io_rocc_imem_finish_bits_header_src ),
       .io_rocc_imem_finish_bits_header_dst( io_rocc_imem_finish_bits_header_dst ),
       .io_rocc_imem_finish_bits_payload_master_xact_id( io_rocc_imem_finish_bits_payload_master_xact_id ),
       //.io_rocc_iptw_req_ready(  )
       .io_rocc_iptw_req_valid( io_rocc_iptw_req_valid ),
       .io_rocc_iptw_req_bits( io_rocc_iptw_req_bits ),
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       .io_rocc_dptw_req_valid( io_rocc_dptw_req_valid ),
       .io_rocc_dptw_req_bits( io_rocc_dptw_req_bits ),
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       .io_rocc_pptw_req_valid( io_rocc_pptw_req_valid ),
       .io_rocc_pptw_req_bits( io_rocc_pptw_req_bits )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  FPU FPU(.clk(clk), .reset(reset),
       .io_ctrl_valid( ctrl_io_fpu_valid ),
       .io_ctrl_fcsr_rdy( FPU_io_ctrl_fcsr_rdy ),
       .io_ctrl_nack_mem( FPU_io_ctrl_nack_mem ),
       .io_ctrl_illegal_rm( FPU_io_ctrl_illegal_rm ),
       .io_ctrl_killx( ctrl_io_fpu_killx ),
       .io_ctrl_killm( ctrl_io_fpu_killm ),
       .io_ctrl_dec_cmd( FPU_io_ctrl_dec_cmd ),
       .io_ctrl_dec_ldst( FPU_io_ctrl_dec_ldst ),
       .io_ctrl_dec_wen( FPU_io_ctrl_dec_wen ),
       .io_ctrl_dec_ren1( FPU_io_ctrl_dec_ren1 ),
       .io_ctrl_dec_ren2( FPU_io_ctrl_dec_ren2 ),
       .io_ctrl_dec_ren3( FPU_io_ctrl_dec_ren3 ),
       .io_ctrl_dec_swap23( FPU_io_ctrl_dec_swap23 ),
       .io_ctrl_dec_single( FPU_io_ctrl_dec_single ),
       .io_ctrl_dec_fromint( FPU_io_ctrl_dec_fromint ),
       .io_ctrl_dec_toint( FPU_io_ctrl_dec_toint ),
       .io_ctrl_dec_fastpipe( FPU_io_ctrl_dec_fastpipe ),
       .io_ctrl_dec_fma( FPU_io_ctrl_dec_fma ),
       .io_ctrl_dec_round( FPU_io_ctrl_dec_round ),
       .io_ctrl_sboard_set( FPU_io_ctrl_sboard_set ),
       .io_ctrl_sboard_clr( FPU_io_ctrl_sboard_clr ),
       .io_ctrl_sboard_clra( FPU_io_ctrl_sboard_clra ),
       .io_dpath_inst( dpath_io_fpu_inst ),
       .io_dpath_fromint_data( dpath_io_fpu_fromint_data ),
       .io_dpath_fcsr_rm( dpath_io_fpu_fcsr_rm ),
       .io_dpath_fcsr_flags_valid( FPU_io_dpath_fcsr_flags_valid ),
       .io_dpath_fcsr_flags_bits( FPU_io_dpath_fcsr_flags_bits ),
       .io_dpath_store_data( FPU_io_dpath_store_data ),
       .io_dpath_toint_data( FPU_io_dpath_toint_data ),
       .io_dpath_dmem_resp_val( dpath_io_fpu_dmem_resp_val ),
       .io_dpath_dmem_resp_type( dpath_io_fpu_dmem_resp_type ),
       .io_dpath_dmem_resp_tag( dpath_io_fpu_dmem_resp_tag ),
       .io_dpath_dmem_resp_data( dpath_io_fpu_dmem_resp_data )
  );
endmodule

module HellaCacheArbiter(input clk,
    output io_requestor_1_req_ready,
    input  io_requestor_1_req_valid,
    input  io_requestor_1_req_bits_kill,
    input [2:0] io_requestor_1_req_bits_typ,
    input  io_requestor_1_req_bits_phys,
    input [43:0] io_requestor_1_req_bits_addr,
    input [63:0] io_requestor_1_req_bits_data,
    input [7:0] io_requestor_1_req_bits_tag,
    input [4:0] io_requestor_1_req_bits_cmd,
    output io_requestor_1_resp_valid,
    output io_requestor_1_resp_bits_nack,
    output io_requestor_1_resp_bits_replay,
    output[2:0] io_requestor_1_resp_bits_typ,
    output io_requestor_1_resp_bits_has_data,
    output[63:0] io_requestor_1_resp_bits_data,
    output[63:0] io_requestor_1_resp_bits_data_subword,
    output[7:0] io_requestor_1_resp_bits_tag,
    output[3:0] io_requestor_1_resp_bits_cmd,
    output[43:0] io_requestor_1_resp_bits_addr,
    output[63:0] io_requestor_1_resp_bits_store_data,
    output io_requestor_1_replay_next_valid,
    output[7:0] io_requestor_1_replay_next_bits,
    output io_requestor_1_xcpt_ma_ld,
    output io_requestor_1_xcpt_ma_st,
    output io_requestor_1_xcpt_pf_ld,
    output io_requestor_1_xcpt_pf_st,
    //input  io_requestor_1_ptw_req_ready
    //output io_requestor_1_ptw_req_valid
    //output[29:0] io_requestor_1_ptw_req_bits
    //input  io_requestor_1_ptw_resp_valid
    //input  io_requestor_1_ptw_resp_bits_error
    //input [18:0] io_requestor_1_ptw_resp_bits_ppn
    //input [5:0] io_requestor_1_ptw_resp_bits_perm
    //input [7:0] io_requestor_1_ptw_status_ip
    //input [7:0] io_requestor_1_ptw_status_im
    //input [6:0] io_requestor_1_ptw_status_zero
    //input  io_requestor_1_ptw_status_er
    //input  io_requestor_1_ptw_status_vm
    //input  io_requestor_1_ptw_status_s64
    //input  io_requestor_1_ptw_status_u64
    //input  io_requestor_1_ptw_status_ef
    //input  io_requestor_1_ptw_status_pei
    //input  io_requestor_1_ptw_status_ei
    //input  io_requestor_1_ptw_status_ps
    //input  io_requestor_1_ptw_status_s
    //input  io_requestor_1_ptw_invalidate
    //input  io_requestor_1_ptw_sret
    output io_requestor_1_ordered,
    output io_requestor_0_req_ready,
    input  io_requestor_0_req_valid,
    input  io_requestor_0_req_bits_kill,
    input [2:0] io_requestor_0_req_bits_typ,
    input  io_requestor_0_req_bits_phys,
    input [43:0] io_requestor_0_req_bits_addr,
    input [63:0] io_requestor_0_req_bits_data,
    input [7:0] io_requestor_0_req_bits_tag,
    input [4:0] io_requestor_0_req_bits_cmd,
    output io_requestor_0_resp_valid,
    output io_requestor_0_resp_bits_nack,
    output io_requestor_0_resp_bits_replay,
    output[2:0] io_requestor_0_resp_bits_typ,
    output io_requestor_0_resp_bits_has_data,
    output[63:0] io_requestor_0_resp_bits_data,
    output[63:0] io_requestor_0_resp_bits_data_subword,
    output[7:0] io_requestor_0_resp_bits_tag,
    output[3:0] io_requestor_0_resp_bits_cmd,
    output[43:0] io_requestor_0_resp_bits_addr,
    output[63:0] io_requestor_0_resp_bits_store_data,
    output io_requestor_0_replay_next_valid,
    output[7:0] io_requestor_0_replay_next_bits,
    output io_requestor_0_xcpt_ma_ld,
    output io_requestor_0_xcpt_ma_st,
    output io_requestor_0_xcpt_pf_ld,
    output io_requestor_0_xcpt_pf_st,
    //input  io_requestor_0_ptw_req_ready
    //output io_requestor_0_ptw_req_valid
    //output[29:0] io_requestor_0_ptw_req_bits
    //input  io_requestor_0_ptw_resp_valid
    //input  io_requestor_0_ptw_resp_bits_error
    //input [18:0] io_requestor_0_ptw_resp_bits_ppn
    //input [5:0] io_requestor_0_ptw_resp_bits_perm
    //input [7:0] io_requestor_0_ptw_status_ip
    //input [7:0] io_requestor_0_ptw_status_im
    //input [6:0] io_requestor_0_ptw_status_zero
    //input  io_requestor_0_ptw_status_er
    //input  io_requestor_0_ptw_status_vm
    //input  io_requestor_0_ptw_status_s64
    //input  io_requestor_0_ptw_status_u64
    //input  io_requestor_0_ptw_status_ef
    //input  io_requestor_0_ptw_status_pei
    //input  io_requestor_0_ptw_status_ei
    //input  io_requestor_0_ptw_status_ps
    //input  io_requestor_0_ptw_status_s
    //input  io_requestor_0_ptw_invalidate
    //input  io_requestor_0_ptw_sret
    output io_requestor_0_ordered,
    input  io_mem_req_ready,
    output io_mem_req_valid,
    output io_mem_req_bits_kill,
    output[2:0] io_mem_req_bits_typ,
    output io_mem_req_bits_phys,
    output[43:0] io_mem_req_bits_addr,
    output[63:0] io_mem_req_bits_data,
    output[7:0] io_mem_req_bits_tag,
    output[4:0] io_mem_req_bits_cmd,
    input  io_mem_resp_valid,
    input  io_mem_resp_bits_nack,
    input  io_mem_resp_bits_replay,
    input [2:0] io_mem_resp_bits_typ,
    input  io_mem_resp_bits_has_data,
    input [63:0] io_mem_resp_bits_data,
    input [63:0] io_mem_resp_bits_data_subword,
    input [7:0] io_mem_resp_bits_tag,
    input [3:0] io_mem_resp_bits_cmd,
    input [43:0] io_mem_resp_bits_addr,
    input [63:0] io_mem_resp_bits_store_data,
    input  io_mem_replay_next_valid,
    input [7:0] io_mem_replay_next_bits,
    input  io_mem_xcpt_ma_ld,
    input  io_mem_xcpt_ma_st,
    input  io_mem_xcpt_pf_ld,
    input  io_mem_xcpt_pf_st,
    //output io_mem_ptw_req_ready
    input  io_mem_ptw_req_valid,
    input [29:0] io_mem_ptw_req_bits,
    //output io_mem_ptw_resp_valid
    //output io_mem_ptw_resp_bits_error
    //output[18:0] io_mem_ptw_resp_bits_ppn
    //output[5:0] io_mem_ptw_resp_bits_perm
    //output[7:0] io_mem_ptw_status_ip
    //output[7:0] io_mem_ptw_status_im
    //output[6:0] io_mem_ptw_status_zero
    //output io_mem_ptw_status_er
    //output io_mem_ptw_status_vm
    //output io_mem_ptw_status_s64
    //output io_mem_ptw_status_u64
    //output io_mem_ptw_status_ef
    //output io_mem_ptw_status_pei
    //output io_mem_ptw_status_ei
    //output io_mem_ptw_status_ps
    //output io_mem_ptw_status_s
    //output io_mem_ptw_invalidate
    //output io_mem_ptw_sret
    input  io_mem_ordered
);

  wire[4:0] T0;
  wire[7:0] T1;
  wire[8:0] T2;
  wire[8:0] T3;
  wire[8:0] T4;
  wire[63:0] T5;
  reg  r_valid_0;
  wire[43:0] T6;
  wire T7;
  wire[2:0] T8;
  wire T9;
  wire T10;
  wire[7:0] T11;
  wire[6:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire[7:0] T16;
  wire[6:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire[7:0] T23;
  wire[6:0] T24;
  wire T25;
  wire T26;
  wire T27;
  wire[7:0] T28;
  wire[6:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    r_valid_0 = {1{$random}};
  end
`endif

  assign io_mem_req_bits_cmd = T0;
  assign T0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign io_mem_req_bits_tag = T1;
  assign T1 = T2[3'h7:1'h0];
  assign T2 = io_requestor_0_req_valid ? T4 : T3;
  assign T3 = {io_requestor_1_req_bits_tag, 1'h1};
  assign T4 = {io_requestor_0_req_bits_tag, 1'h0};
  assign io_mem_req_bits_data = T5;
  assign T5 = r_valid_0 ? io_requestor_0_req_bits_data : io_requestor_1_req_bits_data;
  assign io_mem_req_bits_addr = T6;
  assign T6 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign io_mem_req_bits_phys = T7;
  assign T7 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign io_mem_req_bits_typ = T8;
  assign T8 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign io_mem_req_bits_kill = T9;
  assign T9 = r_valid_0 ? io_requestor_0_req_bits_kill : io_requestor_1_req_bits_kill;
  assign io_mem_req_valid = T10;
  assign T10 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_replay_next_bits = T11;
  assign T11 = {1'h0, T12};
  assign T12 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_0_replay_next_valid = T13;
  assign T13 = io_mem_replay_next_valid & T14;
  assign T14 = T15 == 1'h0;
  assign T15 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_tag = T16;
  assign T16 = {1'h0, T17};
  assign T17 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_0_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_replay = T18;
  assign T18 = io_mem_resp_bits_replay & T19;
  assign T19 = T20 == 1'h0;
  assign T20 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_0_resp_bits_nack = T21;
  assign T21 = io_mem_resp_bits_nack & T19;
  assign io_requestor_0_resp_valid = T22;
  assign T22 = io_mem_resp_valid & T19;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_replay_next_bits = T23;
  assign T23 = {1'h0, T24};
  assign T24 = io_mem_replay_next_bits >> 1'h1;
  assign io_requestor_1_replay_next_valid = T25;
  assign T25 = io_mem_replay_next_valid & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = io_mem_replay_next_bits[1'h0:1'h0];
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_tag = T28;
  assign T28 = {1'h0, T29};
  assign T29 = io_mem_resp_bits_tag >> 1'h1;
  assign io_requestor_1_resp_bits_data_subword = io_mem_resp_bits_data_subword;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_replay = T30;
  assign T30 = io_mem_resp_bits_replay & T31;
  assign T31 = T32 == 1'h1;
  assign T32 = io_mem_resp_bits_tag[1'h0:1'h0];
  assign io_requestor_1_resp_bits_nack = T33;
  assign T33 = io_mem_resp_bits_nack & T31;
  assign io_requestor_1_resp_valid = T34;
  assign T34 = io_mem_resp_valid & T31;
  assign io_requestor_1_req_ready = T35;
  assign T35 = io_requestor_0_req_ready & T36;
  assign T36 = io_requestor_0_req_valid ^ 1'h1;

  always @(posedge clk) begin
    r_valid_0 <= io_requestor_0_req_valid;
  end
endmodule

module RRArbiter_1(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[3:0] T9;
  wire T10;
  wire[2:0] T11;
  wire[5:0] T12;
  wire[2:0] T13;
  wire[511:0] T14;
  wire[1:0] T15;
  wire[25:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_atomic_opcode = T9;
  assign T9 = T10 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T10 = T0;
  assign io_out_bits_payload_subword_addr = T11;
  assign T11 = T10 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign io_out_bits_payload_write_mask = T12;
  assign T12 = T10 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign io_out_bits_payload_a_type = T13;
  assign T13 = T10 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign io_out_bits_payload_data = T14;
  assign T14 = T10 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign io_out_bits_payload_client_xact_id = T15;
  assign T15 = T10 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign io_out_bits_payload_addr = T16;
  assign T16 = T10 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign io_out_bits_header_dst = T17;
  assign T17 = T10 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T18;
  assign T18 = T10 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T19;
  assign T19 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T20;
  assign T20 = T21 & io_out_ready;
  assign T21 = T28 | T22;
  assign T22 = T23 ^ 1'h1;
  assign T23 = T26 | T24;
  assign T24 = io_in_1_valid & T25;
  assign T25 = R5 < 1'h1;
  assign T26 = io_in_0_valid & T27;
  assign T27 = R5 < 1'h0;
  assign T28 = R5 < 1'h0;
  assign io_in_1_ready = T29;
  assign T29 = T30 & io_out_ready;
  assign T30 = T34 | T31;
  assign T31 = T32 ^ 1'h1;
  assign T32 = T33 | io_in_0_valid;
  assign T33 = T26 | T24;
  assign T34 = T36 & T35;
  assign T35 = R5 < 1'h1;
  assign T36 = T26 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module RRArbiter_2(input clk, input reset,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output io_chosen
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire[2:0] T9;
  wire T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R5 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T3 ? 1'h1 : T2;
  assign T2 = io_in_0_valid == 1'h0;
  assign T3 = io_in_1_valid & T4;
  assign T4 = R5 < 1'h1;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = T8 ? T0 : R5;
  assign T8 = io_out_ready & io_out_valid;
  assign io_out_bits_payload_master_xact_id = T9;
  assign T9 = T10 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T10 = T0;
  assign io_out_bits_header_dst = T11;
  assign T11 = T10 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign io_out_bits_header_src = T12;
  assign T12 = T10 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign io_out_valid = T13;
  assign T13 = T10 ? io_in_1_valid : io_in_0_valid;
  assign io_in_0_ready = T14;
  assign T14 = T15 & io_out_ready;
  assign T15 = T22 | T16;
  assign T16 = T17 ^ 1'h1;
  assign T17 = T20 | T18;
  assign T18 = io_in_1_valid & T19;
  assign T19 = R5 < 1'h1;
  assign T20 = io_in_0_valid & T21;
  assign T21 = R5 < 1'h0;
  assign T22 = R5 < 1'h0;
  assign io_in_1_ready = T23;
  assign T23 = T24 & io_out_ready;
  assign T24 = T28 | T25;
  assign T25 = T26 ^ 1'h1;
  assign T26 = T27 | io_in_0_valid;
  assign T27 = T20 | T18;
  assign T28 = T30 & T29;
  assign T29 = R5 < 1'h1;
  assign T30 = T20 ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      R5 <= 1'h0;
    end else if(T8) begin
      R5 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatAppendsArbiterId(input clk, input reset,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire[1:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire[2:0] T3;
  wire[2:0] RRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire RRArbiter_1_io_out_valid;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[1:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire RRArbiter_0_io_out_valid;
  wire RRArbiter_1_io_in_0_ready;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_1_io_in_1_ready;
  wire[1:0] T15;
  wire T16;
  wire T17;
  wire RRArbiter_0_io_in_1_ready;


  assign T0 = T1[1'h1:1'h0];
  assign T1 = {io_in_0_acquire_bits_payload_client_xact_id, 1'h0};
  assign T2 = T3[1'h1:1'h0];
  assign T3 = {io_in_1_acquire_bits_payload_client_xact_id, 1'h1};
  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T4;
  assign T4 = T9 ? io_in_1_grant_ready : T5;
  assign T5 = T6 ? io_in_0_grant_ready : 1'h0;
  assign T6 = T7 == 1'h0;
  assign T7 = T8;
  assign T8 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign T9 = T10 == 1'h1;
  assign T10 = T11;
  assign T11 = io_out_grant_bits_payload_client_xact_id[1'h0:1'h0];
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = T12;
  assign T12 = {1'h0, T13};
  assign T13 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T14;
  assign T14 = T6 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = T15;
  assign T15 = {1'h0, T16};
  assign T16 = io_out_grant_bits_payload_client_xact_id >> 1'h1;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T17;
  assign T17 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  RRArbiter_1 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( T2 ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( T0 ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_2 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module Tile(input clk, input reset,
    input  io_tilelink_acquire_ready,
    output io_tilelink_acquire_valid,
    output[1:0] io_tilelink_acquire_bits_header_src,
    output[1:0] io_tilelink_acquire_bits_header_dst,
    output[25:0] io_tilelink_acquire_bits_payload_addr,
    output[1:0] io_tilelink_acquire_bits_payload_client_xact_id,
    output[511:0] io_tilelink_acquire_bits_payload_data,
    output[2:0] io_tilelink_acquire_bits_payload_a_type,
    output[5:0] io_tilelink_acquire_bits_payload_write_mask,
    output[2:0] io_tilelink_acquire_bits_payload_subword_addr,
    output[3:0] io_tilelink_acquire_bits_payload_atomic_opcode,
    output io_tilelink_grant_ready,
    input  io_tilelink_grant_valid,
    input [1:0] io_tilelink_grant_bits_header_src,
    input [1:0] io_tilelink_grant_bits_header_dst,
    input [511:0] io_tilelink_grant_bits_payload_data,
    input [1:0] io_tilelink_grant_bits_payload_client_xact_id,
    input [2:0] io_tilelink_grant_bits_payload_master_xact_id,
    input [3:0] io_tilelink_grant_bits_payload_g_type,
    input  io_tilelink_finish_ready,
    output io_tilelink_finish_valid,
    output[1:0] io_tilelink_finish_bits_header_src,
    output[1:0] io_tilelink_finish_bits_header_dst,
    output[2:0] io_tilelink_finish_bits_payload_master_xact_id,
    output io_tilelink_probe_ready,
    input  io_tilelink_probe_valid,
    input [1:0] io_tilelink_probe_bits_header_src,
    input [1:0] io_tilelink_probe_bits_header_dst,
    input [25:0] io_tilelink_probe_bits_payload_addr,
    input [2:0] io_tilelink_probe_bits_payload_master_xact_id,
    input [1:0] io_tilelink_probe_bits_payload_p_type,
    input  io_tilelink_release_ready,
    output io_tilelink_release_valid,
    output[1:0] io_tilelink_release_bits_header_src,
    output[1:0] io_tilelink_release_bits_header_dst,
    output[25:0] io_tilelink_release_bits_payload_addr,
    output[1:0] io_tilelink_release_bits_payload_client_xact_id,
    output[2:0] io_tilelink_release_bits_payload_master_xact_id,
    output[511:0] io_tilelink_release_bits_payload_data,
    output[2:0] io_tilelink_release_bits_payload_r_type,
    input  io_host_reset,
    input  io_host_id,
    output io_host_pcr_req_ready,
    input  io_host_pcr_req_valid,
    input  io_host_pcr_req_bits_rw,
    input [4:0] io_host_pcr_req_bits_addr,
    input [63:0] io_host_pcr_req_bits_data,
    input  io_host_pcr_rep_ready,
    output io_host_pcr_rep_valid,
    output[63:0] io_host_pcr_rep_bits,
    input  io_host_ipi_req_ready,
    output io_host_ipi_req_valid,
    output io_host_ipi_req_bits,
    output io_host_ipi_rep_ready,
    input  io_host_ipi_rep_valid,
    input  io_host_ipi_rep_bits,
    output io_host_debug_stats_pcr
);

  wire[2:0] dcache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] dcache_io_mem_finish_bits_header_dst;
  wire[1:0] dcache_io_mem_finish_bits_header_src;
  wire dcache_io_mem_finish_valid;
  wire dcache_io_mem_grant_ready;
  wire[3:0] dcache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] dcache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] dcache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] dcache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] dcache_io_mem_acquire_bits_payload_data;
  wire[1:0] dcache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] dcache_io_mem_acquire_bits_payload_addr;
  wire[1:0] dcache_io_mem_acquire_bits_header_dst;
  wire[1:0] dcache_io_mem_acquire_bits_header_src;
  wire dcache_io_mem_acquire_valid;
  wire[2:0] icache_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] icache_io_mem_finish_bits_header_dst;
  wire[1:0] icache_io_mem_finish_bits_header_src;
  wire icache_io_mem_finish_valid;
  wire icache_io_mem_grant_ready;
  wire[3:0] icache_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] icache_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] icache_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] icache_io_mem_acquire_bits_payload_a_type;
  wire[511:0] icache_io_mem_acquire_bits_payload_data;
  wire[1:0] icache_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] icache_io_mem_acquire_bits_payload_addr;
  wire icache_io_mem_acquire_valid;
  wire dcache_io_cpu_ordered;
  wire[29:0] dcache_io_cpu_ptw_req_bits;
  wire dcache_io_cpu_ptw_req_valid;
  wire dcache_io_cpu_xcpt_pf_st;
  wire dcache_io_cpu_xcpt_pf_ld;
  wire dcache_io_cpu_xcpt_ma_st;
  wire dcache_io_cpu_xcpt_ma_ld;
  wire[7:0] dcache_io_cpu_replay_next_bits;
  wire dcache_io_cpu_replay_next_valid;
  wire[63:0] dcache_io_cpu_resp_bits_store_data;
  wire[43:0] dcache_io_cpu_resp_bits_addr;
  wire[3:0] dcache_io_cpu_resp_bits_cmd;
  wire[7:0] dcache_io_cpu_resp_bits_tag;
  wire[63:0] dcache_io_cpu_resp_bits_data_subword;
  wire[63:0] dcache_io_cpu_resp_bits_data;
  wire dcache_io_cpu_resp_bits_has_data;
  wire[2:0] dcache_io_cpu_resp_bits_typ;
  wire dcache_io_cpu_resp_bits_replay;
  wire dcache_io_cpu_resp_bits_nack;
  wire dcache_io_cpu_resp_valid;
  wire dcache_io_cpu_req_ready;
  wire[4:0] ptw_io_mem_req_bits_cmd;
  wire[43:0] ptw_io_mem_req_bits_addr;
  wire ptw_io_mem_req_bits_phys;
  wire[2:0] ptw_io_mem_req_bits_typ;
  wire ptw_io_mem_req_bits_kill;
  wire ptw_io_mem_req_valid;
  wire[4:0] core_io_dmem_req_bits_cmd;
  wire[7:0] core_io_dmem_req_bits_tag;
  wire[63:0] core_io_dmem_req_bits_data;
  wire[43:0] core_io_dmem_req_bits_addr;
  wire core_io_dmem_req_bits_phys;
  wire[2:0] core_io_dmem_req_bits_typ;
  wire core_io_dmem_req_bits_kill;
  wire core_io_dmem_req_valid;
  wire dcArb_io_requestor_1_ordered;
  wire dcArb_io_requestor_1_xcpt_pf_st;
  wire dcArb_io_requestor_1_xcpt_pf_ld;
  wire dcArb_io_requestor_1_xcpt_ma_st;
  wire dcArb_io_requestor_1_xcpt_ma_ld;
  wire[7:0] dcArb_io_requestor_1_replay_next_bits;
  wire dcArb_io_requestor_1_replay_next_valid;
  wire[63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire[43:0] dcArb_io_requestor_1_resp_bits_addr;
  wire[3:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire[7:0] dcArb_io_requestor_1_resp_bits_tag;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data_subword;
  wire[63:0] dcArb_io_requestor_1_resp_bits_data;
  wire dcArb_io_requestor_1_resp_bits_has_data;
  wire[2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire dcArb_io_requestor_1_resp_bits_replay;
  wire dcArb_io_requestor_1_resp_bits_nack;
  wire dcArb_io_requestor_1_resp_valid;
  wire dcArb_io_requestor_1_req_ready;
  wire[29:0] icache_io_cpu_ptw_req_bits;
  wire icache_io_cpu_ptw_req_valid;
  wire[1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire[3:0] icache_io_cpu_btb_resp_bits_bht_index;
  wire[2:0] icache_io_cpu_btb_resp_bits_entry;
  wire[42:0] icache_io_cpu_btb_resp_bits_target;
  wire icache_io_cpu_btb_resp_bits_taken;
  wire icache_io_cpu_btb_resp_valid;
  wire icache_io_cpu_resp_bits_xcpt_if;
  wire icache_io_cpu_resp_bits_xcpt_ma;
  wire[31:0] icache_io_cpu_resp_bits_data;
  wire[43:0] icache_io_cpu_resp_bits_pc;
  wire icache_io_cpu_resp_valid;
  wire core_io_ptw_status_s;
  wire core_io_ptw_status_ps;
  wire core_io_ptw_status_ei;
  wire core_io_ptw_status_pei;
  wire core_io_ptw_status_ef;
  wire core_io_ptw_status_u64;
  wire core_io_ptw_status_s64;
  wire core_io_ptw_status_vm;
  wire core_io_ptw_status_er;
  wire[6:0] core_io_ptw_status_zero;
  wire[7:0] core_io_ptw_status_im;
  wire[7:0] core_io_ptw_status_ip;
  wire core_io_ptw_sret;
  wire core_io_ptw_invalidate;
  wire[31:0] core_io_ptw_ptbr;
  wire dcArb_io_requestor_0_ordered;
  wire dcArb_io_requestor_0_xcpt_pf_st;
  wire dcArb_io_requestor_0_xcpt_pf_ld;
  wire dcArb_io_requestor_0_xcpt_ma_st;
  wire dcArb_io_requestor_0_xcpt_ma_ld;
  wire[7:0] dcArb_io_requestor_0_replay_next_bits;
  wire dcArb_io_requestor_0_replay_next_valid;
  wire[63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire[43:0] dcArb_io_requestor_0_resp_bits_addr;
  wire[3:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire[7:0] dcArb_io_requestor_0_resp_bits_tag;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data_subword;
  wire[63:0] dcArb_io_requestor_0_resp_bits_data;
  wire dcArb_io_requestor_0_resp_bits_has_data;
  wire[2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire dcArb_io_requestor_0_resp_bits_replay;
  wire dcArb_io_requestor_0_resp_bits_nack;
  wire dcArb_io_requestor_0_resp_valid;
  wire dcArb_io_requestor_0_req_ready;
  wire memArb_io_in_0_finish_ready;
  wire[3:0] memArb_io_in_0_grant_bits_payload_g_type;
  wire[2:0] memArb_io_in_0_grant_bits_payload_master_xact_id;
  wire[1:0] memArb_io_in_0_grant_bits_payload_client_xact_id;
  wire[511:0] memArb_io_in_0_grant_bits_payload_data;
  wire[1:0] memArb_io_in_0_grant_bits_header_dst;
  wire[1:0] memArb_io_in_0_grant_bits_header_src;
  wire memArb_io_in_0_grant_valid;
  wire memArb_io_in_0_acquire_ready;
  wire ptw_io_requestor_1_sret;
  wire ptw_io_requestor_1_invalidate;
  wire ptw_io_requestor_1_status_s;
  wire ptw_io_requestor_1_status_ps;
  wire ptw_io_requestor_1_status_ei;
  wire ptw_io_requestor_1_status_pei;
  wire ptw_io_requestor_1_status_ef;
  wire ptw_io_requestor_1_status_u64;
  wire ptw_io_requestor_1_status_s64;
  wire ptw_io_requestor_1_status_vm;
  wire ptw_io_requestor_1_status_er;
  wire[6:0] ptw_io_requestor_1_status_zero;
  wire[7:0] ptw_io_requestor_1_status_im;
  wire[7:0] ptw_io_requestor_1_status_ip;
  wire[5:0] ptw_io_requestor_1_resp_bits_perm;
  wire[18:0] ptw_io_requestor_1_resp_bits_ppn;
  wire ptw_io_requestor_1_resp_bits_error;
  wire ptw_io_requestor_1_resp_valid;
  wire ptw_io_requestor_1_req_ready;
  wire[4:0] dcArb_io_mem_req_bits_cmd;
  wire[7:0] dcArb_io_mem_req_bits_tag;
  wire[63:0] dcArb_io_mem_req_bits_data;
  wire[43:0] dcArb_io_mem_req_bits_addr;
  wire dcArb_io_mem_req_bits_phys;
  wire[2:0] dcArb_io_mem_req_bits_typ;
  wire dcArb_io_mem_req_bits_kill;
  wire dcArb_io_mem_req_valid;
  wire memArb_io_in_1_finish_ready;
  wire[3:0] memArb_io_in_1_grant_bits_payload_g_type;
  wire[2:0] memArb_io_in_1_grant_bits_payload_master_xact_id;
  wire[1:0] memArb_io_in_1_grant_bits_payload_client_xact_id;
  wire[511:0] memArb_io_in_1_grant_bits_payload_data;
  wire[1:0] memArb_io_in_1_grant_bits_header_dst;
  wire[1:0] memArb_io_in_1_grant_bits_header_src;
  wire memArb_io_in_1_grant_valid;
  wire memArb_io_in_1_acquire_ready;
  wire core_io_imem_invalidate;
  wire ptw_io_requestor_0_sret;
  wire ptw_io_requestor_0_invalidate;
  wire ptw_io_requestor_0_status_s;
  wire ptw_io_requestor_0_status_ps;
  wire ptw_io_requestor_0_status_ei;
  wire ptw_io_requestor_0_status_pei;
  wire ptw_io_requestor_0_status_ef;
  wire ptw_io_requestor_0_status_u64;
  wire ptw_io_requestor_0_status_s64;
  wire ptw_io_requestor_0_status_vm;
  wire ptw_io_requestor_0_status_er;
  wire[6:0] ptw_io_requestor_0_status_zero;
  wire[7:0] ptw_io_requestor_0_status_im;
  wire[7:0] ptw_io_requestor_0_status_ip;
  wire[5:0] ptw_io_requestor_0_resp_bits_perm;
  wire[18:0] ptw_io_requestor_0_resp_bits_ppn;
  wire ptw_io_requestor_0_resp_bits_error;
  wire ptw_io_requestor_0_resp_valid;
  wire ptw_io_requestor_0_req_ready;
  wire core_io_imem_btb_update_bits_incorrectTarget;
  wire core_io_imem_btb_update_bits_isReturn;
  wire core_io_imem_btb_update_bits_isCall;
  wire core_io_imem_btb_update_bits_isJump;
  wire core_io_imem_btb_update_bits_taken;
  wire[42:0] core_io_imem_btb_update_bits_returnAddr;
  wire[42:0] core_io_imem_btb_update_bits_target;
  wire[42:0] core_io_imem_btb_update_bits_pc;
  wire[1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire[3:0] core_io_imem_btb_update_bits_prediction_bits_bht_index;
  wire[2:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire[42:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire core_io_imem_btb_update_bits_prediction_bits_taken;
  wire core_io_imem_btb_update_bits_prediction_valid;
  wire core_io_imem_btb_update_valid;
  wire core_io_imem_resp_ready;
  wire[43:0] core_io_imem_req_bits_pc;
  wire core_io_imem_req_valid;
  wire core_io_host_debug_stats_pcr;
  wire core_io_host_ipi_rep_ready;
  wire core_io_host_ipi_req_bits;
  wire core_io_host_ipi_req_valid;
  wire[63:0] core_io_host_pcr_rep_bits;
  wire core_io_host_pcr_rep_valid;
  wire core_io_host_pcr_req_ready;
  wire[2:0] dcache_io_mem_release_bits_payload_r_type;
  wire[511:0] dcache_io_mem_release_bits_payload_data;
  wire[2:0] dcache_io_mem_release_bits_payload_master_xact_id;
  wire[1:0] T0;
  wire[2:0] T1;
  wire[1:0] dcache_io_mem_release_bits_payload_client_xact_id;
  wire[25:0] dcache_io_mem_release_bits_payload_addr;
  wire[1:0] dcache_io_mem_release_bits_header_dst;
  wire[1:0] dcache_io_mem_release_bits_header_src;
  wire dcache_io_mem_release_valid;
  wire dcache_io_mem_probe_ready;
  wire[2:0] memArb_io_out_finish_bits_payload_master_xact_id;
  wire[1:0] memArb_io_out_finish_bits_header_dst;
  wire[1:0] memArb_io_out_finish_bits_header_src;
  wire memArb_io_out_finish_valid;
  wire memArb_io_out_grant_ready;
  wire[3:0] memArb_io_out_acquire_bits_payload_atomic_opcode;
  wire[2:0] memArb_io_out_acquire_bits_payload_subword_addr;
  wire[5:0] memArb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] memArb_io_out_acquire_bits_payload_a_type;
  wire[511:0] memArb_io_out_acquire_bits_payload_data;
  wire[1:0] memArb_io_out_acquire_bits_payload_client_xact_id;
  wire[25:0] memArb_io_out_acquire_bits_payload_addr;
  wire[1:0] memArb_io_out_acquire_bits_header_dst;
  wire[1:0] memArb_io_out_acquire_bits_header_src;
  wire memArb_io_out_acquire_valid;


  assign io_host_debug_stats_pcr = core_io_host_debug_stats_pcr;
  assign io_host_ipi_rep_ready = core_io_host_ipi_rep_ready;
  assign io_host_ipi_req_bits = core_io_host_ipi_req_bits;
  assign io_host_ipi_req_valid = core_io_host_ipi_req_valid;
  assign io_host_pcr_rep_bits = core_io_host_pcr_rep_bits;
  assign io_host_pcr_rep_valid = core_io_host_pcr_rep_valid;
  assign io_host_pcr_req_ready = core_io_host_pcr_req_ready;
  assign io_tilelink_release_bits_payload_r_type = dcache_io_mem_release_bits_payload_r_type;
  assign io_tilelink_release_bits_payload_data = dcache_io_mem_release_bits_payload_data;
  assign io_tilelink_release_bits_payload_master_xact_id = dcache_io_mem_release_bits_payload_master_xact_id;
  assign io_tilelink_release_bits_payload_client_xact_id = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = {dcache_io_mem_release_bits_payload_client_xact_id, 1'h0};
  assign io_tilelink_release_bits_payload_addr = dcache_io_mem_release_bits_payload_addr;
  assign io_tilelink_release_bits_header_dst = dcache_io_mem_release_bits_header_dst;
  assign io_tilelink_release_bits_header_src = dcache_io_mem_release_bits_header_src;
  assign io_tilelink_release_valid = dcache_io_mem_release_valid;
  assign io_tilelink_probe_ready = dcache_io_mem_probe_ready;
  assign io_tilelink_finish_bits_payload_master_xact_id = memArb_io_out_finish_bits_payload_master_xact_id;
  assign io_tilelink_finish_bits_header_dst = memArb_io_out_finish_bits_header_dst;
  assign io_tilelink_finish_bits_header_src = memArb_io_out_finish_bits_header_src;
  assign io_tilelink_finish_valid = memArb_io_out_finish_valid;
  assign io_tilelink_grant_ready = memArb_io_out_grant_ready;
  assign io_tilelink_acquire_bits_payload_atomic_opcode = memArb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_tilelink_acquire_bits_payload_subword_addr = memArb_io_out_acquire_bits_payload_subword_addr;
  assign io_tilelink_acquire_bits_payload_write_mask = memArb_io_out_acquire_bits_payload_write_mask;
  assign io_tilelink_acquire_bits_payload_a_type = memArb_io_out_acquire_bits_payload_a_type;
  assign io_tilelink_acquire_bits_payload_data = memArb_io_out_acquire_bits_payload_data;
  assign io_tilelink_acquire_bits_payload_client_xact_id = memArb_io_out_acquire_bits_payload_client_xact_id;
  assign io_tilelink_acquire_bits_payload_addr = memArb_io_out_acquire_bits_payload_addr;
  assign io_tilelink_acquire_bits_header_dst = memArb_io_out_acquire_bits_header_dst;
  assign io_tilelink_acquire_bits_header_src = memArb_io_out_acquire_bits_header_src;
  assign io_tilelink_acquire_valid = memArb_io_out_acquire_valid;
  Frontend icache(.clk(clk), .reset(reset),
       .io_cpu_req_valid( core_io_imem_req_valid ),
       .io_cpu_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_cpu_resp_ready( core_io_imem_resp_ready ),
       .io_cpu_resp_valid( icache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_cpu_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_cpu_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_cpu_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_cpu_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_cpu_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_cpu_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_cpu_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_cpu_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_cpu_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_cpu_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_cpu_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_cpu_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_cpu_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_cpu_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_cpu_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_cpu_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_cpu_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_cpu_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_cpu_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_cpu_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_cpu_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_cpu_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_cpu_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_0_req_ready ),
       .io_cpu_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_0_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_0_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_0_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_0_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_0_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_0_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_0_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_0_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_0_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_0_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_0_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_0_sret ),
       .io_cpu_invalidate( core_io_imem_invalidate ),
       .io_mem_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_mem_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( icache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_1_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_1_finish_ready ),
       .io_mem_finish_valid( icache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id )
  );
  HellaCache dcache(.clk(clk), .reset(reset),
       .io_cpu_req_ready( dcache_io_cpu_req_ready ),
       .io_cpu_req_valid( dcArb_io_mem_req_valid ),
       .io_cpu_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_cpu_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_cpu_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_cpu_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_cpu_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_cpu_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_cpu_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_cpu_resp_valid( dcache_io_cpu_resp_valid ),
       .io_cpu_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_cpu_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_cpu_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_cpu_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_cpu_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_cpu_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_cpu_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_cpu_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_cpu_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_cpu_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_cpu_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_cpu_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_cpu_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_cpu_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_cpu_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       .io_cpu_ptw_req_ready( ptw_io_requestor_1_req_ready ),
       .io_cpu_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_cpu_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_cpu_ptw_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_cpu_ptw_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_cpu_ptw_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_cpu_ptw_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_cpu_ptw_status_ip( ptw_io_requestor_1_status_ip ),
       .io_cpu_ptw_status_im( ptw_io_requestor_1_status_im ),
       .io_cpu_ptw_status_zero( ptw_io_requestor_1_status_zero ),
       .io_cpu_ptw_status_er( ptw_io_requestor_1_status_er ),
       .io_cpu_ptw_status_vm( ptw_io_requestor_1_status_vm ),
       .io_cpu_ptw_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_cpu_ptw_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_cpu_ptw_status_ef( ptw_io_requestor_1_status_ef ),
       .io_cpu_ptw_status_pei( ptw_io_requestor_1_status_pei ),
       .io_cpu_ptw_status_ei( ptw_io_requestor_1_status_ei ),
       .io_cpu_ptw_status_ps( ptw_io_requestor_1_status_ps ),
       .io_cpu_ptw_status_s( ptw_io_requestor_1_status_s ),
       .io_cpu_ptw_invalidate( ptw_io_requestor_1_invalidate ),
       .io_cpu_ptw_sret( ptw_io_requestor_1_sret ),
       .io_cpu_ordered( dcache_io_cpu_ordered ),
       .io_mem_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_mem_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_mem_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_mem_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_mem_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( dcache_io_mem_grant_ready ),
       .io_mem_grant_valid( memArb_io_in_0_grant_valid ),
       .io_mem_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_mem_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_mem_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_mem_finish_ready( memArb_io_in_0_finish_ready ),
       .io_mem_finish_valid( dcache_io_mem_finish_valid ),
       .io_mem_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_mem_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( dcache_io_mem_probe_ready ),
       .io_mem_probe_valid( io_tilelink_probe_valid ),
       .io_mem_probe_bits_header_src( io_tilelink_probe_bits_header_src ),
       .io_mem_probe_bits_header_dst( io_tilelink_probe_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( io_tilelink_probe_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( io_tilelink_probe_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( io_tilelink_probe_bits_payload_p_type ),
       .io_mem_release_ready( io_tilelink_release_ready ),
       .io_mem_release_valid( dcache_io_mem_release_valid ),
       .io_mem_release_bits_header_src( dcache_io_mem_release_bits_header_src ),
       .io_mem_release_bits_header_dst( dcache_io_mem_release_bits_header_dst ),
       .io_mem_release_bits_payload_addr( dcache_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( dcache_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( dcache_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( dcache_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( dcache_io_mem_release_bits_payload_r_type )
  );
  PTW ptw(.clk(clk), .reset(reset),
       .io_requestor_1_req_ready( ptw_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_requestor_1_req_bits( dcache_io_cpu_ptw_req_bits ),
       .io_requestor_1_resp_valid( ptw_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_error( ptw_io_requestor_1_resp_bits_error ),
       .io_requestor_1_resp_bits_ppn( ptw_io_requestor_1_resp_bits_ppn ),
       .io_requestor_1_resp_bits_perm( ptw_io_requestor_1_resp_bits_perm ),
       .io_requestor_1_status_ip( ptw_io_requestor_1_status_ip ),
       .io_requestor_1_status_im( ptw_io_requestor_1_status_im ),
       .io_requestor_1_status_zero( ptw_io_requestor_1_status_zero ),
       .io_requestor_1_status_er( ptw_io_requestor_1_status_er ),
       .io_requestor_1_status_vm( ptw_io_requestor_1_status_vm ),
       .io_requestor_1_status_s64( ptw_io_requestor_1_status_s64 ),
       .io_requestor_1_status_u64( ptw_io_requestor_1_status_u64 ),
       .io_requestor_1_status_ef( ptw_io_requestor_1_status_ef ),
       .io_requestor_1_status_pei( ptw_io_requestor_1_status_pei ),
       .io_requestor_1_status_ei( ptw_io_requestor_1_status_ei ),
       .io_requestor_1_status_ps( ptw_io_requestor_1_status_ps ),
       .io_requestor_1_status_s( ptw_io_requestor_1_status_s ),
       .io_requestor_1_invalidate( ptw_io_requestor_1_invalidate ),
       .io_requestor_1_sret( ptw_io_requestor_1_sret ),
       .io_requestor_0_req_ready( ptw_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_requestor_0_req_bits( icache_io_cpu_ptw_req_bits ),
       .io_requestor_0_resp_valid( ptw_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_error( ptw_io_requestor_0_resp_bits_error ),
       .io_requestor_0_resp_bits_ppn( ptw_io_requestor_0_resp_bits_ppn ),
       .io_requestor_0_resp_bits_perm( ptw_io_requestor_0_resp_bits_perm ),
       .io_requestor_0_status_ip( ptw_io_requestor_0_status_ip ),
       .io_requestor_0_status_im( ptw_io_requestor_0_status_im ),
       .io_requestor_0_status_zero( ptw_io_requestor_0_status_zero ),
       .io_requestor_0_status_er( ptw_io_requestor_0_status_er ),
       .io_requestor_0_status_vm( ptw_io_requestor_0_status_vm ),
       .io_requestor_0_status_s64( ptw_io_requestor_0_status_s64 ),
       .io_requestor_0_status_u64( ptw_io_requestor_0_status_u64 ),
       .io_requestor_0_status_ef( ptw_io_requestor_0_status_ef ),
       .io_requestor_0_status_pei( ptw_io_requestor_0_status_pei ),
       .io_requestor_0_status_ei( ptw_io_requestor_0_status_ei ),
       .io_requestor_0_status_ps( ptw_io_requestor_0_status_ps ),
       .io_requestor_0_status_s( ptw_io_requestor_0_status_s ),
       .io_requestor_0_invalidate( ptw_io_requestor_0_invalidate ),
       .io_requestor_0_sret( ptw_io_requestor_0_sret ),
       .io_mem_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_mem_req_valid( ptw_io_mem_req_valid ),
       .io_mem_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_mem_req_bits_data(  )
       //.io_mem_req_bits_tag(  )
       .io_mem_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_mem_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_mem_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       //.io_mem_ptw_req_valid(  )
       //.io_mem_ptw_req_bits(  )
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcArb_io_requestor_0_ordered ),
       .io_dpath_ptbr( core_io_ptw_ptbr ),
       .io_dpath_invalidate( core_io_ptw_invalidate ),
       .io_dpath_sret( core_io_ptw_sret ),
       .io_dpath_status_ip( core_io_ptw_status_ip ),
       .io_dpath_status_im( core_io_ptw_status_im ),
       .io_dpath_status_zero( core_io_ptw_status_zero ),
       .io_dpath_status_er( core_io_ptw_status_er ),
       .io_dpath_status_vm( core_io_ptw_status_vm ),
       .io_dpath_status_s64( core_io_ptw_status_s64 ),
       .io_dpath_status_u64( core_io_ptw_status_u64 ),
       .io_dpath_status_ef( core_io_ptw_status_ef ),
       .io_dpath_status_pei( core_io_ptw_status_pei ),
       .io_dpath_status_ei( core_io_ptw_status_ei ),
       .io_dpath_status_ps( core_io_ptw_status_ps ),
       .io_dpath_status_s( core_io_ptw_status_s )
  );
  Core core(.clk(clk), .reset(reset),
       .io_host_reset( io_host_reset ),
       .io_host_id( io_host_id ),
       .io_host_pcr_req_ready( core_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( io_host_pcr_req_valid ),
       .io_host_pcr_req_bits_rw( io_host_pcr_req_bits_rw ),
       .io_host_pcr_req_bits_addr( io_host_pcr_req_bits_addr ),
       .io_host_pcr_req_bits_data( io_host_pcr_req_bits_data ),
       .io_host_pcr_rep_ready( io_host_pcr_rep_ready ),
       .io_host_pcr_rep_valid( core_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( core_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( io_host_ipi_req_ready ),
       .io_host_ipi_req_valid( core_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( core_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( core_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( io_host_ipi_rep_valid ),
       .io_host_ipi_rep_bits( io_host_ipi_rep_bits ),
       .io_host_debug_stats_pcr( core_io_host_debug_stats_pcr ),
       .io_imem_req_valid( core_io_imem_req_valid ),
       .io_imem_req_bits_pc( core_io_imem_req_bits_pc ),
       .io_imem_resp_ready( core_io_imem_resp_ready ),
       .io_imem_resp_valid( icache_io_cpu_resp_valid ),
       .io_imem_resp_bits_pc( icache_io_cpu_resp_bits_pc ),
       .io_imem_resp_bits_data( icache_io_cpu_resp_bits_data ),
       .io_imem_resp_bits_xcpt_ma( icache_io_cpu_resp_bits_xcpt_ma ),
       .io_imem_resp_bits_xcpt_if( icache_io_cpu_resp_bits_xcpt_if ),
       .io_imem_btb_resp_valid( icache_io_cpu_btb_resp_valid ),
       .io_imem_btb_resp_bits_taken( icache_io_cpu_btb_resp_bits_taken ),
       .io_imem_btb_resp_bits_target( icache_io_cpu_btb_resp_bits_target ),
       .io_imem_btb_resp_bits_entry( icache_io_cpu_btb_resp_bits_entry ),
       .io_imem_btb_resp_bits_bht_index( icache_io_cpu_btb_resp_bits_bht_index ),
       .io_imem_btb_resp_bits_bht_value( icache_io_cpu_btb_resp_bits_bht_value ),
       .io_imem_btb_update_valid( core_io_imem_btb_update_valid ),
       .io_imem_btb_update_bits_prediction_valid( core_io_imem_btb_update_bits_prediction_valid ),
       .io_imem_btb_update_bits_prediction_bits_taken( core_io_imem_btb_update_bits_prediction_bits_taken ),
       .io_imem_btb_update_bits_prediction_bits_target( core_io_imem_btb_update_bits_prediction_bits_target ),
       .io_imem_btb_update_bits_prediction_bits_entry( core_io_imem_btb_update_bits_prediction_bits_entry ),
       .io_imem_btb_update_bits_prediction_bits_bht_index( core_io_imem_btb_update_bits_prediction_bits_bht_index ),
       .io_imem_btb_update_bits_prediction_bits_bht_value( core_io_imem_btb_update_bits_prediction_bits_bht_value ),
       .io_imem_btb_update_bits_pc( core_io_imem_btb_update_bits_pc ),
       .io_imem_btb_update_bits_target( core_io_imem_btb_update_bits_target ),
       .io_imem_btb_update_bits_returnAddr( core_io_imem_btb_update_bits_returnAddr ),
       .io_imem_btb_update_bits_taken( core_io_imem_btb_update_bits_taken ),
       .io_imem_btb_update_bits_isJump( core_io_imem_btb_update_bits_isJump ),
       .io_imem_btb_update_bits_isCall( core_io_imem_btb_update_bits_isCall ),
       .io_imem_btb_update_bits_isReturn( core_io_imem_btb_update_bits_isReturn ),
       .io_imem_btb_update_bits_incorrectTarget( core_io_imem_btb_update_bits_incorrectTarget ),
       //.io_imem_ptw_req_ready(  )
       .io_imem_ptw_req_valid( icache_io_cpu_ptw_req_valid ),
       .io_imem_ptw_req_bits( icache_io_cpu_ptw_req_bits ),
       //.io_imem_ptw_resp_valid(  )
       //.io_imem_ptw_resp_bits_error(  )
       //.io_imem_ptw_resp_bits_ppn(  )
       //.io_imem_ptw_resp_bits_perm(  )
       //.io_imem_ptw_status_ip(  )
       //.io_imem_ptw_status_im(  )
       //.io_imem_ptw_status_zero(  )
       //.io_imem_ptw_status_er(  )
       //.io_imem_ptw_status_vm(  )
       //.io_imem_ptw_status_s64(  )
       //.io_imem_ptw_status_u64(  )
       //.io_imem_ptw_status_ef(  )
       //.io_imem_ptw_status_pei(  )
       //.io_imem_ptw_status_ei(  )
       //.io_imem_ptw_status_ps(  )
       //.io_imem_ptw_status_s(  )
       //.io_imem_ptw_invalidate(  )
       //.io_imem_ptw_sret(  )
       .io_imem_invalidate( core_io_imem_invalidate ),
       .io_dmem_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_dmem_req_valid( core_io_dmem_req_valid ),
       .io_dmem_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_dmem_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_dmem_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_dmem_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_dmem_req_bits_data( core_io_dmem_req_bits_data ),
       .io_dmem_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_dmem_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_dmem_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_dmem_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_dmem_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_dmem_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_dmem_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_dmem_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_dmem_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_dmem_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_dmem_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_dmem_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_dmem_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_dmem_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_dmem_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_dmem_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_dmem_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_dmem_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_dmem_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_dmem_ptw_req_ready(  )
       //.io_dmem_ptw_req_valid(  )
       //.io_dmem_ptw_req_bits(  )
       //.io_dmem_ptw_resp_valid(  )
       //.io_dmem_ptw_resp_bits_error(  )
       //.io_dmem_ptw_resp_bits_ppn(  )
       //.io_dmem_ptw_resp_bits_perm(  )
       //.io_dmem_ptw_status_ip(  )
       //.io_dmem_ptw_status_im(  )
       //.io_dmem_ptw_status_zero(  )
       //.io_dmem_ptw_status_er(  )
       //.io_dmem_ptw_status_vm(  )
       //.io_dmem_ptw_status_s64(  )
       //.io_dmem_ptw_status_u64(  )
       //.io_dmem_ptw_status_ef(  )
       //.io_dmem_ptw_status_pei(  )
       //.io_dmem_ptw_status_ei(  )
       //.io_dmem_ptw_status_ps(  )
       //.io_dmem_ptw_status_s(  )
       //.io_dmem_ptw_invalidate(  )
       //.io_dmem_ptw_sret(  )
       .io_dmem_ordered( dcArb_io_requestor_1_ordered ),
       .io_ptw_ptbr( core_io_ptw_ptbr ),
       .io_ptw_invalidate( core_io_ptw_invalidate ),
       .io_ptw_sret( core_io_ptw_sret ),
       .io_ptw_status_ip( core_io_ptw_status_ip ),
       .io_ptw_status_im( core_io_ptw_status_im ),
       .io_ptw_status_zero( core_io_ptw_status_zero ),
       .io_ptw_status_er( core_io_ptw_status_er ),
       .io_ptw_status_vm( core_io_ptw_status_vm ),
       .io_ptw_status_s64( core_io_ptw_status_s64 ),
       .io_ptw_status_u64( core_io_ptw_status_u64 ),
       .io_ptw_status_ef( core_io_ptw_status_ef ),
       .io_ptw_status_pei( core_io_ptw_status_pei ),
       .io_ptw_status_ei( core_io_ptw_status_ei ),
       .io_ptw_status_ps( core_io_ptw_status_ps ),
       .io_ptw_status_s( core_io_ptw_status_s )
       //.io_rocc_cmd_ready(  )
       //.io_rocc_cmd_valid(  )
       //.io_rocc_cmd_bits_inst_funct(  )
       //.io_rocc_cmd_bits_inst_rs2(  )
       //.io_rocc_cmd_bits_inst_rs1(  )
       //.io_rocc_cmd_bits_inst_xd(  )
       //.io_rocc_cmd_bits_inst_xs1(  )
       //.io_rocc_cmd_bits_inst_xs2(  )
       //.io_rocc_cmd_bits_inst_rd(  )
       //.io_rocc_cmd_bits_inst_opcode(  )
       //.io_rocc_cmd_bits_rs1(  )
       //.io_rocc_cmd_bits_rs2(  )
       //.io_rocc_resp_ready(  )
       //.io_rocc_resp_valid(  )
       //.io_rocc_resp_bits_rd(  )
       //.io_rocc_resp_bits_data(  )
       //.io_rocc_mem_req_ready(  )
       //.io_rocc_mem_req_valid(  )
       //.io_rocc_mem_req_bits_kill(  )
       //.io_rocc_mem_req_bits_typ(  )
       //.io_rocc_mem_req_bits_phys(  )
       //.io_rocc_mem_req_bits_addr(  )
       //.io_rocc_mem_req_bits_data(  )
       //.io_rocc_mem_req_bits_tag(  )
       //.io_rocc_mem_req_bits_cmd(  )
       //.io_rocc_mem_resp_valid(  )
       //.io_rocc_mem_resp_bits_nack(  )
       //.io_rocc_mem_resp_bits_replay(  )
       //.io_rocc_mem_resp_bits_typ(  )
       //.io_rocc_mem_resp_bits_has_data(  )
       //.io_rocc_mem_resp_bits_data(  )
       //.io_rocc_mem_resp_bits_data_subword(  )
       //.io_rocc_mem_resp_bits_tag(  )
       //.io_rocc_mem_resp_bits_cmd(  )
       //.io_rocc_mem_resp_bits_addr(  )
       //.io_rocc_mem_resp_bits_store_data(  )
       //.io_rocc_mem_replay_next_valid(  )
       //.io_rocc_mem_replay_next_bits(  )
       //.io_rocc_mem_xcpt_ma_ld(  )
       //.io_rocc_mem_xcpt_ma_st(  )
       //.io_rocc_mem_xcpt_pf_ld(  )
       //.io_rocc_mem_xcpt_pf_st(  )
       //.io_rocc_mem_ptw_req_ready(  )
       //.io_rocc_mem_ptw_req_valid(  )
       //.io_rocc_mem_ptw_req_bits(  )
       //.io_rocc_mem_ptw_resp_valid(  )
       //.io_rocc_mem_ptw_resp_bits_error(  )
       //.io_rocc_mem_ptw_resp_bits_ppn(  )
       //.io_rocc_mem_ptw_resp_bits_perm(  )
       //.io_rocc_mem_ptw_status_ip(  )
       //.io_rocc_mem_ptw_status_im(  )
       //.io_rocc_mem_ptw_status_zero(  )
       //.io_rocc_mem_ptw_status_er(  )
       //.io_rocc_mem_ptw_status_vm(  )
       //.io_rocc_mem_ptw_status_s64(  )
       //.io_rocc_mem_ptw_status_u64(  )
       //.io_rocc_mem_ptw_status_ef(  )
       //.io_rocc_mem_ptw_status_pei(  )
       //.io_rocc_mem_ptw_status_ei(  )
       //.io_rocc_mem_ptw_status_ps(  )
       //.io_rocc_mem_ptw_status_s(  )
       //.io_rocc_mem_ptw_invalidate(  )
       //.io_rocc_mem_ptw_sret(  )
       //.io_rocc_mem_ordered(  )
       //.io_rocc_busy(  )
       //.io_rocc_s(  )
       //.io_rocc_interrupt(  )
       //.io_rocc_imem_acquire_ready(  )
       //.io_rocc_imem_acquire_valid(  )
       //.io_rocc_imem_acquire_bits_header_src(  )
       //.io_rocc_imem_acquire_bits_header_dst(  )
       //.io_rocc_imem_acquire_bits_payload_addr(  )
       //.io_rocc_imem_acquire_bits_payload_client_xact_id(  )
       //.io_rocc_imem_acquire_bits_payload_data(  )
       //.io_rocc_imem_acquire_bits_payload_a_type(  )
       //.io_rocc_imem_acquire_bits_payload_write_mask(  )
       //.io_rocc_imem_acquire_bits_payload_subword_addr(  )
       //.io_rocc_imem_acquire_bits_payload_atomic_opcode(  )
       //.io_rocc_imem_grant_ready(  )
       //.io_rocc_imem_grant_valid(  )
       //.io_rocc_imem_grant_bits_header_src(  )
       //.io_rocc_imem_grant_bits_header_dst(  )
       //.io_rocc_imem_grant_bits_payload_data(  )
       //.io_rocc_imem_grant_bits_payload_client_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_master_xact_id(  )
       //.io_rocc_imem_grant_bits_payload_g_type(  )
       //.io_rocc_imem_finish_ready(  )
       //.io_rocc_imem_finish_valid(  )
       //.io_rocc_imem_finish_bits_header_src(  )
       //.io_rocc_imem_finish_bits_header_dst(  )
       //.io_rocc_imem_finish_bits_payload_master_xact_id(  )
       //.io_rocc_iptw_req_ready(  )
       //.io_rocc_iptw_req_valid(  )
       //.io_rocc_iptw_req_bits(  )
       //.io_rocc_iptw_resp_valid(  )
       //.io_rocc_iptw_resp_bits_error(  )
       //.io_rocc_iptw_resp_bits_ppn(  )
       //.io_rocc_iptw_resp_bits_perm(  )
       //.io_rocc_iptw_status_ip(  )
       //.io_rocc_iptw_status_im(  )
       //.io_rocc_iptw_status_zero(  )
       //.io_rocc_iptw_status_er(  )
       //.io_rocc_iptw_status_vm(  )
       //.io_rocc_iptw_status_s64(  )
       //.io_rocc_iptw_status_u64(  )
       //.io_rocc_iptw_status_ef(  )
       //.io_rocc_iptw_status_pei(  )
       //.io_rocc_iptw_status_ei(  )
       //.io_rocc_iptw_status_ps(  )
       //.io_rocc_iptw_status_s(  )
       //.io_rocc_iptw_invalidate(  )
       //.io_rocc_iptw_sret(  )
       //.io_rocc_dptw_req_ready(  )
       //.io_rocc_dptw_req_valid(  )
       //.io_rocc_dptw_req_bits(  )
       //.io_rocc_dptw_resp_valid(  )
       //.io_rocc_dptw_resp_bits_error(  )
       //.io_rocc_dptw_resp_bits_ppn(  )
       //.io_rocc_dptw_resp_bits_perm(  )
       //.io_rocc_dptw_status_ip(  )
       //.io_rocc_dptw_status_im(  )
       //.io_rocc_dptw_status_zero(  )
       //.io_rocc_dptw_status_er(  )
       //.io_rocc_dptw_status_vm(  )
       //.io_rocc_dptw_status_s64(  )
       //.io_rocc_dptw_status_u64(  )
       //.io_rocc_dptw_status_ef(  )
       //.io_rocc_dptw_status_pei(  )
       //.io_rocc_dptw_status_ei(  )
       //.io_rocc_dptw_status_ps(  )
       //.io_rocc_dptw_status_s(  )
       //.io_rocc_dptw_invalidate(  )
       //.io_rocc_dptw_sret(  )
       //.io_rocc_pptw_req_ready(  )
       //.io_rocc_pptw_req_valid(  )
       //.io_rocc_pptw_req_bits(  )
       //.io_rocc_pptw_resp_valid(  )
       //.io_rocc_pptw_resp_bits_error(  )
       //.io_rocc_pptw_resp_bits_ppn(  )
       //.io_rocc_pptw_resp_bits_perm(  )
       //.io_rocc_pptw_status_ip(  )
       //.io_rocc_pptw_status_im(  )
       //.io_rocc_pptw_status_zero(  )
       //.io_rocc_pptw_status_er(  )
       //.io_rocc_pptw_status_vm(  )
       //.io_rocc_pptw_status_s64(  )
       //.io_rocc_pptw_status_u64(  )
       //.io_rocc_pptw_status_ef(  )
       //.io_rocc_pptw_status_pei(  )
       //.io_rocc_pptw_status_ei(  )
       //.io_rocc_pptw_status_ps(  )
       //.io_rocc_pptw_status_s(  )
       //.io_rocc_pptw_invalidate(  )
       //.io_rocc_pptw_sret(  )
       //.io_rocc_exception(  )
  );
  `ifndef SYNTHESIS
    assign core.io_dmem_ptw_req_valid = {1{$random}};
    assign core.io_dmem_ptw_req_bits = {1{$random}};
    assign core.io_rocc_cmd_ready = {1{$random}};
    assign core.io_rocc_resp_valid = {1{$random}};
    assign core.io_rocc_resp_bits_rd = {1{$random}};
    assign core.io_rocc_resp_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_valid = {1{$random}};
    assign core.io_rocc_mem_req_bits_kill = {1{$random}};
    assign core.io_rocc_mem_req_bits_typ = {1{$random}};
    assign core.io_rocc_mem_req_bits_phys = {1{$random}};
    assign core.io_rocc_mem_req_bits_addr = {2{$random}};
    assign core.io_rocc_mem_req_bits_data = {2{$random}};
    assign core.io_rocc_mem_req_bits_tag = {1{$random}};
    assign core.io_rocc_mem_req_bits_cmd = {1{$random}};
    assign core.io_rocc_mem_ptw_req_ready = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_valid = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_error = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_ppn = {1{$random}};
    assign core.io_rocc_mem_ptw_resp_bits_perm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ip = {1{$random}};
    assign core.io_rocc_mem_ptw_status_im = {1{$random}};
    assign core.io_rocc_mem_ptw_status_zero = {1{$random}};
    assign core.io_rocc_mem_ptw_status_er = {1{$random}};
    assign core.io_rocc_mem_ptw_status_vm = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_u64 = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ef = {1{$random}};
    assign core.io_rocc_mem_ptw_status_pei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ei = {1{$random}};
    assign core.io_rocc_mem_ptw_status_ps = {1{$random}};
    assign core.io_rocc_mem_ptw_status_s = {1{$random}};
    assign core.io_rocc_mem_ptw_invalidate = {1{$random}};
    assign core.io_rocc_mem_ptw_sret = {1{$random}};
    assign core.io_rocc_busy = {1{$random}};
    assign core.io_rocc_interrupt = {1{$random}};
    assign core.io_rocc_imem_acquire_valid = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_client_xact_id = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_data = {16{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_a_type = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_write_mask = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_subword_addr = {1{$random}};
    assign core.io_rocc_imem_acquire_bits_payload_atomic_opcode = {1{$random}};
    assign core.io_rocc_imem_grant_ready = {1{$random}};
    assign core.io_rocc_imem_finish_valid = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_src = {1{$random}};
    assign core.io_rocc_imem_finish_bits_header_dst = {1{$random}};
    assign core.io_rocc_imem_finish_bits_payload_master_xact_id = {1{$random}};
    assign core.io_rocc_iptw_req_valid = {1{$random}};
    assign core.io_rocc_iptw_req_bits = {1{$random}};
    assign core.io_rocc_dptw_req_valid = {1{$random}};
    assign core.io_rocc_dptw_req_bits = {1{$random}};
    assign core.io_rocc_pptw_req_valid = {1{$random}};
    assign core.io_rocc_pptw_req_bits = {1{$random}};
  `endif
  HellaCacheArbiter dcArb(.clk(clk),
       .io_requestor_1_req_ready( dcArb_io_requestor_1_req_ready ),
       .io_requestor_1_req_valid( core_io_dmem_req_valid ),
       .io_requestor_1_req_bits_kill( core_io_dmem_req_bits_kill ),
       .io_requestor_1_req_bits_typ( core_io_dmem_req_bits_typ ),
       .io_requestor_1_req_bits_phys( core_io_dmem_req_bits_phys ),
       .io_requestor_1_req_bits_addr( core_io_dmem_req_bits_addr ),
       .io_requestor_1_req_bits_data( core_io_dmem_req_bits_data ),
       .io_requestor_1_req_bits_tag( core_io_dmem_req_bits_tag ),
       .io_requestor_1_req_bits_cmd( core_io_dmem_req_bits_cmd ),
       .io_requestor_1_resp_valid( dcArb_io_requestor_1_resp_valid ),
       .io_requestor_1_resp_bits_nack( dcArb_io_requestor_1_resp_bits_nack ),
       .io_requestor_1_resp_bits_replay( dcArb_io_requestor_1_resp_bits_replay ),
       .io_requestor_1_resp_bits_typ( dcArb_io_requestor_1_resp_bits_typ ),
       .io_requestor_1_resp_bits_has_data( dcArb_io_requestor_1_resp_bits_has_data ),
       .io_requestor_1_resp_bits_data( dcArb_io_requestor_1_resp_bits_data ),
       .io_requestor_1_resp_bits_data_subword( dcArb_io_requestor_1_resp_bits_data_subword ),
       .io_requestor_1_resp_bits_tag( dcArb_io_requestor_1_resp_bits_tag ),
       .io_requestor_1_resp_bits_cmd( dcArb_io_requestor_1_resp_bits_cmd ),
       .io_requestor_1_resp_bits_addr( dcArb_io_requestor_1_resp_bits_addr ),
       .io_requestor_1_resp_bits_store_data( dcArb_io_requestor_1_resp_bits_store_data ),
       .io_requestor_1_replay_next_valid( dcArb_io_requestor_1_replay_next_valid ),
       .io_requestor_1_replay_next_bits( dcArb_io_requestor_1_replay_next_bits ),
       .io_requestor_1_xcpt_ma_ld( dcArb_io_requestor_1_xcpt_ma_ld ),
       .io_requestor_1_xcpt_ma_st( dcArb_io_requestor_1_xcpt_ma_st ),
       .io_requestor_1_xcpt_pf_ld( dcArb_io_requestor_1_xcpt_pf_ld ),
       .io_requestor_1_xcpt_pf_st( dcArb_io_requestor_1_xcpt_pf_st ),
       //.io_requestor_1_ptw_req_ready(  )
       //.io_requestor_1_ptw_req_valid(  )
       //.io_requestor_1_ptw_req_bits(  )
       //.io_requestor_1_ptw_resp_valid(  )
       //.io_requestor_1_ptw_resp_bits_error(  )
       //.io_requestor_1_ptw_resp_bits_ppn(  )
       //.io_requestor_1_ptw_resp_bits_perm(  )
       //.io_requestor_1_ptw_status_ip(  )
       //.io_requestor_1_ptw_status_im(  )
       //.io_requestor_1_ptw_status_zero(  )
       //.io_requestor_1_ptw_status_er(  )
       //.io_requestor_1_ptw_status_vm(  )
       //.io_requestor_1_ptw_status_s64(  )
       //.io_requestor_1_ptw_status_u64(  )
       //.io_requestor_1_ptw_status_ef(  )
       //.io_requestor_1_ptw_status_pei(  )
       //.io_requestor_1_ptw_status_ei(  )
       //.io_requestor_1_ptw_status_ps(  )
       //.io_requestor_1_ptw_status_s(  )
       //.io_requestor_1_ptw_invalidate(  )
       //.io_requestor_1_ptw_sret(  )
       .io_requestor_1_ordered( dcArb_io_requestor_1_ordered ),
       .io_requestor_0_req_ready( dcArb_io_requestor_0_req_ready ),
       .io_requestor_0_req_valid( ptw_io_mem_req_valid ),
       .io_requestor_0_req_bits_kill( ptw_io_mem_req_bits_kill ),
       .io_requestor_0_req_bits_typ( ptw_io_mem_req_bits_typ ),
       .io_requestor_0_req_bits_phys( ptw_io_mem_req_bits_phys ),
       .io_requestor_0_req_bits_addr( ptw_io_mem_req_bits_addr ),
       //.io_requestor_0_req_bits_data(  )
       //.io_requestor_0_req_bits_tag(  )
       .io_requestor_0_req_bits_cmd( ptw_io_mem_req_bits_cmd ),
       .io_requestor_0_resp_valid( dcArb_io_requestor_0_resp_valid ),
       .io_requestor_0_resp_bits_nack( dcArb_io_requestor_0_resp_bits_nack ),
       .io_requestor_0_resp_bits_replay( dcArb_io_requestor_0_resp_bits_replay ),
       .io_requestor_0_resp_bits_typ( dcArb_io_requestor_0_resp_bits_typ ),
       .io_requestor_0_resp_bits_has_data( dcArb_io_requestor_0_resp_bits_has_data ),
       .io_requestor_0_resp_bits_data( dcArb_io_requestor_0_resp_bits_data ),
       .io_requestor_0_resp_bits_data_subword( dcArb_io_requestor_0_resp_bits_data_subword ),
       .io_requestor_0_resp_bits_tag( dcArb_io_requestor_0_resp_bits_tag ),
       .io_requestor_0_resp_bits_cmd( dcArb_io_requestor_0_resp_bits_cmd ),
       .io_requestor_0_resp_bits_addr( dcArb_io_requestor_0_resp_bits_addr ),
       .io_requestor_0_resp_bits_store_data( dcArb_io_requestor_0_resp_bits_store_data ),
       .io_requestor_0_replay_next_valid( dcArb_io_requestor_0_replay_next_valid ),
       .io_requestor_0_replay_next_bits( dcArb_io_requestor_0_replay_next_bits ),
       .io_requestor_0_xcpt_ma_ld( dcArb_io_requestor_0_xcpt_ma_ld ),
       .io_requestor_0_xcpt_ma_st( dcArb_io_requestor_0_xcpt_ma_st ),
       .io_requestor_0_xcpt_pf_ld( dcArb_io_requestor_0_xcpt_pf_ld ),
       .io_requestor_0_xcpt_pf_st( dcArb_io_requestor_0_xcpt_pf_st ),
       //.io_requestor_0_ptw_req_ready(  )
       //.io_requestor_0_ptw_req_valid(  )
       //.io_requestor_0_ptw_req_bits(  )
       //.io_requestor_0_ptw_resp_valid(  )
       //.io_requestor_0_ptw_resp_bits_error(  )
       //.io_requestor_0_ptw_resp_bits_ppn(  )
       //.io_requestor_0_ptw_resp_bits_perm(  )
       //.io_requestor_0_ptw_status_ip(  )
       //.io_requestor_0_ptw_status_im(  )
       //.io_requestor_0_ptw_status_zero(  )
       //.io_requestor_0_ptw_status_er(  )
       //.io_requestor_0_ptw_status_vm(  )
       //.io_requestor_0_ptw_status_s64(  )
       //.io_requestor_0_ptw_status_u64(  )
       //.io_requestor_0_ptw_status_ef(  )
       //.io_requestor_0_ptw_status_pei(  )
       //.io_requestor_0_ptw_status_ei(  )
       //.io_requestor_0_ptw_status_ps(  )
       //.io_requestor_0_ptw_status_s(  )
       //.io_requestor_0_ptw_invalidate(  )
       //.io_requestor_0_ptw_sret(  )
       .io_requestor_0_ordered( dcArb_io_requestor_0_ordered ),
       .io_mem_req_ready( dcache_io_cpu_req_ready ),
       .io_mem_req_valid( dcArb_io_mem_req_valid ),
       .io_mem_req_bits_kill( dcArb_io_mem_req_bits_kill ),
       .io_mem_req_bits_typ( dcArb_io_mem_req_bits_typ ),
       .io_mem_req_bits_phys( dcArb_io_mem_req_bits_phys ),
       .io_mem_req_bits_addr( dcArb_io_mem_req_bits_addr ),
       .io_mem_req_bits_data( dcArb_io_mem_req_bits_data ),
       .io_mem_req_bits_tag( dcArb_io_mem_req_bits_tag ),
       .io_mem_req_bits_cmd( dcArb_io_mem_req_bits_cmd ),
       .io_mem_resp_valid( dcache_io_cpu_resp_valid ),
       .io_mem_resp_bits_nack( dcache_io_cpu_resp_bits_nack ),
       .io_mem_resp_bits_replay( dcache_io_cpu_resp_bits_replay ),
       .io_mem_resp_bits_typ( dcache_io_cpu_resp_bits_typ ),
       .io_mem_resp_bits_has_data( dcache_io_cpu_resp_bits_has_data ),
       .io_mem_resp_bits_data( dcache_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_data_subword( dcache_io_cpu_resp_bits_data_subword ),
       .io_mem_resp_bits_tag( dcache_io_cpu_resp_bits_tag ),
       .io_mem_resp_bits_cmd( dcache_io_cpu_resp_bits_cmd ),
       .io_mem_resp_bits_addr( dcache_io_cpu_resp_bits_addr ),
       .io_mem_resp_bits_store_data( dcache_io_cpu_resp_bits_store_data ),
       .io_mem_replay_next_valid( dcache_io_cpu_replay_next_valid ),
       .io_mem_replay_next_bits( dcache_io_cpu_replay_next_bits ),
       .io_mem_xcpt_ma_ld( dcache_io_cpu_xcpt_ma_ld ),
       .io_mem_xcpt_ma_st( dcache_io_cpu_xcpt_ma_st ),
       .io_mem_xcpt_pf_ld( dcache_io_cpu_xcpt_pf_ld ),
       .io_mem_xcpt_pf_st( dcache_io_cpu_xcpt_pf_st ),
       //.io_mem_ptw_req_ready(  )
       .io_mem_ptw_req_valid( dcache_io_cpu_ptw_req_valid ),
       .io_mem_ptw_req_bits( dcache_io_cpu_ptw_req_bits ),
       //.io_mem_ptw_resp_valid(  )
       //.io_mem_ptw_resp_bits_error(  )
       //.io_mem_ptw_resp_bits_ppn(  )
       //.io_mem_ptw_resp_bits_perm(  )
       //.io_mem_ptw_status_ip(  )
       //.io_mem_ptw_status_im(  )
       //.io_mem_ptw_status_zero(  )
       //.io_mem_ptw_status_er(  )
       //.io_mem_ptw_status_vm(  )
       //.io_mem_ptw_status_s64(  )
       //.io_mem_ptw_status_u64(  )
       //.io_mem_ptw_status_ef(  )
       //.io_mem_ptw_status_pei(  )
       //.io_mem_ptw_status_ei(  )
       //.io_mem_ptw_status_ps(  )
       //.io_mem_ptw_status_s(  )
       //.io_mem_ptw_invalidate(  )
       //.io_mem_ptw_sret(  )
       .io_mem_ordered( dcache_io_cpu_ordered )
  );
  `ifndef SYNTHESIS
    assign dcArb.io_requestor_0_req_bits_data = {2{$random}};
    assign dcArb.io_requestor_0_req_bits_tag = {1{$random}};
  `endif
  UncachedTileLinkIOArbiterThatAppendsArbiterId memArb(.clk(clk), .reset(reset),
       .io_in_1_acquire_ready( memArb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( icache_io_mem_acquire_valid ),
       //.io_in_1_acquire_bits_header_src(  )
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( icache_io_mem_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( icache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( icache_io_mem_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( icache_io_mem_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( icache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( icache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( icache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( icache_io_mem_grant_ready ),
       .io_in_1_grant_valid( memArb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( memArb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( memArb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( memArb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( memArb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( memArb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( memArb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( memArb_io_in_1_finish_ready ),
       .io_in_1_finish_valid( icache_io_mem_finish_valid ),
       .io_in_1_finish_bits_header_src( icache_io_mem_finish_bits_header_src ),
       .io_in_1_finish_bits_header_dst( icache_io_mem_finish_bits_header_dst ),
       .io_in_1_finish_bits_payload_master_xact_id( icache_io_mem_finish_bits_payload_master_xact_id ),
       .io_in_0_acquire_ready( memArb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( dcache_io_mem_acquire_valid ),
       .io_in_0_acquire_bits_header_src( dcache_io_mem_acquire_bits_header_src ),
       .io_in_0_acquire_bits_header_dst( dcache_io_mem_acquire_bits_header_dst ),
       .io_in_0_acquire_bits_payload_addr( dcache_io_mem_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( dcache_io_mem_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( dcache_io_mem_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( dcache_io_mem_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( dcache_io_mem_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( dcache_io_mem_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( dcache_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( dcache_io_mem_grant_ready ),
       .io_in_0_grant_valid( memArb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( memArb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( memArb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( memArb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( memArb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( memArb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( memArb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( memArb_io_in_0_finish_ready ),
       .io_in_0_finish_valid( dcache_io_mem_finish_valid ),
       .io_in_0_finish_bits_header_src( dcache_io_mem_finish_bits_header_src ),
       .io_in_0_finish_bits_header_dst( dcache_io_mem_finish_bits_header_dst ),
       .io_in_0_finish_bits_payload_master_xact_id( dcache_io_mem_finish_bits_payload_master_xact_id ),
       .io_out_acquire_ready( io_tilelink_acquire_ready ),
       .io_out_acquire_valid( memArb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( memArb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( memArb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( memArb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( memArb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( memArb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( memArb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( memArb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( memArb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( memArb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( memArb_io_out_grant_ready ),
       .io_out_grant_valid( io_tilelink_grant_valid ),
       .io_out_grant_bits_header_src( io_tilelink_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_tilelink_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_tilelink_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_tilelink_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_tilelink_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_tilelink_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_tilelink_finish_ready ),
       .io_out_finish_valid( memArb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( memArb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( memArb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( memArb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign memArb.io_in_1_acquire_bits_header_src = {1{$random}};
    assign memArb.io_in_1_acquire_bits_header_dst = {1{$random}};
  `endif
endmodule

module Queue_2(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [1:0] io_enq_bits_client_xact_id,
    input [511:0] io_enq_bits_data,
    input [2:0] io_enq_bits_a_type,
    input [5:0] io_enq_bits_write_mask,
    input [2:0] io_enq_bits_subword_addr,
    input [3:0] io_enq_bits_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[1:0] io_deq_bits_client_xact_id,
    output[511:0] io_deq_bits_data,
    output[2:0] io_deq_bits_a_type,
    output[5:0] io_deq_bits_write_mask,
    output[2:0] io_deq_bits_subword_addr,
    output[3:0] io_deq_bits_atomic_opcode,
    output io_count
);

  wire T0;
  wire[1:0] T1;
  reg  maybe_full;
  wire T2;
  wire T3;
  wire do_enq;
  wire T4;
  wire do_deq;
  wire[3:0] T5;
  wire[555:0] T6;
  reg [555:0] ram [0:0];
  wire[555:0] T7;
  wire[555:0] T8;
  wire[555:0] T9;
  wire[15:0] T10;
  wire[6:0] T11;
  wire[8:0] T12;
  wire[539:0] T13;
  wire[513:0] T14;
  wire[2:0] T15;
  wire[5:0] T16;
  wire[2:0] T17;
  wire[511:0] T18;
  wire[1:0] T19;
  wire[25:0] T20;
  wire T21;
  wire empty;
  wire T22;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {18{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = {maybe_full, 1'h0};
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = T4 ? do_enq : maybe_full;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T4 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_atomic_opcode = T5;
  assign T5 = T6[2'h3:1'h0];
  assign T6 = ram[1'h0];
  assign T8 = T9;
  assign T9 = {T13, T10};
  assign T10 = {T12, T11};
  assign T11 = {io_enq_bits_subword_addr, io_enq_bits_atomic_opcode};
  assign T12 = {io_enq_bits_a_type, io_enq_bits_write_mask};
  assign T13 = {io_enq_bits_addr, T14};
  assign T14 = {io_enq_bits_client_xact_id, io_enq_bits_data};
  assign io_deq_bits_subword_addr = T15;
  assign T15 = T6[3'h6:3'h4];
  assign io_deq_bits_write_mask = T16;
  assign T16 = T6[4'hc:3'h7];
  assign io_deq_bits_a_type = T17;
  assign T17 = T6[4'hf:4'hd];
  assign io_deq_bits_data = T18;
  assign T18 = T6[10'h20f:5'h10];
  assign io_deq_bits_client_xact_id = T19;
  assign T19 = T6[10'h211:10'h210];
  assign io_deq_bits_addr = T20;
  assign T20 = T6[10'h22b:10'h212];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign io_enq_ready = T22;
  assign T22 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T4) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[1'h0] <= T8;
  end
endmodule

module HTIF(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    output io_cpu_0_reset,
    //output io_cpu_0_id
    input  io_cpu_0_pcr_req_ready,
    output io_cpu_0_pcr_req_valid,
    output io_cpu_0_pcr_req_bits_rw,
    output[4:0] io_cpu_0_pcr_req_bits_addr,
    output[63:0] io_cpu_0_pcr_req_bits_data,
    output io_cpu_0_pcr_rep_ready,
    input  io_cpu_0_pcr_rep_valid,
    input [63:0] io_cpu_0_pcr_rep_bits,
    output io_cpu_0_ipi_req_ready,
    input  io_cpu_0_ipi_req_valid,
    input  io_cpu_0_ipi_req_bits,
    input  io_cpu_0_ipi_rep_ready,
    output io_cpu_0_ipi_rep_valid,
    //output io_cpu_0_ipi_rep_bits
    input  io_cpu_0_debug_stats_pcr,
    input  io_mem_acquire_ready,
    output io_mem_acquire_valid,
    output[1:0] io_mem_acquire_bits_header_src,
    output[1:0] io_mem_acquire_bits_header_dst,
    output[25:0] io_mem_acquire_bits_payload_addr,
    output[1:0] io_mem_acquire_bits_payload_client_xact_id,
    output[511:0] io_mem_acquire_bits_payload_data,
    output[2:0] io_mem_acquire_bits_payload_a_type,
    output[5:0] io_mem_acquire_bits_payload_write_mask,
    output[2:0] io_mem_acquire_bits_payload_subword_addr,
    output[3:0] io_mem_acquire_bits_payload_atomic_opcode,
    output io_mem_grant_ready,
    input  io_mem_grant_valid,
    input [1:0] io_mem_grant_bits_header_src,
    input [1:0] io_mem_grant_bits_header_dst,
    input [511:0] io_mem_grant_bits_payload_data,
    input [1:0] io_mem_grant_bits_payload_client_xact_id,
    input [2:0] io_mem_grant_bits_payload_master_xact_id,
    input [3:0] io_mem_grant_bits_payload_g_type,
    input  io_mem_finish_ready,
    output io_mem_finish_valid,
    //output[1:0] io_mem_finish_bits_header_src
    output[1:0] io_mem_finish_bits_header_dst,
    output[2:0] io_mem_finish_bits_payload_master_xact_id,
    output io_mem_probe_ready,
    input  io_mem_probe_valid,
    input [1:0] io_mem_probe_bits_header_src,
    input [1:0] io_mem_probe_bits_header_dst,
    input [25:0] io_mem_probe_bits_payload_addr,
    input [2:0] io_mem_probe_bits_payload_master_xact_id,
    input [1:0] io_mem_probe_bits_payload_p_type,
    input  io_mem_release_ready,
    output io_mem_release_valid,
    //output[1:0] io_mem_release_bits_header_src
    //output[1:0] io_mem_release_bits_header_dst
    output[25:0] io_mem_release_bits_payload_addr,
    output[1:0] io_mem_release_bits_payload_client_xact_id,
    output[2:0] io_mem_release_bits_payload_master_xact_id,
    output[511:0] io_mem_release_bits_payload_data,
    output[2:0] io_mem_release_bits_payload_r_type,
    input [63:0] io_scr_rdata_63,
    input [63:0] io_scr_rdata_62,
    input [63:0] io_scr_rdata_61,
    input [63:0] io_scr_rdata_60,
    input [63:0] io_scr_rdata_59,
    input [63:0] io_scr_rdata_58,
    input [63:0] io_scr_rdata_57,
    input [63:0] io_scr_rdata_56,
    input [63:0] io_scr_rdata_55,
    input [63:0] io_scr_rdata_54,
    input [63:0] io_scr_rdata_53,
    input [63:0] io_scr_rdata_52,
    input [63:0] io_scr_rdata_51,
    input [63:0] io_scr_rdata_50,
    input [63:0] io_scr_rdata_49,
    input [63:0] io_scr_rdata_48,
    input [63:0] io_scr_rdata_47,
    input [63:0] io_scr_rdata_46,
    input [63:0] io_scr_rdata_45,
    input [63:0] io_scr_rdata_44,
    input [63:0] io_scr_rdata_43,
    input [63:0] io_scr_rdata_42,
    input [63:0] io_scr_rdata_41,
    input [63:0] io_scr_rdata_40,
    input [63:0] io_scr_rdata_39,
    input [63:0] io_scr_rdata_38,
    input [63:0] io_scr_rdata_37,
    input [63:0] io_scr_rdata_36,
    input [63:0] io_scr_rdata_35,
    input [63:0] io_scr_rdata_34,
    input [63:0] io_scr_rdata_33,
    input [63:0] io_scr_rdata_32,
    input [63:0] io_scr_rdata_31,
    input [63:0] io_scr_rdata_30,
    input [63:0] io_scr_rdata_29,
    input [63:0] io_scr_rdata_28,
    input [63:0] io_scr_rdata_27,
    input [63:0] io_scr_rdata_26,
    input [63:0] io_scr_rdata_25,
    input [63:0] io_scr_rdata_24,
    input [63:0] io_scr_rdata_23,
    input [63:0] io_scr_rdata_22,
    input [63:0] io_scr_rdata_21,
    input [63:0] io_scr_rdata_20,
    input [63:0] io_scr_rdata_19,
    input [63:0] io_scr_rdata_18,
    input [63:0] io_scr_rdata_17,
    input [63:0] io_scr_rdata_16,
    input [63:0] io_scr_rdata_15,
    input [63:0] io_scr_rdata_14,
    input [63:0] io_scr_rdata_13,
    input [63:0] io_scr_rdata_12,
    input [63:0] io_scr_rdata_11,
    input [63:0] io_scr_rdata_10,
    input [63:0] io_scr_rdata_9,
    input [63:0] io_scr_rdata_8,
    input [63:0] io_scr_rdata_7,
    input [63:0] io_scr_rdata_6,
    input [63:0] io_scr_rdata_5,
    input [63:0] io_scr_rdata_4,
    input [63:0] io_scr_rdata_3,
    input [63:0] io_scr_rdata_2,
    //input [63:0] io_scr_rdata_1
    //input [63:0] io_scr_rdata_0
    output io_scr_wen,
    output[5:0] io_scr_waddr,
    output[63:0] io_scr_wdata
);

  wire[3:0] T0;
  wire[3:0] T1;
  wire[3:0] T2;
  wire T3;
  reg [3:0] cmd;
  wire[3:0] T4;
  wire[3:0] T5;
  wire[63:0] rx_shifter_in;
  wire[47:0] T6;
  reg [63:0] rx_shifter;
  wire[63:0] T7;
  wire T8;
  wire T9;
  wire T10;
  reg [14:0] rx_count;
  wire[14:0] T11;
  wire[14:0] T12;
  wire[14:0] T13;
  wire[14:0] T14;
  wire T15;
  wire T16;
  wire[12:0] T17;
  wire[11:0] tx_size;
  reg [11:0] size;
  wire[11:0] T18;
  wire[11:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire nack;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire bad_mem_packet;
  wire T32;
  wire[2:0] T33;
  reg [39:0] addr;
  wire[39:0] T34;
  wire[39:0] T35;
  wire[39:0] T36;
  wire[39:0] T37;
  wire T38;
  wire T39;
  reg [3:0] state;
  wire[3:0] T40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire[3:0] T43;
  wire[3:0] T44;
  wire[3:0] T45;
  wire[3:0] T46;
  wire[3:0] T47;
  wire[3:0] T48;
  wire[3:0] T49;
  wire[3:0] T50;
  wire[3:0] T51;
  wire[3:0] T52;
  wire[3:0] T53;
  wire[3:0] T54;
  wire T55;
  wire T56;
  wire[3:0] rx_cmd;
  wire T57;
  wire[12:0] rx_word_count;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire rx_done;
  wire T62;
  wire T63;
  wire T64;
  wire[2:0] T65;
  wire T66;
  wire[12:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire rx_word_done;
  wire T72;
  wire[1:0] T73;
  wire T74;
  wire T75;
  wire acq_q_io_enq_ready;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  reg  mem_acked;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire[3:0] T87;
  wire T88;
  wire T89;
  reg [8:0] pos;
  wire[8:0] T90;
  wire[8:0] T91;
  wire[8:0] T92;
  wire[8:0] T93;
  wire T94;
  wire[3:0] T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire tx_done;
  wire T100;
  wire T101;
  wire T102;
  wire[2:0] packet_ram_raddr;
  wire[2:0] T103;
  wire[12:0] T104;
  reg [14:0] tx_count;
  wire[14:0] T105;
  wire[14:0] T106;
  wire[14:0] T107;
  wire[14:0] T108;
  wire T109;
  wire T110;
  wire T111;
  wire[12:0] T112;
  wire T113;
  wire T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire[4:0] T120;
  wire T121;
  wire T122;
  wire[1:0] T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[2:0] T129;
  wire T130;
  wire T131;
  wire T132;
  wire[2:0] T133;
  wire[2:0] T134;
  wire[2:0] T135;
  wire[5:0] T136;
  wire[5:0] T137;
  wire[5:0] T138;
  wire[2:0] T139;
  wire[2:0] T140;
  wire[2:0] T141;
  wire[511:0] T142;
  wire[511:0] T143;
  wire[511:0] T144;
  wire[1:0] T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire[25:0] T150;
  wire[36:0] init_addr;
  wire[39:0] T151;
  wire[25:0] T152;
  wire[25:0] T153;
  wire T154;
  wire T155;
  wire T156;
  wire[63:0] T157;
  reg [63:0] packet_ram [7:0];
  wire[63:0] T158;
  wire[63:0] T159;
  wire T160;
  wire T161;
  wire[63:0] T162;
  wire[63:0] T163;
  wire T164;
  wire T165;
  wire[63:0] T166;
  wire[63:0] T167;
  wire T168;
  wire T169;
  wire[63:0] T170;
  wire[63:0] T171;
  wire T172;
  wire T173;
  wire[63:0] T174;
  wire[63:0] T175;
  wire T176;
  wire T177;
  wire[63:0] T178;
  wire[63:0] T179;
  wire T180;
  wire T181;
  wire[63:0] T182;
  wire[63:0] T183;
  wire T184;
  wire T185;
  wire[63:0] T186;
  wire[63:0] T187;
  wire T188;
  wire T189;
  wire[63:0] T190;
  wire T191;
  wire[2:0] T192;
  wire[2:0] T193;
  wire[5:0] T194;
  wire[5:0] T195;
  wire T196;
  wire T197;
  reg [2:0] mem_gxid;
  wire[2:0] T198;
  reg [1:0] mem_gsrc;
  wire[1:0] T199;
  wire T200;
  reg  mem_needs_ack;
  wire T201;
  wire T202;
  wire T203;
  wire[3:0] acq_q_io_deq_bits_atomic_opcode;
  wire[2:0] acq_q_io_deq_bits_subword_addr;
  wire[5:0] acq_q_io_deq_bits_write_mask;
  wire[2:0] acq_q_io_deq_bits_a_type;
  wire[511:0] mem_req_data;
  wire[447:0] T204;
  wire[383:0] T205;
  wire[319:0] T206;
  wire[255:0] T207;
  wire[191:0] T208;
  wire[127:0] T209;
  wire[63:0] T210;
  wire[63:0] T211;
  wire[63:0] T212;
  wire[63:0] T213;
  wire[63:0] T214;
  wire[63:0] T215;
  wire[63:0] T216;
  wire[63:0] T217;
  wire[1:0] acq_q_io_deq_bits_client_xact_id;
  wire[25:0] acq_q_io_deq_bits_addr;
  wire acq_q_io_deq_valid;
  reg  R218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  reg  R229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire[15:0] T235;
  wire[63:0] T236;
  wire[5:0] T237;
  wire[1:0] T238;
  wire[63:0] tx_data;
  wire[63:0] T239;
  wire[63:0] T240;
  reg [63:0] pcrReadData;
  wire[63:0] T241;
  wire[63:0] T242;
  wire[63:0] T243;
  wire[63:0] T244;
  wire[63:0] T245;
  wire[63:0] T246;
  wire[63:0] T247;
  wire[63:0] T248;
  wire[63:0] T249;
  wire[63:0] T250;
  wire[63:0] scr_rdata_0;
  wire[63:0] scr_rdata_1;
  wire T251;
  wire[5:0] T252;
  wire[63:0] T253;
  wire[63:0] scr_rdata_2;
  wire[63:0] scr_rdata_3;
  wire T254;
  wire T255;
  wire[63:0] T256;
  wire[63:0] T257;
  wire[63:0] scr_rdata_4;
  wire[63:0] scr_rdata_5;
  wire T258;
  wire[63:0] T259;
  wire[63:0] scr_rdata_6;
  wire[63:0] scr_rdata_7;
  wire T260;
  wire T261;
  wire T262;
  wire[63:0] T263;
  wire[63:0] T264;
  wire[63:0] T265;
  wire[63:0] scr_rdata_8;
  wire[63:0] scr_rdata_9;
  wire T266;
  wire[63:0] T267;
  wire[63:0] scr_rdata_10;
  wire[63:0] scr_rdata_11;
  wire T268;
  wire T269;
  wire[63:0] T270;
  wire[63:0] T271;
  wire[63:0] scr_rdata_12;
  wire[63:0] scr_rdata_13;
  wire T272;
  wire[63:0] T273;
  wire[63:0] scr_rdata_14;
  wire[63:0] scr_rdata_15;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[63:0] T278;
  wire[63:0] T279;
  wire[63:0] T280;
  wire[63:0] T281;
  wire[63:0] scr_rdata_16;
  wire[63:0] scr_rdata_17;
  wire T282;
  wire[63:0] T283;
  wire[63:0] scr_rdata_18;
  wire[63:0] scr_rdata_19;
  wire T284;
  wire T285;
  wire[63:0] T286;
  wire[63:0] T287;
  wire[63:0] scr_rdata_20;
  wire[63:0] scr_rdata_21;
  wire T288;
  wire[63:0] T289;
  wire[63:0] scr_rdata_22;
  wire[63:0] scr_rdata_23;
  wire T290;
  wire T291;
  wire T292;
  wire[63:0] T293;
  wire[63:0] T294;
  wire[63:0] T295;
  wire[63:0] scr_rdata_24;
  wire[63:0] scr_rdata_25;
  wire T296;
  wire[63:0] T297;
  wire[63:0] scr_rdata_26;
  wire[63:0] scr_rdata_27;
  wire T298;
  wire T299;
  wire[63:0] T300;
  wire[63:0] T301;
  wire[63:0] scr_rdata_28;
  wire[63:0] scr_rdata_29;
  wire T302;
  wire[63:0] T303;
  wire[63:0] scr_rdata_30;
  wire[63:0] scr_rdata_31;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire[63:0] T309;
  wire[63:0] T310;
  wire[63:0] T311;
  wire[63:0] T312;
  wire[63:0] T313;
  wire[63:0] scr_rdata_32;
  wire[63:0] scr_rdata_33;
  wire T314;
  wire[63:0] T315;
  wire[63:0] scr_rdata_34;
  wire[63:0] scr_rdata_35;
  wire T316;
  wire T317;
  wire[63:0] T318;
  wire[63:0] T319;
  wire[63:0] scr_rdata_36;
  wire[63:0] scr_rdata_37;
  wire T320;
  wire[63:0] T321;
  wire[63:0] scr_rdata_38;
  wire[63:0] scr_rdata_39;
  wire T322;
  wire T323;
  wire T324;
  wire[63:0] T325;
  wire[63:0] T326;
  wire[63:0] T327;
  wire[63:0] scr_rdata_40;
  wire[63:0] scr_rdata_41;
  wire T328;
  wire[63:0] T329;
  wire[63:0] scr_rdata_42;
  wire[63:0] scr_rdata_43;
  wire T330;
  wire T331;
  wire[63:0] T332;
  wire[63:0] T333;
  wire[63:0] scr_rdata_44;
  wire[63:0] scr_rdata_45;
  wire T334;
  wire[63:0] T335;
  wire[63:0] scr_rdata_46;
  wire[63:0] scr_rdata_47;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire[63:0] T340;
  wire[63:0] T341;
  wire[63:0] T342;
  wire[63:0] T343;
  wire[63:0] scr_rdata_48;
  wire[63:0] scr_rdata_49;
  wire T344;
  wire[63:0] T345;
  wire[63:0] scr_rdata_50;
  wire[63:0] scr_rdata_51;
  wire T346;
  wire T347;
  wire[63:0] T348;
  wire[63:0] T349;
  wire[63:0] scr_rdata_52;
  wire[63:0] scr_rdata_53;
  wire T350;
  wire[63:0] T351;
  wire[63:0] scr_rdata_54;
  wire[63:0] scr_rdata_55;
  wire T352;
  wire T353;
  wire T354;
  wire[63:0] T355;
  wire[63:0] T356;
  wire[63:0] T357;
  wire[63:0] scr_rdata_56;
  wire[63:0] scr_rdata_57;
  wire T358;
  wire[63:0] T359;
  wire[63:0] scr_rdata_58;
  wire[63:0] scr_rdata_59;
  wire T360;
  wire T361;
  wire[63:0] T362;
  wire[63:0] T363;
  wire[63:0] scr_rdata_60;
  wire[63:0] scr_rdata_61;
  wire T364;
  wire[63:0] T365;
  wire[63:0] scr_rdata_62;
  wire[63:0] scr_rdata_63;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire[63:0] tx_header;
  wire[15:0] T375;
  wire[3:0] tx_cmd_ext;
  wire[2:0] tx_cmd;
  wire[47:0] T376;
  reg [7:0] seqno;
  wire[7:0] T377;
  wire[7:0] T378;
  wire T379;
  wire T380;
  wire T381;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    cmd = {1{$random}};
    rx_shifter = {2{$random}};
    rx_count = {1{$random}};
    size = {1{$random}};
    addr = {2{$random}};
    state = {1{$random}};
    mem_acked = {1{$random}};
    pos = {1{$random}};
    tx_count = {1{$random}};
    for (initvar = 0; initvar < 8; initvar = initvar+1)
      packet_ram[initvar] = {2{$random}};
    mem_gxid = {1{$random}};
    mem_gsrc = {1{$random}};
    mem_needs_ack = {1{$random}};
    R218 = {1{$random}};
    R229 = {1{$random}};
    pcrReadData = {2{$random}};
    seqno = {1{$random}};
  end
`endif

  assign T0 = T3 ? T2 : T1;
  assign T1 = 4'h0;
  assign T2 = 4'h0;
  assign T3 = cmd == 4'h1;
  assign T4 = T9 ? T5 : cmd;
  assign T5 = rx_shifter_in[2'h3:1'h0];
  assign rx_shifter_in = {io_host_in_bits, T6};
  assign T6 = rx_shifter[6'h3f:5'h10];
  assign T7 = T8 ? rx_shifter_in : rx_shifter;
  assign T8 = io_host_in_valid & io_host_in_ready;
  assign T9 = T8 & T10;
  assign T10 = rx_count == 15'h3;
  assign T11 = reset ? 15'h0 : T12;
  assign T12 = T15 ? 15'h0 : T13;
  assign T13 = T8 ? T14 : rx_count;
  assign T14 = rx_count + 15'h1;
  assign T15 = T99 & T16;
  assign T16 = T104 == T17;
  assign T17 = {1'h0, tx_size};
  assign tx_size = T20 ? size : 12'h0;
  assign T18 = T9 ? T19 : size;
  assign T19 = rx_shifter_in[4'hf:3'h4];
  assign T20 = T26 & T21;
  assign T21 = T23 | T22;
  assign T22 = cmd == 4'h3;
  assign T23 = T25 | T24;
  assign T24 = cmd == 4'h2;
  assign T25 = cmd == 4'h0;
  assign T26 = nack ^ 1'h1;
  assign nack = T130 ? bad_mem_packet : T27;
  assign T27 = T29 ? T28 : 1'h1;
  assign T28 = size != 12'h1;
  assign T29 = T31 | T30;
  assign T30 = cmd == 4'h3;
  assign T31 = cmd == 4'h2;
  assign bad_mem_packet = T128 | T32;
  assign T32 = T33 != 3'h0;
  assign T33 = addr[2'h2:1'h0];
  assign T34 = T38 ? T37 : T35;
  assign T35 = T9 ? T36 : addr;
  assign T36 = rx_shifter_in[6'h3f:5'h18];
  assign T37 = addr + 40'h8;
  assign T38 = T39 & io_mem_finish_ready;
  assign T39 = state == 4'h7;
  assign T40 = reset ? 4'h0 : T41;
  assign T41 = T125 ? 4'h8 : T42;
  assign T42 = io_cpu_0_pcr_rep_valid ? 4'h8 : T43;
  assign T43 = T118 ? 4'h8 : T44;
  assign T44 = T117 ? 4'h2 : T45;
  assign T45 = T99 ? T95 : T46;
  assign T46 = T38 ? T87 : T47;
  assign T47 = T86 ? 4'h7 : T48;
  assign T48 = T79 ? 4'h7 : T49;
  assign T49 = T77 ? 4'h5 : T50;
  assign T50 = T75 ? 4'h6 : T51;
  assign T51 = T61 ? T52 : state;
  assign T52 = T60 ? 4'h3 : T53;
  assign T53 = T59 ? 4'h4 : T54;
  assign T54 = T55 ? 4'h1 : 4'h8;
  assign T55 = T58 | T56;
  assign T56 = rx_cmd == 4'h3;
  assign rx_cmd = T57 ? T5 : cmd;
  assign T57 = rx_word_count == 13'h0;
  assign rx_word_count = rx_count >> 2'h2;
  assign T58 = rx_cmd == 4'h2;
  assign T59 = rx_cmd == 4'h1;
  assign T60 = rx_cmd == 4'h0;
  assign T61 = T74 & rx_done;
  assign rx_done = rx_word_done & T62;
  assign T62 = T71 ? T68 : T63;
  assign T63 = T66 | T64;
  assign T64 = T65 == 3'h0;
  assign T65 = rx_word_count[2'h2:1'h0];
  assign T66 = rx_word_count == T67;
  assign T67 = {1'h0, size};
  assign T68 = T70 & T69;
  assign T69 = T5 != 4'h3;
  assign T70 = T5 != 4'h1;
  assign T71 = rx_word_count == 13'h0;
  assign rx_word_done = io_host_in_valid & T72;
  assign T72 = T73 == 2'h3;
  assign T73 = rx_count[1'h1:1'h0];
  assign T74 = state == 4'h0;
  assign T75 = T76 & acq_q_io_enq_ready;
  assign T76 = state == 4'h4;
  assign T77 = T78 & acq_q_io_enq_ready;
  assign T78 = state == 4'h3;
  assign T79 = T85 & mem_acked;
  assign T80 = reset ? 1'h0 : T81;
  assign T81 = T84 ? 1'h0 : T82;
  assign T82 = T79 ? 1'h0 : T83;
  assign T83 = io_mem_grant_valid ? 1'h1 : mem_acked;
  assign T84 = state == 4'h5;
  assign T85 = state == 4'h6;
  assign T86 = T84 & io_mem_grant_valid;
  assign T87 = T88 ? 4'h8 : 4'h0;
  assign T88 = T94 | T89;
  assign T89 = pos == 9'h1;
  assign T90 = T38 ? T93 : T91;
  assign T91 = T9 ? T92 : pos;
  assign T92 = rx_shifter_in[4'hf:3'h7];
  assign T93 = pos - 9'h1;
  assign T94 = cmd == 4'h0;
  assign T95 = T96 ? 4'h3 : 4'h0;
  assign T96 = T98 & T97;
  assign T97 = pos != 9'h0;
  assign T98 = cmd == 4'h0;
  assign T99 = T116 & tx_done;
  assign tx_done = T113 & T100;
  assign T100 = T111 | T101;
  assign T101 = T110 & T102;
  assign T102 = packet_ram_raddr == 3'h7;
  assign packet_ram_raddr = T103 - 3'h1;
  assign T103 = T104[2'h2:1'h0];
  assign T104 = tx_count[4'he:2'h2];
  assign T105 = reset ? 15'h0 : T106;
  assign T106 = T15 ? 15'h0 : T107;
  assign T107 = T109 ? T108 : tx_count;
  assign T108 = tx_count + 15'h1;
  assign T109 = io_host_out_valid & io_host_out_ready;
  assign T110 = 13'h0 < T104;
  assign T111 = T104 == T112;
  assign T112 = {1'h0, tx_size};
  assign T113 = io_host_out_ready & T114;
  assign T114 = T115 == 2'h3;
  assign T115 = tx_count[1'h1:1'h0];
  assign T116 = state == 4'h8;
  assign T117 = io_cpu_0_pcr_req_valid & io_cpu_0_pcr_req_ready;
  assign T118 = T121 & T119;
  assign T119 = T120 == 5'h1d;
  assign T120 = addr[3'h4:1'h0];
  assign T121 = T124 & T122;
  assign T122 = T123 == 2'h0;
  assign T123 = addr[5'h15:5'h14];
  assign T124 = state == 4'h1;
  assign T125 = T127 & T126;
  assign T126 = T123 == 2'h3;
  assign T127 = state == 4'h1;
  assign T128 = T129 != 3'h0;
  assign T129 = size[2'h2:1'h0];
  assign T130 = T132 | T131;
  assign T131 = cmd == 4'h1;
  assign T132 = cmd == 4'h0;
  assign T133 = T3 ? T135 : T134;
  assign T134 = 3'h0;
  assign T135 = 3'h0;
  assign T136 = T3 ? T138 : T137;
  assign T137 = 6'h0;
  assign T138 = 6'h0;
  assign T139 = T3 ? T141 : T140;
  assign T140 = 3'h2;
  assign T141 = 3'h3;
  assign T142 = T3 ? T144 : T143;
  assign T143 = 512'h0;
  assign T144 = 512'h0;
  assign T145 = T3 ? T147 : T146;
  assign T146 = 2'h0;
  assign T147 = 2'h0;
  assign T148 = T3 ? T152 : T149;
  assign T149 = T150;
  assign T150 = init_addr[5'h19:1'h0];
  assign init_addr = T151 >> 2'h3;
  assign T151 = addr;
  assign T152 = T153;
  assign T153 = init_addr[5'h19:1'h0];
  assign T154 = T156 | T155;
  assign T155 = state == 4'h4;
  assign T156 = state == 4'h3;
  assign io_scr_wdata = T157;
  assign T157 = packet_ram[3'h0];
  assign T159 = io_mem_grant_bits_payload_data[9'h1ff:9'h1c0];
  assign T160 = T161 & io_mem_grant_valid;
  assign T161 = state == 4'h5;
  assign T163 = io_mem_grant_bits_payload_data[9'h1bf:9'h180];
  assign T164 = T165 & io_mem_grant_valid;
  assign T165 = state == 4'h5;
  assign T167 = io_mem_grant_bits_payload_data[9'h17f:9'h140];
  assign T168 = T169 & io_mem_grant_valid;
  assign T169 = state == 4'h5;
  assign T171 = io_mem_grant_bits_payload_data[9'h13f:9'h100];
  assign T172 = T173 & io_mem_grant_valid;
  assign T173 = state == 4'h5;
  assign T175 = io_mem_grant_bits_payload_data[8'hff:8'hc0];
  assign T176 = T177 & io_mem_grant_valid;
  assign T177 = state == 4'h5;
  assign T179 = io_mem_grant_bits_payload_data[8'hbf:8'h80];
  assign T180 = T181 & io_mem_grant_valid;
  assign T181 = state == 4'h5;
  assign T183 = io_mem_grant_bits_payload_data[7'h7f:7'h40];
  assign T184 = T185 & io_mem_grant_valid;
  assign T185 = state == 4'h5;
  assign T187 = io_mem_grant_bits_payload_data[6'h3f:1'h0];
  assign T188 = T189 & io_mem_grant_valid;
  assign T189 = state == 4'h5;
  assign T191 = rx_word_done & io_host_in_ready;
  assign T192 = T193 - 3'h1;
  assign T193 = rx_word_count[2'h2:1'h0];
  assign io_scr_waddr = T194;
  assign T194 = T195;
  assign T195 = addr[3'h5:1'h0];
  assign io_scr_wen = T196;
  assign T196 = T125 ? T197 : 1'h0;
  assign T197 = cmd == 4'h3;
  assign io_mem_release_valid = 1'h0;
  assign io_mem_probe_ready = 1'h0;
  assign io_mem_finish_bits_payload_master_xact_id = mem_gxid;
  assign T198 = io_mem_grant_valid ? io_mem_grant_bits_payload_master_xact_id : mem_gxid;
  assign io_mem_finish_bits_header_dst = mem_gsrc;
  assign T199 = io_mem_grant_valid ? io_mem_grant_bits_header_src : mem_gsrc;
  assign io_mem_finish_valid = T200;
  assign T200 = T203 & mem_needs_ack;
  assign T201 = io_mem_grant_valid ? T202 : mem_needs_ack;
  assign T202 = io_mem_grant_bits_payload_g_type != 4'h0;
  assign T203 = state == 4'h7;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_acquire_bits_payload_atomic_opcode = acq_q_io_deq_bits_atomic_opcode;
  assign io_mem_acquire_bits_payload_subword_addr = acq_q_io_deq_bits_subword_addr;
  assign io_mem_acquire_bits_payload_write_mask = acq_q_io_deq_bits_write_mask;
  assign io_mem_acquire_bits_payload_a_type = acq_q_io_deq_bits_a_type;
  assign io_mem_acquire_bits_payload_data = mem_req_data;
  assign mem_req_data = {T217, T204};
  assign T204 = {T216, T205};
  assign T205 = {T215, T206};
  assign T206 = {T214, T207};
  assign T207 = {T213, T208};
  assign T208 = {T212, T209};
  assign T209 = {T211, T210};
  assign T210 = packet_ram[3'h0];
  assign T211 = packet_ram[3'h1];
  assign T212 = packet_ram[3'h2];
  assign T213 = packet_ram[3'h3];
  assign T214 = packet_ram[3'h4];
  assign T215 = packet_ram[3'h5];
  assign T216 = packet_ram[3'h6];
  assign T217 = packet_ram[3'h7];
  assign io_mem_acquire_bits_payload_client_xact_id = acq_q_io_deq_bits_client_xact_id;
  assign io_mem_acquire_bits_payload_addr = acq_q_io_deq_bits_addr;
  assign io_mem_acquire_bits_header_dst = 2'h0;
  assign io_mem_acquire_bits_header_src = 2'h2;
  assign io_mem_acquire_valid = acq_q_io_deq_valid;
  assign io_cpu_0_ipi_rep_valid = R218;
  assign T219 = reset ? 1'h0 : T220;
  assign T220 = T222 ? 1'h1 : T221;
  assign T221 = io_cpu_0_ipi_rep_ready ? 1'h0 : R218;
  assign T222 = io_cpu_0_ipi_req_valid & T223;
  assign T223 = io_cpu_0_ipi_req_bits == 1'h0;
  assign io_cpu_0_ipi_req_ready = 1'h1;
  assign io_cpu_0_pcr_rep_ready = 1'h1;
  assign io_cpu_0_pcr_req_bits_data = T157;
  assign io_cpu_0_pcr_req_bits_addr = T120;
  assign io_cpu_0_pcr_req_bits_rw = T224;
  assign T224 = cmd == 4'h3;
  assign io_cpu_0_pcr_req_valid = T225;
  assign T225 = T227 & T226;
  assign T226 = T120 != 5'h1d;
  assign T227 = T228 & T122;
  assign T228 = state == 4'h1;
  assign io_cpu_0_reset = R229;
  assign T230 = reset ? 1'h1 : T231;
  assign T231 = T233 ? T232 : R229;
  assign T232 = T157[1'h0:1'h0];
  assign T233 = T118 & T234;
  assign T234 = cmd == 4'h3;
  assign io_host_debug_stats_pcr = io_cpu_0_debug_stats_pcr;
  assign io_host_out_bits = T235;
  assign T235 = T236[4'hf:1'h0];
  assign T236 = tx_data >> T237;
  assign T237 = {T238, 4'h0};
  assign T238 = tx_count[1'h1:1'h0];
  assign tx_data = T379 ? tx_header : T239;
  assign T239 = T372 ? pcrReadData : T240;
  assign T240 = packet_ram[packet_ram_raddr];
  assign T241 = T125 ? T245 : T242;
  assign T242 = io_cpu_0_pcr_rep_valid ? io_cpu_0_pcr_rep_bits : T243;
  assign T243 = T118 ? T244 : pcrReadData;
  assign T244 = {63'h0, R229};
  assign T245 = T371 ? T309 : T246;
  assign T246 = T308 ? T278 : T247;
  assign T247 = T277 ? T263 : T248;
  assign T248 = T262 ? T256 : T249;
  assign T249 = T255 ? T253 : T250;
  assign T250 = T251 ? scr_rdata_1 : scr_rdata_0;
  assign scr_rdata_0 = 64'h1;
  assign scr_rdata_1 = 64'h1000;
  assign T251 = T252[1'h0:1'h0];
  assign T252 = T195;
  assign T253 = T254 ? scr_rdata_3 : scr_rdata_2;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign T254 = T252[1'h0:1'h0];
  assign T255 = T252[1'h1:1'h1];
  assign T256 = T261 ? T259 : T257;
  assign T257 = T258 ? scr_rdata_5 : scr_rdata_4;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign T258 = T252[1'h0:1'h0];
  assign T259 = T260 ? scr_rdata_7 : scr_rdata_6;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign T260 = T252[1'h0:1'h0];
  assign T261 = T252[1'h1:1'h1];
  assign T262 = T252[2'h2:2'h2];
  assign T263 = T276 ? T270 : T264;
  assign T264 = T269 ? T267 : T265;
  assign T265 = T266 ? scr_rdata_9 : scr_rdata_8;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign T266 = T252[1'h0:1'h0];
  assign T267 = T268 ? scr_rdata_11 : scr_rdata_10;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign T268 = T252[1'h0:1'h0];
  assign T269 = T252[1'h1:1'h1];
  assign T270 = T275 ? T273 : T271;
  assign T271 = T272 ? scr_rdata_13 : scr_rdata_12;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign T272 = T252[1'h0:1'h0];
  assign T273 = T274 ? scr_rdata_15 : scr_rdata_14;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign T274 = T252[1'h0:1'h0];
  assign T275 = T252[1'h1:1'h1];
  assign T276 = T252[2'h2:2'h2];
  assign T277 = T252[2'h3:2'h3];
  assign T278 = T307 ? T293 : T279;
  assign T279 = T292 ? T286 : T280;
  assign T280 = T285 ? T283 : T281;
  assign T281 = T282 ? scr_rdata_17 : scr_rdata_16;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign T282 = T252[1'h0:1'h0];
  assign T283 = T284 ? scr_rdata_19 : scr_rdata_18;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign T284 = T252[1'h0:1'h0];
  assign T285 = T252[1'h1:1'h1];
  assign T286 = T291 ? T289 : T287;
  assign T287 = T288 ? scr_rdata_21 : scr_rdata_20;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign T288 = T252[1'h0:1'h0];
  assign T289 = T290 ? scr_rdata_23 : scr_rdata_22;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign T290 = T252[1'h0:1'h0];
  assign T291 = T252[1'h1:1'h1];
  assign T292 = T252[2'h2:2'h2];
  assign T293 = T306 ? T300 : T294;
  assign T294 = T299 ? T297 : T295;
  assign T295 = T296 ? scr_rdata_25 : scr_rdata_24;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign T296 = T252[1'h0:1'h0];
  assign T297 = T298 ? scr_rdata_27 : scr_rdata_26;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign T298 = T252[1'h0:1'h0];
  assign T299 = T252[1'h1:1'h1];
  assign T300 = T305 ? T303 : T301;
  assign T301 = T302 ? scr_rdata_29 : scr_rdata_28;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign T302 = T252[1'h0:1'h0];
  assign T303 = T304 ? scr_rdata_31 : scr_rdata_30;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign T304 = T252[1'h0:1'h0];
  assign T305 = T252[1'h1:1'h1];
  assign T306 = T252[2'h2:2'h2];
  assign T307 = T252[2'h3:2'h3];
  assign T308 = T252[3'h4:3'h4];
  assign T309 = T370 ? T340 : T310;
  assign T310 = T339 ? T325 : T311;
  assign T311 = T324 ? T318 : T312;
  assign T312 = T317 ? T315 : T313;
  assign T313 = T314 ? scr_rdata_33 : scr_rdata_32;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign T314 = T252[1'h0:1'h0];
  assign T315 = T316 ? scr_rdata_35 : scr_rdata_34;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign T316 = T252[1'h0:1'h0];
  assign T317 = T252[1'h1:1'h1];
  assign T318 = T323 ? T321 : T319;
  assign T319 = T320 ? scr_rdata_37 : scr_rdata_36;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign T320 = T252[1'h0:1'h0];
  assign T321 = T322 ? scr_rdata_39 : scr_rdata_38;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign T322 = T252[1'h0:1'h0];
  assign T323 = T252[1'h1:1'h1];
  assign T324 = T252[2'h2:2'h2];
  assign T325 = T338 ? T332 : T326;
  assign T326 = T331 ? T329 : T327;
  assign T327 = T328 ? scr_rdata_41 : scr_rdata_40;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign T328 = T252[1'h0:1'h0];
  assign T329 = T330 ? scr_rdata_43 : scr_rdata_42;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign T330 = T252[1'h0:1'h0];
  assign T331 = T252[1'h1:1'h1];
  assign T332 = T337 ? T335 : T333;
  assign T333 = T334 ? scr_rdata_45 : scr_rdata_44;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign T334 = T252[1'h0:1'h0];
  assign T335 = T336 ? scr_rdata_47 : scr_rdata_46;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign T336 = T252[1'h0:1'h0];
  assign T337 = T252[1'h1:1'h1];
  assign T338 = T252[2'h2:2'h2];
  assign T339 = T252[2'h3:2'h3];
  assign T340 = T369 ? T355 : T341;
  assign T341 = T354 ? T348 : T342;
  assign T342 = T347 ? T345 : T343;
  assign T343 = T344 ? scr_rdata_49 : scr_rdata_48;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign T344 = T252[1'h0:1'h0];
  assign T345 = T346 ? scr_rdata_51 : scr_rdata_50;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign T346 = T252[1'h0:1'h0];
  assign T347 = T252[1'h1:1'h1];
  assign T348 = T353 ? T351 : T349;
  assign T349 = T350 ? scr_rdata_53 : scr_rdata_52;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign T350 = T252[1'h0:1'h0];
  assign T351 = T352 ? scr_rdata_55 : scr_rdata_54;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign T352 = T252[1'h0:1'h0];
  assign T353 = T252[1'h1:1'h1];
  assign T354 = T252[2'h2:2'h2];
  assign T355 = T368 ? T362 : T356;
  assign T356 = T361 ? T359 : T357;
  assign T357 = T358 ? scr_rdata_57 : scr_rdata_56;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign T358 = T252[1'h0:1'h0];
  assign T359 = T360 ? scr_rdata_59 : scr_rdata_58;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign T360 = T252[1'h0:1'h0];
  assign T361 = T252[1'h1:1'h1];
  assign T362 = T367 ? T365 : T363;
  assign T363 = T364 ? scr_rdata_61 : scr_rdata_60;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign T364 = T252[1'h0:1'h0];
  assign T365 = T366 ? scr_rdata_63 : scr_rdata_62;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T366 = T252[1'h0:1'h0];
  assign T367 = T252[1'h1:1'h1];
  assign T368 = T252[2'h2:2'h2];
  assign T369 = T252[2'h3:2'h3];
  assign T370 = T252[3'h4:3'h4];
  assign T371 = T252[3'h5:3'h5];
  assign T372 = T374 | T373;
  assign T373 = cmd == 4'h3;
  assign T374 = cmd == 4'h2;
  assign tx_header = {T376, T375};
  assign T375 = {tx_size, tx_cmd_ext};
  assign tx_cmd_ext = {1'h0, tx_cmd};
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign T376 = {addr, seqno};
  assign T377 = T9 ? T378 : seqno;
  assign T378 = rx_shifter_in[5'h17:5'h10];
  assign T379 = T104 == 13'h0;
  assign io_host_out_valid = T380;
  assign T380 = state == 4'h8;
  assign io_host_in_ready = T381;
  assign T381 = state == 4'h0;
  Queue_2 acq_q(.clk(clk), .reset(reset),
       .io_enq_ready( acq_q_io_enq_ready ),
       .io_enq_valid( T154 ),
       .io_enq_bits_addr( T148 ),
       .io_enq_bits_client_xact_id( T145 ),
       .io_enq_bits_data( T142 ),
       .io_enq_bits_a_type( T139 ),
       .io_enq_bits_write_mask( T136 ),
       .io_enq_bits_subword_addr( T133 ),
       .io_enq_bits_atomic_opcode( T0 ),
       .io_deq_ready( io_mem_acquire_ready ),
       .io_deq_valid( acq_q_io_deq_valid ),
       .io_deq_bits_addr( acq_q_io_deq_bits_addr ),
       .io_deq_bits_client_xact_id( acq_q_io_deq_bits_client_xact_id ),
       //.io_deq_bits_data(  )
       .io_deq_bits_a_type( acq_q_io_deq_bits_a_type ),
       .io_deq_bits_write_mask( acq_q_io_deq_bits_write_mask ),
       .io_deq_bits_subword_addr( acq_q_io_deq_bits_subword_addr ),
       .io_deq_bits_atomic_opcode( acq_q_io_deq_bits_atomic_opcode )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T9) begin
      cmd <= T5;
    end
    if(T8) begin
      rx_shifter <= rx_shifter_in;
    end
    if(reset) begin
      rx_count <= 15'h0;
    end else if(T15) begin
      rx_count <= 15'h0;
    end else if(T8) begin
      rx_count <= T14;
    end
    if(T9) begin
      size <= T19;
    end
    if(T38) begin
      addr <= T37;
    end else if(T9) begin
      addr <= T36;
    end
    if(reset) begin
      state <= 4'h0;
    end else if(T125) begin
      state <= 4'h8;
    end else if(io_cpu_0_pcr_rep_valid) begin
      state <= 4'h8;
    end else if(T118) begin
      state <= 4'h8;
    end else if(T117) begin
      state <= 4'h2;
    end else if(T99) begin
      state <= T95;
    end else if(T38) begin
      state <= T87;
    end else if(T86) begin
      state <= 4'h7;
    end else if(T79) begin
      state <= 4'h7;
    end else if(T77) begin
      state <= 4'h5;
    end else if(T75) begin
      state <= 4'h6;
    end else if(T61) begin
      state <= T52;
    end
    if(reset) begin
      mem_acked <= 1'h0;
    end else if(T84) begin
      mem_acked <= 1'h0;
    end else if(T79) begin
      mem_acked <= 1'h0;
    end else if(io_mem_grant_valid) begin
      mem_acked <= 1'h1;
    end
    if(T38) begin
      pos <= T93;
    end else if(T9) begin
      pos <= T92;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else if(T15) begin
      tx_count <= 15'h0;
    end else if(T109) begin
      tx_count <= T108;
    end
    if (T160)
      packet_ram[3'h7] <= T159;
    if (T164)
      packet_ram[3'h6] <= T163;
    if (T168)
      packet_ram[3'h5] <= T167;
    if (T172)
      packet_ram[3'h4] <= T171;
    if (T176)
      packet_ram[3'h3] <= T175;
    if (T180)
      packet_ram[3'h2] <= T179;
    if (T184)
      packet_ram[3'h1] <= T183;
    if (T188)
      packet_ram[3'h0] <= T187;
    if (T191)
      packet_ram[T192] <= rx_shifter_in;
    if(io_mem_grant_valid) begin
      mem_gxid <= io_mem_grant_bits_payload_master_xact_id;
    end
    if(io_mem_grant_valid) begin
      mem_gsrc <= io_mem_grant_bits_header_src;
    end
    if(io_mem_grant_valid) begin
      mem_needs_ack <= T202;
    end
    if(reset) begin
      R218 <= 1'h0;
    end else if(T222) begin
      R218 <= 1'h1;
    end else if(io_cpu_0_ipi_rep_ready) begin
      R218 <= 1'h0;
    end
    if(reset) begin
      R229 <= 1'h1;
    end else if(T233) begin
      R229 <= T232;
    end
    if(T125) begin
      pcrReadData <= T245;
    end else if(io_cpu_0_pcr_rep_valid) begin
      pcrReadData <= io_cpu_0_pcr_rep_bits;
    end else if(T118) begin
      pcrReadData <= T244;
    end
    if(T9) begin
      seqno <= T378;
    end
  end
endmodule

module LockingRRArbiter_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[5:0] T20;
  wire[5:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire T27;
  wire[511:0] T28;
  wire[511:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[25:0] T36;
  wire[25:0] T37;
  wire T38;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_atomic_opcode = T11;
  assign T11 = T15 ? io_in_2_bits_payload_atomic_opcode : T12;
  assign T12 = T13 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_subword_addr = T16;
  assign T16 = T19 ? io_in_2_bits_payload_subword_addr : T17;
  assign T17 = T18 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_write_mask = T20;
  assign T20 = T23 ? io_in_2_bits_payload_write_mask : T21;
  assign T21 = T22 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_a_type = T24;
  assign T24 = T27 ? io_in_2_bits_payload_a_type : T25;
  assign T25 = T26 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T28;
  assign T28 = T31 ? io_in_2_bits_payload_data : T29;
  assign T29 = T30 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T32;
  assign T32 = T35 ? io_in_2_bits_payload_client_xact_id : T33;
  assign T33 = T34 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T36;
  assign T36 = T39 ? io_in_2_bits_payload_addr : T37;
  assign T37 = T38 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T40;
  assign T40 = T43 ? io_in_2_bits_header_dst : T41;
  assign T41 = T42 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T42 = T14[1'h0:1'h0];
  assign T43 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T44;
  assign T44 = T47 ? io_in_2_bits_header_src : T45;
  assign T45 = T46 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T46 = T14[1'h0:1'h0];
  assign T47 = T14[1'h1:1'h1];
  assign io_out_valid = T48;
  assign T48 = T51 ? io_in_2_valid : T49;
  assign T49 = T50 ? io_in_1_valid : io_in_0_valid;
  assign T50 = T14[1'h0:1'h0];
  assign T51 = T14[1'h1:1'h1];
  assign io_in_0_ready = T52;
  assign T52 = T53 & io_out_ready;
  assign T53 = T63 | T54;
  assign T54 = T55 ^ 1'h1;
  assign T55 = T58 | T56;
  assign T56 = io_in_2_valid & T57;
  assign T57 = last_grant < 2'h2;
  assign T58 = T61 | T59;
  assign T59 = io_in_1_valid & T60;
  assign T60 = last_grant < 2'h1;
  assign T61 = io_in_0_valid & T62;
  assign T62 = last_grant < 2'h0;
  assign T63 = last_grant < 2'h0;
  assign io_in_1_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T70 | T66;
  assign T66 = T67 ^ 1'h1;
  assign T67 = T68 | io_in_0_valid;
  assign T68 = T69 | T56;
  assign T69 = T61 | T59;
  assign T70 = T72 & T71;
  assign T71 = last_grant < 2'h1;
  assign T72 = T61 ^ 1'h1;
  assign io_in_2_ready = T73;
  assign T73 = T74 & io_out_ready;
  assign T74 = T80 | T75;
  assign T75 = T76 ^ 1'h1;
  assign T76 = T77 | io_in_1_valid;
  assign T77 = T78 | io_in_0_valid;
  assign T78 = T79 | T56;
  assign T79 = T61 | T59;
  assign T80 = T82 & T81;
  assign T81 = last_grant < 2'h2;
  assign T82 = T83 ^ 1'h1;
  assign T83 = T61 | T59;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_0(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_a_type,
    output[5:0] io_out_2_bits_payload_write_mask,
    output[2:0] io_out_2_bits_payload_subword_addr,
    output[3:0] io_out_2_bits_payload_atomic_opcode,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_a_type,
    output[5:0] io_out_1_bits_payload_write_mask,
    output[2:0] io_out_1_bits_payload_subword_addr,
    output[3:0] io_out_1_bits_payload_atomic_opcode,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_a_type,
    output[5:0] io_out_0_bits_payload_write_mask,
    output[2:0] io_out_0_bits_payload_subword_addr,
    output[3:0] io_out_0_bits_payload_atomic_opcode
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_1_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  wire[5:0] LockingRRArbiter_2_io_out_bits_payload_write_mask;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_a_type;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_atomic_opcode = LockingRRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_0_bits_payload_subword_addr = LockingRRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_0_bits_payload_write_mask = LockingRRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_0_bits_payload_a_type = LockingRRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_atomic_opcode = LockingRRArbiter_1_io_out_bits_payload_atomic_opcode;
  assign io_out_1_bits_payload_subword_addr = LockingRRArbiter_1_io_out_bits_payload_subword_addr;
  assign io_out_1_bits_payload_write_mask = LockingRRArbiter_1_io_out_bits_payload_write_mask;
  assign io_out_1_bits_payload_a_type = LockingRRArbiter_1_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_atomic_opcode = LockingRRArbiter_2_io_out_bits_payload_atomic_opcode;
  assign io_out_2_bits_payload_subword_addr = LockingRRArbiter_2_io_out_bits_payload_subword_addr;
  assign io_out_2_bits_payload_write_mask = LockingRRArbiter_2_io_out_bits_payload_write_mask;
  assign io_out_2_bits_payload_a_type = LockingRRArbiter_2_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_0 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_1_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_1_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_1_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_1_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  LockingRRArbiter_0 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_bits_payload_atomic_opcode ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_bits_payload_atomic_opcode ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( LockingRRArbiter_2_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( LockingRRArbiter_2_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( LockingRRArbiter_2_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( LockingRRArbiter_2_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_r_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[511:0] T16;
  wire[511:0] T17;
  wire T18;
  wire T19;
  wire[2:0] T20;
  wire[2:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[25:0] T28;
  wire[25:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_r_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_r_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T16;
  assign T16 = T19 ? io_in_2_bits_payload_data : T17;
  assign T17 = T18 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T20;
  assign T20 = T23 ? io_in_2_bits_payload_master_xact_id : T21;
  assign T21 = T22 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T24;
  assign T24 = T27 ? io_in_2_bits_payload_client_xact_id : T25;
  assign T25 = T26 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T28;
  assign T28 = T31 ? io_in_2_bits_payload_addr : T29;
  assign T29 = T30 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T32;
  assign T32 = T35 ? io_in_2_bits_header_dst : T33;
  assign T33 = T34 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T36;
  assign T36 = T39 ? io_in_2_bits_header_src : T37;
  assign T37 = T38 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_out_valid = T40;
  assign T40 = T43 ? io_in_2_valid : T41;
  assign T41 = T42 ? io_in_1_valid : io_in_0_valid;
  assign T42 = T14[1'h0:1'h0];
  assign T43 = T14[1'h1:1'h1];
  assign io_in_0_ready = T44;
  assign T44 = T45 & io_out_ready;
  assign T45 = T55 | T46;
  assign T46 = T47 ^ 1'h1;
  assign T47 = T50 | T48;
  assign T48 = io_in_2_valid & T49;
  assign T49 = last_grant < 2'h2;
  assign T50 = T53 | T51;
  assign T51 = io_in_1_valid & T52;
  assign T52 = last_grant < 2'h1;
  assign T53 = io_in_0_valid & T54;
  assign T54 = last_grant < 2'h0;
  assign T55 = last_grant < 2'h0;
  assign io_in_1_ready = T56;
  assign T56 = T57 & io_out_ready;
  assign T57 = T62 | T58;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_0_valid;
  assign T60 = T61 | T48;
  assign T61 = T53 | T51;
  assign T62 = T64 & T63;
  assign T63 = last_grant < 2'h1;
  assign T64 = T53 ^ 1'h1;
  assign io_in_2_ready = T65;
  assign T65 = T66 & io_out_ready;
  assign T66 = T72 | T67;
  assign T67 = T68 ^ 1'h1;
  assign T68 = T69 | io_in_1_valid;
  assign T69 = T70 | io_in_0_valid;
  assign T70 = T71 | T48;
  assign T71 = T53 | T51;
  assign T72 = T74 & T73;
  assign T73 = last_grant < 2'h2;
  assign T74 = T75 ^ 1'h1;
  assign T75 = T53 | T51;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_1(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_r_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_r_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_r_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[511:0] io_out_2_bits_payload_data,
    output[2:0] io_out_2_bits_payload_r_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[511:0] io_out_1_bits_payload_data,
    output[2:0] io_out_1_bits_payload_r_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[511:0] io_out_0_bits_payload_data,
    output[2:0] io_out_0_bits_payload_r_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_r_type;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_r_type = LockingRRArbiter_0_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_r_type = LockingRRArbiter_1_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_r_type = LockingRRArbiter_2_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_1 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_0_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_1_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_1 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_r_type( io_in_2_bits_payload_r_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_r_type( io_in_1_bits_payload_r_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_r_type( io_in_0_bits_payload_r_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_r_type( LockingRRArbiter_2_io_out_bits_payload_r_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[1:0] T11;
  wire[1:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[25:0] T20;
  wire[25:0] T21;
  wire T22;
  wire T23;
  wire[1:0] T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_p_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_p_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = T19 ? io_in_2_bits_payload_master_xact_id : T17;
  assign T17 = T18 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_addr = T20;
  assign T20 = T23 ? io_in_2_bits_payload_addr : T21;
  assign T21 = T22 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T24;
  assign T24 = T27 ? io_in_2_bits_header_dst : T25;
  assign T25 = T26 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T28;
  assign T28 = T31 ? io_in_2_bits_header_src : T29;
  assign T29 = T30 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_valid = T32;
  assign T32 = T35 ? io_in_2_valid : T33;
  assign T33 = T34 ? io_in_1_valid : io_in_0_valid;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_in_0_ready = T36;
  assign T36 = T37 & io_out_ready;
  assign T37 = T47 | T38;
  assign T38 = T39 ^ 1'h1;
  assign T39 = T42 | T40;
  assign T40 = io_in_2_valid & T41;
  assign T41 = last_grant < 2'h2;
  assign T42 = T45 | T43;
  assign T43 = io_in_1_valid & T44;
  assign T44 = last_grant < 2'h1;
  assign T45 = io_in_0_valid & T46;
  assign T46 = last_grant < 2'h0;
  assign T47 = last_grant < 2'h0;
  assign io_in_1_ready = T48;
  assign T48 = T49 & io_out_ready;
  assign T49 = T54 | T50;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T52 | io_in_0_valid;
  assign T52 = T53 | T40;
  assign T53 = T45 | T43;
  assign T54 = T56 & T55;
  assign T55 = last_grant < 2'h1;
  assign T56 = T45 ^ 1'h1;
  assign io_in_2_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = T64 | T59;
  assign T59 = T60 ^ 1'h1;
  assign T60 = T61 | io_in_1_valid;
  assign T61 = T62 | io_in_0_valid;
  assign T62 = T63 | T40;
  assign T63 = T45 | T43;
  assign T64 = T66 & T65;
  assign T65 = last_grant < 2'h2;
  assign T66 = T67 ^ 1'h1;
  assign T67 = T45 | T43;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_2(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[25:0] io_out_2_bits_payload_addr,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[1:0] io_out_2_bits_payload_p_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[25:0] io_out_1_bits_payload_addr,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[1:0] io_out_1_bits_payload_p_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[25:0] io_out_0_bits_payload_addr,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[1:0] io_out_0_bits_payload_p_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_p_type;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_p_type;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_1_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_p_type;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[25:0] LockingRRArbiter_2_io_out_bits_payload_addr;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_p_type = LockingRRArbiter_0_io_out_bits_payload_p_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_addr = LockingRRArbiter_0_io_out_bits_payload_addr;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_p_type = LockingRRArbiter_1_io_out_bits_payload_p_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_addr = LockingRRArbiter_1_io_out_bits_payload_addr;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_p_type = LockingRRArbiter_2_io_out_bits_payload_p_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_addr = LockingRRArbiter_2_io_out_bits_payload_addr;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_2 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_0_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_1_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_1_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_2 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( io_in_2_bits_payload_p_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( io_in_1_bits_payload_p_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_bits_payload_addr ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_p_type( io_in_0_bits_payload_p_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( LockingRRArbiter_2_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( LockingRRArbiter_2_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[3:0] T11;
  wire[3:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[511:0] T24;
  wire[511:0] T25;
  wire T26;
  wire T27;
  wire[1:0] T28;
  wire[1:0] T29;
  wire T30;
  wire T31;
  wire[1:0] T32;
  wire[1:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_g_type = T11;
  assign T11 = T15 ? io_in_2_bits_payload_g_type : T12;
  assign T12 = T13 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_payload_master_xact_id = T16;
  assign T16 = T19 ? io_in_2_bits_payload_master_xact_id : T17;
  assign T17 = T18 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_payload_client_xact_id = T20;
  assign T20 = T23 ? io_in_2_bits_payload_client_xact_id : T21;
  assign T21 = T22 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_bits_payload_data = T24;
  assign T24 = T27 ? io_in_2_bits_payload_data : T25;
  assign T25 = T26 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T28;
  assign T28 = T31 ? io_in_2_bits_header_dst : T29;
  assign T29 = T30 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T30 = T14[1'h0:1'h0];
  assign T31 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T32;
  assign T32 = T35 ? io_in_2_bits_header_src : T33;
  assign T33 = T34 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T34 = T14[1'h0:1'h0];
  assign T35 = T14[1'h1:1'h1];
  assign io_out_valid = T36;
  assign T36 = T39 ? io_in_2_valid : T37;
  assign T37 = T38 ? io_in_1_valid : io_in_0_valid;
  assign T38 = T14[1'h0:1'h0];
  assign T39 = T14[1'h1:1'h1];
  assign io_in_0_ready = T40;
  assign T40 = T41 & io_out_ready;
  assign T41 = T51 | T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T46 | T44;
  assign T44 = io_in_2_valid & T45;
  assign T45 = last_grant < 2'h2;
  assign T46 = T49 | T47;
  assign T47 = io_in_1_valid & T48;
  assign T48 = last_grant < 2'h1;
  assign T49 = io_in_0_valid & T50;
  assign T50 = last_grant < 2'h0;
  assign T51 = last_grant < 2'h0;
  assign io_in_1_ready = T52;
  assign T52 = T53 & io_out_ready;
  assign T53 = T58 | T54;
  assign T54 = T55 ^ 1'h1;
  assign T55 = T56 | io_in_0_valid;
  assign T56 = T57 | T44;
  assign T57 = T49 | T47;
  assign T58 = T60 & T59;
  assign T59 = last_grant < 2'h1;
  assign T60 = T49 ^ 1'h1;
  assign io_in_2_ready = T61;
  assign T61 = T62 & io_out_ready;
  assign T62 = T68 | T63;
  assign T63 = T64 ^ 1'h1;
  assign T64 = T65 | io_in_1_valid;
  assign T65 = T66 | io_in_0_valid;
  assign T66 = T67 | T44;
  assign T67 = T49 | T47;
  assign T68 = T70 & T69;
  assign T69 = last_grant < 2'h2;
  assign T70 = T71 ^ 1'h1;
  assign T71 = T49 | T47;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_3(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[511:0] io_out_2_bits_payload_data,
    output[1:0] io_out_2_bits_payload_client_xact_id,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    output[3:0] io_out_2_bits_payload_g_type,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[511:0] io_out_1_bits_payload_data,
    output[1:0] io_out_1_bits_payload_client_xact_id,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    output[3:0] io_out_1_bits_payload_g_type,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[511:0] io_out_0_bits_payload_data,
    output[1:0] io_out_0_bits_payload_client_xact_id,
    output[2:0] io_out_0_bits_payload_master_xact_id,
    output[3:0] io_out_0_bits_payload_g_type
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[3:0] LockingRRArbiter_0_io_out_bits_payload_g_type;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_0_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[3:0] LockingRRArbiter_1_io_out_bits_payload_g_type;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_1_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[3:0] LockingRRArbiter_2_io_out_bits_payload_g_type;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  wire[511:0] LockingRRArbiter_2_io_out_bits_payload_data;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_g_type = LockingRRArbiter_0_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_payload_client_xact_id = LockingRRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_data = LockingRRArbiter_0_io_out_bits_payload_data;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_g_type = LockingRRArbiter_1_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_payload_client_xact_id = LockingRRArbiter_1_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_data = LockingRRArbiter_1_io_out_bits_payload_data;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_g_type = LockingRRArbiter_2_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_payload_client_xact_id = LockingRRArbiter_2_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_data = LockingRRArbiter_2_io_out_bits_payload_data;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_3 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_0_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_1_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_1_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_1_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  LockingRRArbiter_3 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_data( io_in_2_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( io_in_2_bits_payload_g_type ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_data( io_in_1_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( io_in_1_bits_payload_g_type ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_data( io_in_0_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( io_in_0_bits_payload_g_type ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_data( LockingRRArbiter_2_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( LockingRRArbiter_2_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( LockingRRArbiter_2_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
endmodule

module LockingRRArbiter_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_chosen
);

  wire[1:0] T0;
  wire[1:0] choose;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire T5;
  reg [1:0] last_grant;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire[1:0] T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    last_grant = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = choose;
  assign choose = T9 ? 2'h1 : T1;
  assign T1 = T4 ? 2'h2 : T2;
  assign T2 = io_in_0_valid ? 2'h0 : T3;
  assign T3 = io_in_1_valid ? 2'h1 : 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = last_grant < 2'h2;
  assign T6 = reset ? 2'h0 : T7;
  assign T7 = T8 ? T0 : last_grant;
  assign T8 = io_out_ready & io_out_valid;
  assign T9 = io_in_1_valid & T10;
  assign T10 = last_grant < 2'h1;
  assign io_out_bits_payload_master_xact_id = T11;
  assign T11 = T15 ? io_in_2_bits_payload_master_xact_id : T12;
  assign T12 = T13 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = T0;
  assign T15 = T14[1'h1:1'h1];
  assign io_out_bits_header_dst = T16;
  assign T16 = T19 ? io_in_2_bits_header_dst : T17;
  assign T17 = T18 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T18 = T14[1'h0:1'h0];
  assign T19 = T14[1'h1:1'h1];
  assign io_out_bits_header_src = T20;
  assign T20 = T23 ? io_in_2_bits_header_src : T21;
  assign T21 = T22 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T22 = T14[1'h0:1'h0];
  assign T23 = T14[1'h1:1'h1];
  assign io_out_valid = T24;
  assign T24 = T27 ? io_in_2_valid : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T14[1'h0:1'h0];
  assign T27 = T14[1'h1:1'h1];
  assign io_in_0_ready = T28;
  assign T28 = T29 & io_out_ready;
  assign T29 = T39 | T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = T34 | T32;
  assign T32 = io_in_2_valid & T33;
  assign T33 = last_grant < 2'h2;
  assign T34 = T37 | T35;
  assign T35 = io_in_1_valid & T36;
  assign T36 = last_grant < 2'h1;
  assign T37 = io_in_0_valid & T38;
  assign T38 = last_grant < 2'h0;
  assign T39 = last_grant < 2'h0;
  assign io_in_1_ready = T40;
  assign T40 = T41 & io_out_ready;
  assign T41 = T46 | T42;
  assign T42 = T43 ^ 1'h1;
  assign T43 = T44 | io_in_0_valid;
  assign T44 = T45 | T32;
  assign T45 = T37 | T35;
  assign T46 = T48 & T47;
  assign T47 = last_grant < 2'h1;
  assign T48 = T37 ^ 1'h1;
  assign io_in_2_ready = T49;
  assign T49 = T50 & io_out_ready;
  assign T50 = T56 | T51;
  assign T51 = T52 ^ 1'h1;
  assign T52 = T53 | io_in_1_valid;
  assign T53 = T54 | io_in_0_valid;
  assign T54 = T55 | T32;
  assign T55 = T37 | T35;
  assign T56 = T58 & T57;
  assign T57 = last_grant < 2'h2;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T37 | T35;

  always @(posedge clk) begin
    if(reset) begin
      last_grant <= 2'h0;
    end else if(T8) begin
      last_grant <= T0;
    end
  end
endmodule

module BasicCrossbar_4(input clk, input reset,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_2_ready,
    output io_out_2_valid,
    output[1:0] io_out_2_bits_header_src,
    output[1:0] io_out_2_bits_header_dst,
    output[2:0] io_out_2_bits_payload_master_xact_id,
    input  io_out_1_ready,
    output io_out_1_valid,
    output[1:0] io_out_1_bits_header_src,
    output[1:0] io_out_1_bits_header_dst,
    output[2:0] io_out_1_bits_payload_master_xact_id,
    input  io_out_0_ready,
    output io_out_0_valid,
    output[1:0] io_out_0_bits_header_src,
    output[1:0] io_out_0_bits_header_dst,
    output[2:0] io_out_0_bits_payload_master_xact_id
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_0_io_out_bits_header_src;
  wire LockingRRArbiter_0_io_out_valid;
  wire[2:0] LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_1_io_out_bits_header_src;
  wire LockingRRArbiter_1_io_out_valid;
  wire[2:0] LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_dst;
  wire[1:0] LockingRRArbiter_2_io_out_bits_header_src;
  wire LockingRRArbiter_2_io_out_valid;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire LockingRRArbiter_2_io_in_0_ready;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire LockingRRArbiter_1_io_in_0_ready;
  wire T26;
  wire T27;
  wire T28;
  wire LockingRRArbiter_0_io_in_0_ready;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire LockingRRArbiter_2_io_in_1_ready;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire LockingRRArbiter_1_io_in_1_ready;
  wire T37;
  wire T38;
  wire T39;
  wire LockingRRArbiter_0_io_in_1_ready;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire LockingRRArbiter_2_io_in_2_ready;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire LockingRRArbiter_1_io_in_2_ready;
  wire T48;
  wire T49;
  wire T50;
  wire LockingRRArbiter_0_io_in_2_ready;


  assign T0 = io_in_0_valid & T1;
  assign T1 = io_in_0_bits_header_dst == 2'h2;
  assign T2 = io_in_1_valid & T3;
  assign T3 = io_in_1_bits_header_dst == 2'h2;
  assign T4 = io_in_2_valid & T5;
  assign T5 = io_in_2_bits_header_dst == 2'h2;
  assign T6 = io_in_0_valid & T7;
  assign T7 = io_in_0_bits_header_dst == 2'h1;
  assign T8 = io_in_1_valid & T9;
  assign T9 = io_in_1_bits_header_dst == 2'h1;
  assign T10 = io_in_2_valid & T11;
  assign T11 = io_in_2_bits_header_dst == 2'h1;
  assign T12 = io_in_0_valid & T13;
  assign T13 = io_in_0_bits_header_dst == 2'h0;
  assign T14 = io_in_1_valid & T15;
  assign T15 = io_in_1_bits_header_dst == 2'h0;
  assign T16 = io_in_2_valid & T17;
  assign T17 = io_in_2_bits_header_dst == 2'h0;
  assign io_out_0_bits_payload_master_xact_id = LockingRRArbiter_0_io_out_bits_payload_master_xact_id;
  assign io_out_0_bits_header_dst = LockingRRArbiter_0_io_out_bits_header_dst;
  assign io_out_0_bits_header_src = LockingRRArbiter_0_io_out_bits_header_src;
  assign io_out_0_valid = LockingRRArbiter_0_io_out_valid;
  assign io_out_1_bits_payload_master_xact_id = LockingRRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_1_bits_header_dst = LockingRRArbiter_1_io_out_bits_header_dst;
  assign io_out_1_bits_header_src = LockingRRArbiter_1_io_out_bits_header_src;
  assign io_out_1_valid = LockingRRArbiter_1_io_out_valid;
  assign io_out_2_bits_payload_master_xact_id = LockingRRArbiter_2_io_out_bits_payload_master_xact_id;
  assign io_out_2_bits_header_dst = LockingRRArbiter_2_io_out_bits_header_dst;
  assign io_out_2_bits_header_src = LockingRRArbiter_2_io_out_bits_header_src;
  assign io_out_2_valid = LockingRRArbiter_2_io_out_valid;
  assign io_in_0_ready = T18;
  assign T18 = T22 | T19;
  assign T19 = T20;
  assign T20 = LockingRRArbiter_2_io_in_0_ready & T21;
  assign T21 = io_in_0_bits_header_dst == 2'h2;
  assign T22 = T26 | T23;
  assign T23 = T24;
  assign T24 = LockingRRArbiter_1_io_in_0_ready & T25;
  assign T25 = io_in_0_bits_header_dst == 2'h1;
  assign T26 = T27;
  assign T27 = LockingRRArbiter_0_io_in_0_ready & T28;
  assign T28 = io_in_0_bits_header_dst == 2'h0;
  assign io_in_1_ready = T29;
  assign T29 = T33 | T30;
  assign T30 = T31;
  assign T31 = LockingRRArbiter_2_io_in_1_ready & T32;
  assign T32 = io_in_1_bits_header_dst == 2'h2;
  assign T33 = T37 | T34;
  assign T34 = T35;
  assign T35 = LockingRRArbiter_1_io_in_1_ready & T36;
  assign T36 = io_in_1_bits_header_dst == 2'h1;
  assign T37 = T38;
  assign T38 = LockingRRArbiter_0_io_in_1_ready & T39;
  assign T39 = io_in_1_bits_header_dst == 2'h0;
  assign io_in_2_ready = T40;
  assign T40 = T44 | T41;
  assign T41 = T42;
  assign T42 = LockingRRArbiter_2_io_in_2_ready & T43;
  assign T43 = io_in_2_bits_header_dst == 2'h2;
  assign T44 = T48 | T45;
  assign T45 = T46;
  assign T46 = LockingRRArbiter_1_io_in_2_ready & T47;
  assign T47 = io_in_2_bits_header_dst == 2'h1;
  assign T48 = T49;
  assign T49 = LockingRRArbiter_0_io_in_2_ready & T50;
  assign T50 = io_in_2_bits_header_dst == 2'h0;
  LockingRRArbiter_4 LockingRRArbiter_0(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( T16 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( T14 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( T12 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_0_ready ),
       .io_out_valid( LockingRRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_0_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_1(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( T8 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( T6 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_1_ready ),
       .io_out_valid( LockingRRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
  LockingRRArbiter_4 LockingRRArbiter_2(.clk(clk), .reset(reset),
       .io_in_2_ready( LockingRRArbiter_2_io_in_2_ready ),
       .io_in_2_valid( T4 ),
       .io_in_2_bits_header_src( io_in_2_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_bits_payload_master_xact_id ),
       .io_in_1_ready( LockingRRArbiter_2_io_in_1_ready ),
       .io_in_1_valid( T2 ),
       .io_in_1_bits_header_src( io_in_1_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_bits_payload_master_xact_id ),
       .io_in_0_ready( LockingRRArbiter_2_io_in_0_ready ),
       .io_in_0_valid( T0 ),
       .io_in_0_bits_header_src( io_in_0_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_bits_payload_master_xact_id ),
       .io_out_ready( io_out_2_ready ),
       .io_out_valid( LockingRRArbiter_2_io_out_valid ),
       .io_out_bits_header_src( LockingRRArbiter_2_io_out_bits_header_src ),
       .io_out_bits_header_dst( LockingRRArbiter_2_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( LockingRRArbiter_2_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module RocketChipCrossbarNetwork(input clk, input reset,
    output io_clients_1_acquire_ready,
    input  io_clients_1_acquire_valid,
    input [1:0] io_clients_1_acquire_bits_header_src,
    input [1:0] io_clients_1_acquire_bits_header_dst,
    input [25:0] io_clients_1_acquire_bits_payload_addr,
    input [1:0] io_clients_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_1_acquire_bits_payload_data,
    input [2:0] io_clients_1_acquire_bits_payload_a_type,
    input [5:0] io_clients_1_acquire_bits_payload_write_mask,
    input [2:0] io_clients_1_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_1_acquire_bits_payload_atomic_opcode,
    input  io_clients_1_grant_ready,
    output io_clients_1_grant_valid,
    output[1:0] io_clients_1_grant_bits_header_src,
    output[1:0] io_clients_1_grant_bits_header_dst,
    output[511:0] io_clients_1_grant_bits_payload_data,
    output[1:0] io_clients_1_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_1_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_1_grant_bits_payload_g_type,
    output io_clients_1_finish_ready,
    input  io_clients_1_finish_valid,
    input [1:0] io_clients_1_finish_bits_header_src,
    input [1:0] io_clients_1_finish_bits_header_dst,
    input [2:0] io_clients_1_finish_bits_payload_master_xact_id,
    input  io_clients_1_probe_ready,
    output io_clients_1_probe_valid,
    output[1:0] io_clients_1_probe_bits_header_src,
    output[1:0] io_clients_1_probe_bits_header_dst,
    output[25:0] io_clients_1_probe_bits_payload_addr,
    output[2:0] io_clients_1_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_1_probe_bits_payload_p_type,
    output io_clients_1_release_ready,
    input  io_clients_1_release_valid,
    input [1:0] io_clients_1_release_bits_header_src,
    input [1:0] io_clients_1_release_bits_header_dst,
    input [25:0] io_clients_1_release_bits_payload_addr,
    input [1:0] io_clients_1_release_bits_payload_client_xact_id,
    input [2:0] io_clients_1_release_bits_payload_master_xact_id,
    input [511:0] io_clients_1_release_bits_payload_data,
    input [2:0] io_clients_1_release_bits_payload_r_type,
    output io_clients_0_acquire_ready,
    input  io_clients_0_acquire_valid,
    input [1:0] io_clients_0_acquire_bits_header_src,
    input [1:0] io_clients_0_acquire_bits_header_dst,
    input [25:0] io_clients_0_acquire_bits_payload_addr,
    input [1:0] io_clients_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_clients_0_acquire_bits_payload_data,
    input [2:0] io_clients_0_acquire_bits_payload_a_type,
    input [5:0] io_clients_0_acquire_bits_payload_write_mask,
    input [2:0] io_clients_0_acquire_bits_payload_subword_addr,
    input [3:0] io_clients_0_acquire_bits_payload_atomic_opcode,
    input  io_clients_0_grant_ready,
    output io_clients_0_grant_valid,
    output[1:0] io_clients_0_grant_bits_header_src,
    output[1:0] io_clients_0_grant_bits_header_dst,
    output[511:0] io_clients_0_grant_bits_payload_data,
    output[1:0] io_clients_0_grant_bits_payload_client_xact_id,
    output[2:0] io_clients_0_grant_bits_payload_master_xact_id,
    output[3:0] io_clients_0_grant_bits_payload_g_type,
    output io_clients_0_finish_ready,
    input  io_clients_0_finish_valid,
    input [1:0] io_clients_0_finish_bits_header_src,
    input [1:0] io_clients_0_finish_bits_header_dst,
    input [2:0] io_clients_0_finish_bits_payload_master_xact_id,
    input  io_clients_0_probe_ready,
    output io_clients_0_probe_valid,
    output[1:0] io_clients_0_probe_bits_header_src,
    output[1:0] io_clients_0_probe_bits_header_dst,
    output[25:0] io_clients_0_probe_bits_payload_addr,
    output[2:0] io_clients_0_probe_bits_payload_master_xact_id,
    output[1:0] io_clients_0_probe_bits_payload_p_type,
    output io_clients_0_release_ready,
    input  io_clients_0_release_valid,
    input [1:0] io_clients_0_release_bits_header_src,
    input [1:0] io_clients_0_release_bits_header_dst,
    input [25:0] io_clients_0_release_bits_payload_addr,
    input [1:0] io_clients_0_release_bits_payload_client_xact_id,
    input [2:0] io_clients_0_release_bits_payload_master_xact_id,
    input [511:0] io_clients_0_release_bits_payload_data,
    input [2:0] io_clients_0_release_bits_payload_r_type,
    input  io_masters_0_acquire_ready,
    output io_masters_0_acquire_valid,
    output[1:0] io_masters_0_acquire_bits_header_src,
    output[1:0] io_masters_0_acquire_bits_header_dst,
    output[25:0] io_masters_0_acquire_bits_payload_addr,
    output[1:0] io_masters_0_acquire_bits_payload_client_xact_id,
    output[511:0] io_masters_0_acquire_bits_payload_data,
    output[2:0] io_masters_0_acquire_bits_payload_a_type,
    output[5:0] io_masters_0_acquire_bits_payload_write_mask,
    output[2:0] io_masters_0_acquire_bits_payload_subword_addr,
    output[3:0] io_masters_0_acquire_bits_payload_atomic_opcode,
    output io_masters_0_grant_ready,
    input  io_masters_0_grant_valid,
    input [1:0] io_masters_0_grant_bits_header_src,
    input [1:0] io_masters_0_grant_bits_header_dst,
    input [511:0] io_masters_0_grant_bits_payload_data,
    input [1:0] io_masters_0_grant_bits_payload_client_xact_id,
    input [2:0] io_masters_0_grant_bits_payload_master_xact_id,
    input [3:0] io_masters_0_grant_bits_payload_g_type,
    input  io_masters_0_finish_ready,
    output io_masters_0_finish_valid,
    output[1:0] io_masters_0_finish_bits_header_src,
    output[1:0] io_masters_0_finish_bits_header_dst,
    output[2:0] io_masters_0_finish_bits_payload_master_xact_id,
    output io_masters_0_probe_ready,
    input  io_masters_0_probe_valid,
    input [1:0] io_masters_0_probe_bits_header_src,
    input [1:0] io_masters_0_probe_bits_header_dst,
    input [25:0] io_masters_0_probe_bits_payload_addr,
    input [2:0] io_masters_0_probe_bits_payload_master_xact_id,
    input [1:0] io_masters_0_probe_bits_payload_p_type,
    input  io_masters_0_release_ready,
    output io_masters_0_release_valid,
    output[1:0] io_masters_0_release_bits_header_src,
    output[1:0] io_masters_0_release_bits_header_dst,
    output[25:0] io_masters_0_release_bits_payload_addr,
    output[1:0] io_masters_0_release_bits_payload_client_xact_id,
    output[2:0] io_masters_0_release_bits_payload_master_xact_id,
    output[511:0] io_masters_0_release_bits_payload_data,
    output[2:0] io_masters_0_release_bits_payload_r_type
);

  wire T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire T5;
  wire[2:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire T10;
  wire T11;
  wire T12;
  wire[3:0] T13;
  wire[2:0] T14;
  wire[1:0] T15;
  wire[511:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[1:0] T23;
  wire[2:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire[1:0] T28;
  wire T29;
  wire T30;
  wire[2:0] T31;
  wire[511:0] T32;
  wire[2:0] T33;
  wire[1:0] T34;
  wire[25:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire T39;
  wire[2:0] T40;
  wire[511:0] T41;
  wire[2:0] T42;
  wire[1:0] T43;
  wire[25:0] T44;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire[3:0] T50;
  wire[2:0] T51;
  wire[5:0] T52;
  wire[2:0] T53;
  wire[511:0] T54;
  wire[1:0] T55;
  wire[25:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[3:0] T61;
  wire[2:0] T62;
  wire[5:0] T63;
  wire[2:0] T64;
  wire[511:0] T65;
  wire[1:0] T66;
  wire[25:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[2:0] T72;
  wire[2:0] relNet_io_out_0_bits_payload_r_type;
  wire[511:0] T73;
  wire[511:0] relNet_io_out_0_bits_payload_data;
  wire[2:0] T74;
  wire[2:0] relNet_io_out_0_bits_payload_master_xact_id;
  wire[1:0] T75;
  wire[1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire[25:0] T76;
  wire[25:0] relNet_io_out_0_bits_payload_addr;
  wire[1:0] T77;
  wire[1:0] relNet_io_out_0_bits_header_dst;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] relNet_io_out_0_bits_header_src;
  wire T80;
  wire relNet_io_out_0_valid;
  wire T81;
  wire prbNet_io_in_0_ready;
  wire[2:0] T82;
  wire[2:0] ackNet_io_out_0_bits_payload_master_xact_id;
  wire[1:0] T83;
  wire[1:0] ackNet_io_out_0_bits_header_dst;
  wire[1:0] T84;
  wire[1:0] T85;
  wire[1:0] ackNet_io_out_0_bits_header_src;
  wire T86;
  wire ackNet_io_out_0_valid;
  wire T87;
  wire gntNet_io_in_0_ready;
  wire[3:0] T88;
  wire[3:0] acqNet_io_out_0_bits_payload_atomic_opcode;
  wire[2:0] T89;
  wire[2:0] acqNet_io_out_0_bits_payload_subword_addr;
  wire[5:0] T90;
  wire[5:0] acqNet_io_out_0_bits_payload_write_mask;
  wire[2:0] T91;
  wire[2:0] acqNet_io_out_0_bits_payload_a_type;
  wire[511:0] T92;
  wire[511:0] acqNet_io_out_0_bits_payload_data;
  wire[1:0] T93;
  wire[1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire[25:0] T94;
  wire[25:0] acqNet_io_out_0_bits_payload_addr;
  wire[1:0] T95;
  wire[1:0] acqNet_io_out_0_bits_header_dst;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] acqNet_io_out_0_bits_header_src;
  wire T98;
  wire acqNet_io_out_0_valid;
  wire T99;
  wire relNet_io_in_1_ready;
  wire[1:0] T100;
  wire[1:0] prbNet_io_out_1_bits_payload_p_type;
  wire[2:0] T101;
  wire[2:0] prbNet_io_out_1_bits_payload_master_xact_id;
  wire[25:0] T102;
  wire[25:0] prbNet_io_out_1_bits_payload_addr;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] prbNet_io_out_1_bits_header_dst;
  wire[1:0] T105;
  wire[1:0] prbNet_io_out_1_bits_header_src;
  wire T106;
  wire prbNet_io_out_1_valid;
  wire T107;
  wire ackNet_io_in_1_ready;
  wire[3:0] T108;
  wire[3:0] gntNet_io_out_1_bits_payload_g_type;
  wire[2:0] T109;
  wire[2:0] gntNet_io_out_1_bits_payload_master_xact_id;
  wire[1:0] T110;
  wire[1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire[511:0] T111;
  wire[511:0] gntNet_io_out_1_bits_payload_data;
  wire[1:0] T112;
  wire[1:0] T113;
  wire[1:0] gntNet_io_out_1_bits_header_dst;
  wire[1:0] T114;
  wire[1:0] gntNet_io_out_1_bits_header_src;
  wire T115;
  wire gntNet_io_out_1_valid;
  wire T116;
  wire acqNet_io_in_1_ready;
  wire T117;
  wire relNet_io_in_2_ready;
  wire[1:0] T118;
  wire[1:0] prbNet_io_out_2_bits_payload_p_type;
  wire[2:0] T119;
  wire[2:0] prbNet_io_out_2_bits_payload_master_xact_id;
  wire[25:0] T120;
  wire[25:0] prbNet_io_out_2_bits_payload_addr;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] prbNet_io_out_2_bits_header_dst;
  wire[1:0] T123;
  wire[1:0] prbNet_io_out_2_bits_header_src;
  wire T124;
  wire prbNet_io_out_2_valid;
  wire T125;
  wire ackNet_io_in_2_ready;
  wire[3:0] T126;
  wire[3:0] gntNet_io_out_2_bits_payload_g_type;
  wire[2:0] T127;
  wire[2:0] gntNet_io_out_2_bits_payload_master_xact_id;
  wire[1:0] T128;
  wire[1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire[511:0] T129;
  wire[511:0] gntNet_io_out_2_bits_payload_data;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] gntNet_io_out_2_bits_header_dst;
  wire[1:0] T132;
  wire[1:0] gntNet_io_out_2_bits_header_src;
  wire T133;
  wire gntNet_io_out_2_valid;
  wire T134;
  wire acqNet_io_in_2_ready;


  assign T0 = io_masters_0_finish_ready;
  assign T1 = io_clients_0_finish_bits_payload_master_xact_id;
  assign T2 = io_clients_0_finish_bits_header_dst;
  assign T3 = T4;
  assign T4 = io_clients_0_finish_bits_header_src + 2'h1;
  assign T5 = io_clients_0_finish_valid;
  assign T6 = io_clients_1_finish_bits_payload_master_xact_id;
  assign T7 = io_clients_1_finish_bits_header_dst;
  assign T8 = T9;
  assign T9 = io_clients_1_finish_bits_header_src + 2'h1;
  assign T10 = io_clients_1_finish_valid;
  assign T11 = io_clients_0_grant_ready;
  assign T12 = io_clients_1_grant_ready;
  assign T13 = io_masters_0_grant_bits_payload_g_type;
  assign T14 = io_masters_0_grant_bits_payload_master_xact_id;
  assign T15 = io_masters_0_grant_bits_payload_client_xact_id;
  assign T16 = io_masters_0_grant_bits_payload_data;
  assign T17 = T18;
  assign T18 = io_masters_0_grant_bits_header_dst + 2'h1;
  assign T19 = io_masters_0_grant_bits_header_src;
  assign T20 = io_masters_0_grant_valid;
  assign T21 = io_clients_0_probe_ready;
  assign T22 = io_clients_1_probe_ready;
  assign T23 = io_masters_0_probe_bits_payload_p_type;
  assign T24 = io_masters_0_probe_bits_payload_master_xact_id;
  assign T25 = io_masters_0_probe_bits_payload_addr;
  assign T26 = T27;
  assign T27 = io_masters_0_probe_bits_header_dst + 2'h1;
  assign T28 = io_masters_0_probe_bits_header_src;
  assign T29 = io_masters_0_probe_valid;
  assign T30 = io_masters_0_release_ready;
  assign T31 = io_clients_0_release_bits_payload_r_type;
  assign T32 = io_clients_0_release_bits_payload_data;
  assign T33 = io_clients_0_release_bits_payload_master_xact_id;
  assign T34 = io_clients_0_release_bits_payload_client_xact_id;
  assign T35 = io_clients_0_release_bits_payload_addr;
  assign T36 = io_clients_0_release_bits_header_dst;
  assign T37 = T38;
  assign T38 = io_clients_0_release_bits_header_src + 2'h1;
  assign T39 = io_clients_0_release_valid;
  assign T40 = io_clients_1_release_bits_payload_r_type;
  assign T41 = io_clients_1_release_bits_payload_data;
  assign T42 = io_clients_1_release_bits_payload_master_xact_id;
  assign T43 = io_clients_1_release_bits_payload_client_xact_id;
  assign T44 = io_clients_1_release_bits_payload_addr;
  assign T45 = io_clients_1_release_bits_header_dst;
  assign T46 = T47;
  assign T47 = io_clients_1_release_bits_header_src + 2'h1;
  assign T48 = io_clients_1_release_valid;
  assign T49 = io_masters_0_acquire_ready;
  assign T50 = io_clients_0_acquire_bits_payload_atomic_opcode;
  assign T51 = io_clients_0_acquire_bits_payload_subword_addr;
  assign T52 = io_clients_0_acquire_bits_payload_write_mask;
  assign T53 = io_clients_0_acquire_bits_payload_a_type;
  assign T54 = io_clients_0_acquire_bits_payload_data;
  assign T55 = io_clients_0_acquire_bits_payload_client_xact_id;
  assign T56 = io_clients_0_acquire_bits_payload_addr;
  assign T57 = io_clients_0_acquire_bits_header_dst;
  assign T58 = T59;
  assign T59 = io_clients_0_acquire_bits_header_src + 2'h1;
  assign T60 = io_clients_0_acquire_valid;
  assign T61 = io_clients_1_acquire_bits_payload_atomic_opcode;
  assign T62 = io_clients_1_acquire_bits_payload_subword_addr;
  assign T63 = io_clients_1_acquire_bits_payload_write_mask;
  assign T64 = io_clients_1_acquire_bits_payload_a_type;
  assign T65 = io_clients_1_acquire_bits_payload_data;
  assign T66 = io_clients_1_acquire_bits_payload_client_xact_id;
  assign T67 = io_clients_1_acquire_bits_payload_addr;
  assign T68 = io_clients_1_acquire_bits_header_dst;
  assign T69 = T70;
  assign T70 = io_clients_1_acquire_bits_header_src + 2'h1;
  assign T71 = io_clients_1_acquire_valid;
  assign io_masters_0_release_bits_payload_r_type = T72;
  assign T72 = relNet_io_out_0_bits_payload_r_type;
  assign io_masters_0_release_bits_payload_data = T73;
  assign T73 = relNet_io_out_0_bits_payload_data;
  assign io_masters_0_release_bits_payload_master_xact_id = T74;
  assign T74 = relNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_release_bits_payload_client_xact_id = T75;
  assign T75 = relNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_release_bits_payload_addr = T76;
  assign T76 = relNet_io_out_0_bits_payload_addr;
  assign io_masters_0_release_bits_header_dst = T77;
  assign T77 = relNet_io_out_0_bits_header_dst;
  assign io_masters_0_release_bits_header_src = T78;
  assign T78 = T79;
  assign T79 = relNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_release_valid = T80;
  assign T80 = relNet_io_out_0_valid;
  assign io_masters_0_probe_ready = T81;
  assign T81 = prbNet_io_in_0_ready;
  assign io_masters_0_finish_bits_payload_master_xact_id = T82;
  assign T82 = ackNet_io_out_0_bits_payload_master_xact_id;
  assign io_masters_0_finish_bits_header_dst = T83;
  assign T83 = ackNet_io_out_0_bits_header_dst;
  assign io_masters_0_finish_bits_header_src = T84;
  assign T84 = T85;
  assign T85 = ackNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_finish_valid = T86;
  assign T86 = ackNet_io_out_0_valid;
  assign io_masters_0_grant_ready = T87;
  assign T87 = gntNet_io_in_0_ready;
  assign io_masters_0_acquire_bits_payload_atomic_opcode = T88;
  assign T88 = acqNet_io_out_0_bits_payload_atomic_opcode;
  assign io_masters_0_acquire_bits_payload_subword_addr = T89;
  assign T89 = acqNet_io_out_0_bits_payload_subword_addr;
  assign io_masters_0_acquire_bits_payload_write_mask = T90;
  assign T90 = acqNet_io_out_0_bits_payload_write_mask;
  assign io_masters_0_acquire_bits_payload_a_type = T91;
  assign T91 = acqNet_io_out_0_bits_payload_a_type;
  assign io_masters_0_acquire_bits_payload_data = T92;
  assign T92 = acqNet_io_out_0_bits_payload_data;
  assign io_masters_0_acquire_bits_payload_client_xact_id = T93;
  assign T93 = acqNet_io_out_0_bits_payload_client_xact_id;
  assign io_masters_0_acquire_bits_payload_addr = T94;
  assign T94 = acqNet_io_out_0_bits_payload_addr;
  assign io_masters_0_acquire_bits_header_dst = T95;
  assign T95 = acqNet_io_out_0_bits_header_dst;
  assign io_masters_0_acquire_bits_header_src = T96;
  assign T96 = T97;
  assign T97 = acqNet_io_out_0_bits_header_src - 2'h1;
  assign io_masters_0_acquire_valid = T98;
  assign T98 = acqNet_io_out_0_valid;
  assign io_clients_0_release_ready = T99;
  assign T99 = relNet_io_in_1_ready;
  assign io_clients_0_probe_bits_payload_p_type = T100;
  assign T100 = prbNet_io_out_1_bits_payload_p_type;
  assign io_clients_0_probe_bits_payload_master_xact_id = T101;
  assign T101 = prbNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_probe_bits_payload_addr = T102;
  assign T102 = prbNet_io_out_1_bits_payload_addr;
  assign io_clients_0_probe_bits_header_dst = T103;
  assign T103 = T104;
  assign T104 = prbNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_probe_bits_header_src = T105;
  assign T105 = prbNet_io_out_1_bits_header_src;
  assign io_clients_0_probe_valid = T106;
  assign T106 = prbNet_io_out_1_valid;
  assign io_clients_0_finish_ready = T107;
  assign T107 = ackNet_io_in_1_ready;
  assign io_clients_0_grant_bits_payload_g_type = T108;
  assign T108 = gntNet_io_out_1_bits_payload_g_type;
  assign io_clients_0_grant_bits_payload_master_xact_id = T109;
  assign T109 = gntNet_io_out_1_bits_payload_master_xact_id;
  assign io_clients_0_grant_bits_payload_client_xact_id = T110;
  assign T110 = gntNet_io_out_1_bits_payload_client_xact_id;
  assign io_clients_0_grant_bits_payload_data = T111;
  assign T111 = gntNet_io_out_1_bits_payload_data;
  assign io_clients_0_grant_bits_header_dst = T112;
  assign T112 = T113;
  assign T113 = gntNet_io_out_1_bits_header_dst - 2'h1;
  assign io_clients_0_grant_bits_header_src = T114;
  assign T114 = gntNet_io_out_1_bits_header_src;
  assign io_clients_0_grant_valid = T115;
  assign T115 = gntNet_io_out_1_valid;
  assign io_clients_0_acquire_ready = T116;
  assign T116 = acqNet_io_in_1_ready;
  assign io_clients_1_release_ready = T117;
  assign T117 = relNet_io_in_2_ready;
  assign io_clients_1_probe_bits_payload_p_type = T118;
  assign T118 = prbNet_io_out_2_bits_payload_p_type;
  assign io_clients_1_probe_bits_payload_master_xact_id = T119;
  assign T119 = prbNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_probe_bits_payload_addr = T120;
  assign T120 = prbNet_io_out_2_bits_payload_addr;
  assign io_clients_1_probe_bits_header_dst = T121;
  assign T121 = T122;
  assign T122 = prbNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_probe_bits_header_src = T123;
  assign T123 = prbNet_io_out_2_bits_header_src;
  assign io_clients_1_probe_valid = T124;
  assign T124 = prbNet_io_out_2_valid;
  assign io_clients_1_finish_ready = T125;
  assign T125 = ackNet_io_in_2_ready;
  assign io_clients_1_grant_bits_payload_g_type = T126;
  assign T126 = gntNet_io_out_2_bits_payload_g_type;
  assign io_clients_1_grant_bits_payload_master_xact_id = T127;
  assign T127 = gntNet_io_out_2_bits_payload_master_xact_id;
  assign io_clients_1_grant_bits_payload_client_xact_id = T128;
  assign T128 = gntNet_io_out_2_bits_payload_client_xact_id;
  assign io_clients_1_grant_bits_payload_data = T129;
  assign T129 = gntNet_io_out_2_bits_payload_data;
  assign io_clients_1_grant_bits_header_dst = T130;
  assign T130 = T131;
  assign T131 = gntNet_io_out_2_bits_header_dst - 2'h1;
  assign io_clients_1_grant_bits_header_src = T132;
  assign T132 = gntNet_io_out_2_bits_header_src;
  assign io_clients_1_grant_valid = T133;
  assign T133 = gntNet_io_out_2_valid;
  assign io_clients_1_acquire_ready = T134;
  assign T134 = acqNet_io_in_2_ready;
  BasicCrossbar_0 acqNet(.clk(clk), .reset(reset),
       .io_in_2_ready( acqNet_io_in_2_ready ),
       .io_in_2_valid( T71 ),
       .io_in_2_bits_header_src( T69 ),
       .io_in_2_bits_header_dst( T68 ),
       .io_in_2_bits_payload_addr( T67 ),
       .io_in_2_bits_payload_client_xact_id( T66 ),
       .io_in_2_bits_payload_data( T65 ),
       .io_in_2_bits_payload_a_type( T64 ),
       .io_in_2_bits_payload_write_mask( T63 ),
       .io_in_2_bits_payload_subword_addr( T62 ),
       .io_in_2_bits_payload_atomic_opcode( T61 ),
       .io_in_1_ready( acqNet_io_in_1_ready ),
       .io_in_1_valid( T60 ),
       .io_in_1_bits_header_src( T58 ),
       .io_in_1_bits_header_dst( T57 ),
       .io_in_1_bits_payload_addr( T56 ),
       .io_in_1_bits_payload_client_xact_id( T55 ),
       .io_in_1_bits_payload_data( T54 ),
       .io_in_1_bits_payload_a_type( T53 ),
       .io_in_1_bits_payload_write_mask( T52 ),
       .io_in_1_bits_payload_subword_addr( T51 ),
       .io_in_1_bits_payload_atomic_opcode( T50 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_a_type(  )
       //.io_in_0_bits_payload_write_mask(  )
       //.io_in_0_bits_payload_subword_addr(  )
       //.io_in_0_bits_payload_atomic_opcode(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_a_type(  )
       //.io_out_2_bits_payload_write_mask(  )
       //.io_out_2_bits_payload_subword_addr(  )
       //.io_out_2_bits_payload_atomic_opcode(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_a_type(  )
       //.io_out_1_bits_payload_write_mask(  )
       //.io_out_1_bits_payload_subword_addr(  )
       //.io_out_1_bits_payload_atomic_opcode(  )
       .io_out_0_ready( T49 ),
       .io_out_0_valid( acqNet_io_out_0_valid ),
       .io_out_0_bits_header_src( acqNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( acqNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( acqNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( acqNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_data( acqNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_a_type( acqNet_io_out_0_bits_payload_a_type ),
       .io_out_0_bits_payload_write_mask( acqNet_io_out_0_bits_payload_write_mask ),
       .io_out_0_bits_payload_subword_addr( acqNet_io_out_0_bits_payload_subword_addr ),
       .io_out_0_bits_payload_atomic_opcode( acqNet_io_out_0_bits_payload_atomic_opcode )
  );
  `ifndef SYNTHESIS
    assign acqNet.io_in_0_bits_header_src = {1{$random}};
    assign acqNet.io_in_0_bits_header_dst = {1{$random}};
    assign acqNet.io_in_0_bits_payload_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign acqNet.io_in_0_bits_payload_data = {16{$random}};
    assign acqNet.io_in_0_bits_payload_a_type = {1{$random}};
    assign acqNet.io_in_0_bits_payload_write_mask = {1{$random}};
    assign acqNet.io_in_0_bits_payload_subword_addr = {1{$random}};
    assign acqNet.io_in_0_bits_payload_atomic_opcode = {1{$random}};
  `endif
  BasicCrossbar_1 relNet(.clk(clk), .reset(reset),
       .io_in_2_ready( relNet_io_in_2_ready ),
       .io_in_2_valid( T48 ),
       .io_in_2_bits_header_src( T46 ),
       .io_in_2_bits_header_dst( T45 ),
       .io_in_2_bits_payload_addr( T44 ),
       .io_in_2_bits_payload_client_xact_id( T43 ),
       .io_in_2_bits_payload_master_xact_id( T42 ),
       .io_in_2_bits_payload_data( T41 ),
       .io_in_2_bits_payload_r_type( T40 ),
       .io_in_1_ready( relNet_io_in_1_ready ),
       .io_in_1_valid( T39 ),
       .io_in_1_bits_header_src( T37 ),
       .io_in_1_bits_header_dst( T36 ),
       .io_in_1_bits_payload_addr( T35 ),
       .io_in_1_bits_payload_client_xact_id( T34 ),
       .io_in_1_bits_payload_master_xact_id( T33 ),
       .io_in_1_bits_payload_data( T32 ),
       .io_in_1_bits_payload_r_type( T31 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_client_xact_id(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_data(  )
       //.io_in_0_bits_payload_r_type(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_addr(  )
       //.io_out_2_bits_payload_client_xact_id(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       //.io_out_2_bits_payload_data(  )
       //.io_out_2_bits_payload_r_type(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_addr(  )
       //.io_out_1_bits_payload_client_xact_id(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       //.io_out_1_bits_payload_data(  )
       //.io_out_1_bits_payload_r_type(  )
       .io_out_0_ready( T30 ),
       .io_out_0_valid( relNet_io_out_0_valid ),
       .io_out_0_bits_header_src( relNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( relNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_addr( relNet_io_out_0_bits_payload_addr ),
       .io_out_0_bits_payload_client_xact_id( relNet_io_out_0_bits_payload_client_xact_id ),
       .io_out_0_bits_payload_master_xact_id( relNet_io_out_0_bits_payload_master_xact_id ),
       .io_out_0_bits_payload_data( relNet_io_out_0_bits_payload_data ),
       .io_out_0_bits_payload_r_type( relNet_io_out_0_bits_payload_r_type )
  );
  `ifndef SYNTHESIS
    assign relNet.io_in_0_bits_header_src = {1{$random}};
    assign relNet.io_in_0_bits_header_dst = {1{$random}};
    assign relNet.io_in_0_bits_payload_addr = {1{$random}};
    assign relNet.io_in_0_bits_payload_client_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign relNet.io_in_0_bits_payload_data = {16{$random}};
    assign relNet.io_in_0_bits_payload_r_type = {1{$random}};
  `endif
  BasicCrossbar_2 prbNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_addr(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_p_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_addr(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_p_type(  )
       .io_in_0_ready( prbNet_io_in_0_ready ),
       .io_in_0_valid( T29 ),
       .io_in_0_bits_header_src( T28 ),
       .io_in_0_bits_header_dst( T26 ),
       .io_in_0_bits_payload_addr( T25 ),
       .io_in_0_bits_payload_master_xact_id( T24 ),
       .io_in_0_bits_payload_p_type( T23 ),
       .io_out_2_ready( T22 ),
       .io_out_2_valid( prbNet_io_out_2_valid ),
       .io_out_2_bits_header_src( prbNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( prbNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_addr( prbNet_io_out_2_bits_payload_addr ),
       .io_out_2_bits_payload_master_xact_id( prbNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_p_type( prbNet_io_out_2_bits_payload_p_type ),
       .io_out_1_ready( T21 ),
       .io_out_1_valid( prbNet_io_out_1_valid ),
       .io_out_1_bits_header_src( prbNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( prbNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_addr( prbNet_io_out_1_bits_payload_addr ),
       .io_out_1_bits_payload_master_xact_id( prbNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_p_type( prbNet_io_out_1_bits_payload_p_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_addr(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_p_type(  )
  );
  `ifndef SYNTHESIS
    assign prbNet.io_in_2_bits_header_src = {1{$random}};
    assign prbNet.io_in_2_bits_header_dst = {1{$random}};
    assign prbNet.io_in_2_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_2_bits_payload_p_type = {1{$random}};
    assign prbNet.io_in_1_bits_header_src = {1{$random}};
    assign prbNet.io_in_1_bits_header_dst = {1{$random}};
    assign prbNet.io_in_1_bits_payload_addr = {1{$random}};
    assign prbNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign prbNet.io_in_1_bits_payload_p_type = {1{$random}};
  `endif
  BasicCrossbar_3 gntNet(.clk(clk), .reset(reset),
       //.io_in_2_ready(  )
       .io_in_2_valid( 1'h0 ),
       //.io_in_2_bits_header_src(  )
       //.io_in_2_bits_header_dst(  )
       //.io_in_2_bits_payload_data(  )
       //.io_in_2_bits_payload_client_xact_id(  )
       //.io_in_2_bits_payload_master_xact_id(  )
       //.io_in_2_bits_payload_g_type(  )
       //.io_in_1_ready(  )
       .io_in_1_valid( 1'h0 ),
       //.io_in_1_bits_header_src(  )
       //.io_in_1_bits_header_dst(  )
       //.io_in_1_bits_payload_data(  )
       //.io_in_1_bits_payload_client_xact_id(  )
       //.io_in_1_bits_payload_master_xact_id(  )
       //.io_in_1_bits_payload_g_type(  )
       .io_in_0_ready( gntNet_io_in_0_ready ),
       .io_in_0_valid( T20 ),
       .io_in_0_bits_header_src( T19 ),
       .io_in_0_bits_header_dst( T17 ),
       .io_in_0_bits_payload_data( T16 ),
       .io_in_0_bits_payload_client_xact_id( T15 ),
       .io_in_0_bits_payload_master_xact_id( T14 ),
       .io_in_0_bits_payload_g_type( T13 ),
       .io_out_2_ready( T12 ),
       .io_out_2_valid( gntNet_io_out_2_valid ),
       .io_out_2_bits_header_src( gntNet_io_out_2_bits_header_src ),
       .io_out_2_bits_header_dst( gntNet_io_out_2_bits_header_dst ),
       .io_out_2_bits_payload_data( gntNet_io_out_2_bits_payload_data ),
       .io_out_2_bits_payload_client_xact_id( gntNet_io_out_2_bits_payload_client_xact_id ),
       .io_out_2_bits_payload_master_xact_id( gntNet_io_out_2_bits_payload_master_xact_id ),
       .io_out_2_bits_payload_g_type( gntNet_io_out_2_bits_payload_g_type ),
       .io_out_1_ready( T11 ),
       .io_out_1_valid( gntNet_io_out_1_valid ),
       .io_out_1_bits_header_src( gntNet_io_out_1_bits_header_src ),
       .io_out_1_bits_header_dst( gntNet_io_out_1_bits_header_dst ),
       .io_out_1_bits_payload_data( gntNet_io_out_1_bits_payload_data ),
       .io_out_1_bits_payload_client_xact_id( gntNet_io_out_1_bits_payload_client_xact_id ),
       .io_out_1_bits_payload_master_xact_id( gntNet_io_out_1_bits_payload_master_xact_id ),
       .io_out_1_bits_payload_g_type( gntNet_io_out_1_bits_payload_g_type ),
       .io_out_0_ready( 1'h0 )
       //.io_out_0_valid(  )
       //.io_out_0_bits_header_src(  )
       //.io_out_0_bits_header_dst(  )
       //.io_out_0_bits_payload_data(  )
       //.io_out_0_bits_payload_client_xact_id(  )
       //.io_out_0_bits_payload_master_xact_id(  )
       //.io_out_0_bits_payload_g_type(  )
  );
  `ifndef SYNTHESIS
    assign gntNet.io_in_2_bits_header_src = {1{$random}};
    assign gntNet.io_in_2_bits_header_dst = {1{$random}};
    assign gntNet.io_in_2_bits_payload_data = {16{$random}};
    assign gntNet.io_in_2_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_2_bits_payload_g_type = {1{$random}};
    assign gntNet.io_in_1_bits_header_src = {1{$random}};
    assign gntNet.io_in_1_bits_header_dst = {1{$random}};
    assign gntNet.io_in_1_bits_payload_data = {16{$random}};
    assign gntNet.io_in_1_bits_payload_client_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_master_xact_id = {1{$random}};
    assign gntNet.io_in_1_bits_payload_g_type = {1{$random}};
  `endif
  BasicCrossbar_4 ackNet(.clk(clk), .reset(reset),
       .io_in_2_ready( ackNet_io_in_2_ready ),
       .io_in_2_valid( T10 ),
       .io_in_2_bits_header_src( T8 ),
       .io_in_2_bits_header_dst( T7 ),
       .io_in_2_bits_payload_master_xact_id( T6 ),
       .io_in_1_ready( ackNet_io_in_1_ready ),
       .io_in_1_valid( T5 ),
       .io_in_1_bits_header_src( T3 ),
       .io_in_1_bits_header_dst( T2 ),
       .io_in_1_bits_payload_master_xact_id( T1 ),
       //.io_in_0_ready(  )
       .io_in_0_valid( 1'h0 ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       .io_out_2_ready( 1'h0 ),
       //.io_out_2_valid(  )
       //.io_out_2_bits_header_src(  )
       //.io_out_2_bits_header_dst(  )
       //.io_out_2_bits_payload_master_xact_id(  )
       .io_out_1_ready( 1'h0 ),
       //.io_out_1_valid(  )
       //.io_out_1_bits_header_src(  )
       //.io_out_1_bits_header_dst(  )
       //.io_out_1_bits_payload_master_xact_id(  )
       .io_out_0_ready( T0 ),
       .io_out_0_valid( ackNet_io_out_0_valid ),
       .io_out_0_bits_header_src( ackNet_io_out_0_bits_header_src ),
       .io_out_0_bits_header_dst( ackNet_io_out_0_bits_header_dst ),
       .io_out_0_bits_payload_master_xact_id( ackNet_io_out_0_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign ackNet.io_in_0_bits_header_src = {1{$random}};
    assign ackNet.io_in_0_bits_header_dst = {1{$random}};
    assign ackNet.io_in_0_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module VoluntaryReleaseTracker(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    //output[1:0] io_inner_probe_bits_header_src
    //output[1:0] io_inner_probe_bits_header_dst
    //output[25:0] io_inner_probe_bits_payload_addr
    //output[2:0] io_inner_probe_bits_payload_master_xact_id
    //output[1:0] io_inner_probe_bits_payload_p_type
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [1:0] state;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  reg [25:0] xact_addr;
  wire[25:0] T21;
  wire[3:0] T22;
  wire[2:0] T23;
  wire[5:0] T24;
  wire[2:0] T25;
  wire[511:0] T26;
  reg [511:0] xact_data;
  wire[511:0] T27;
  wire[1:0] T28;
  wire[25:0] T29;
  wire[3:0] T30;
  wire[3:0] T31;
  wire T32;
  reg [2:0] xact_r_type;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[1:0] T35;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T36;
  wire[511:0] T37;
  wire[1:0] T38;
  reg  init_client_id;
  wire T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    xact_r_type = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T20 & T1;
  assign T1 = state != 2'h0;
  assign T2 = reset ? 2'h0 : T3;
  assign T3 = T18 ? 2'h0 : T4;
  assign T4 = T16 ? 2'h2 : T5;
  assign T5 = T14 ? T6 : state;
  assign T6 = T7 ? 2'h1 : 2'h2;
  assign T7 = T9 | T8;
  assign T8 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T9 = T11 | T10;
  assign T10 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T11 = T13 | T12;
  assign T12 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T13 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T14 = T15 & io_inner_release_valid;
  assign T15 = 2'h0 == state;
  assign T16 = T17 & io_outer_acquire_ready;
  assign T17 = 2'h1 == state;
  assign T18 = T19 & io_inner_grant_ready;
  assign T19 = 2'h2 == state;
  assign T20 = xact_addr == io_inner_release_bits_payload_addr;
  assign T21 = T14 ? io_inner_release_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = 1'h0;
  assign io_outer_grant_ready = 1'h0;
  assign io_outer_acquire_bits_payload_atomic_opcode = T22;
  assign T22 = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T23;
  assign T23 = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T24;
  assign T24 = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T25;
  assign T25 = 3'h3;
  assign io_outer_acquire_bits_payload_data = T26;
  assign T26 = xact_data;
  assign T27 = T14 ? io_inner_release_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T28;
  assign T28 = 2'h0;
  assign io_outer_acquire_bits_payload_addr = T29;
  assign T29 = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T17;
  assign io_inner_release_ready = T15;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_grant_bits_payload_g_type = T30;
  assign T30 = T31;
  assign T31 = T32 ? 4'h0 : 4'h3;
  assign T32 = xact_r_type == 3'h0;
  assign T33 = T14 ? io_inner_release_bits_payload_r_type : xact_r_type;
  assign io_inner_grant_bits_payload_master_xact_id = T34;
  assign T34 = 3'h0;
  assign io_inner_grant_bits_payload_client_xact_id = T35;
  assign T35 = xact_client_xact_id;
  assign T36 = T14 ? io_inner_release_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T37;
  assign T37 = 512'h0;
  assign io_inner_grant_bits_header_dst = T38;
  assign T38 = {1'h0, init_client_id};
  assign T39 = T40[1'h0:1'h0];
  assign T40 = reset ? 2'h0 : T41;
  assign T41 = T14 ? io_inner_release_bits_header_src : T42;
  assign T42 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T19;
  assign io_inner_acquire_ready = 1'h0;

  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else if(T18) begin
      state <= 2'h0;
    end else if(T16) begin
      state <= 2'h2;
    end else if(T14) begin
      state <= T6;
    end
    if(T14) begin
      xact_addr <= io_inner_release_bits_payload_addr;
    end
    if(T14) begin
      xact_data <= io_inner_release_bits_payload_data;
    end
    if(T14) begin
      xact_r_type <= io_inner_release_bits_payload_r_type;
    end
    if(T14) begin
      xact_client_xact_id <= io_inner_release_bits_payload_client_xact_id;
    end
    init_client_id <= T39;
  end
endmodule

module AcquireTracker_0(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h1;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h1;
  assign outer_write_rel_client_xact_id = 2'h1;
  assign outer_write_acq_client_xact_id = 2'h1;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h1;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h1;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 2'h1;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_1(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h2;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h2;
  assign outer_write_rel_client_xact_id = 2'h2;
  assign outer_write_acq_client_xact_id = 2'h2;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h2;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h2;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 2'h2;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_2(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h3;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h3;
  assign outer_write_rel_client_xact_id = 2'h3;
  assign outer_write_acq_client_xact_id = 2'h3;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h3;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h3;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = io_outer_grant_bits_payload_client_xact_id == 2'h3;
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_3(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[2:0] T173;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h4;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h0;
  assign outer_write_rel_client_xact_id = 2'h0;
  assign outer_write_acq_client_xact_id = 2'h0;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h4;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h4;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = T173 == 3'h4;
  assign T173 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_4(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[2:0] T173;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h5;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h1;
  assign outer_write_rel_client_xact_id = 2'h1;
  assign outer_write_acq_client_xact_id = 2'h1;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h5;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h5;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = T173 == 3'h5;
  assign T173 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_5(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[2:0] T173;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h6;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h2;
  assign outer_write_rel_client_xact_id = 2'h2;
  assign outer_write_acq_client_xact_id = 2'h2;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h6;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h6;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = T173 == 3'h6;
  assign T173 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module AcquireTracker_6(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    //output io_inner_finish_ready
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    //output[1:0] io_outer_acquire_bits_header_dst
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    //output io_outer_finish_valid
    //output[1:0] io_outer_finish_bits_header_src
    //output[1:0] io_outer_finish_bits_header_dst
    //output[2:0] io_outer_finish_bits_payload_master_xact_id
    input [1:0] io_tile_incoherent,
    output io_has_acquire_conflict,
    output io_has_release_conflict
);

  wire T0;
  wire T1;
  reg [2:0] state;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire[1:0] probe_initial_flags;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  reg [2:0] xact_a_type;
  wire[2:0] T27;
  wire pending_outer_write;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  reg  release_count;
  wire T34;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire[1:0] T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[2:0] T62;
  wire[2:0] T63;
  wire T64;
  wire T65;
  wire[2:0] T66;
  wire T67;
  wire[3:0] grant_type;
  wire[3:0] T68;
  wire[3:0] T69;
  wire[3:0] T70;
  wire[3:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  reg  init_sharer_cnt;
  wire T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[2:0] T89;
  wire T90;
  wire T91;
  wire[2:0] T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg [25:0] xact_addr;
  wire[25:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] outer_read_atomic_opcode;
  wire[3:0] outer_write_rel_atomic_opcode;
  wire[3:0] outer_write_acq_atomic_opcode;
  wire[2:0] T108;
  wire[2:0] T109;
  wire[2:0] T110;
  wire[2:0] outer_read_subword_addr;
  wire[2:0] outer_write_rel_subword_addr;
  wire[2:0] outer_write_acq_subword_addr;
  wire[5:0] T111;
  wire[5:0] T112;
  wire[5:0] T113;
  wire[5:0] outer_read_write_mask;
  wire[5:0] outer_write_rel_write_mask;
  wire[5:0] outer_write_acq_write_mask;
  wire[2:0] T114;
  wire[2:0] T115;
  wire[2:0] T116;
  wire[2:0] outer_read_a_type;
  wire[2:0] outer_write_rel_a_type;
  wire[2:0] outer_write_acq_a_type;
  wire[511:0] T117;
  wire[511:0] T118;
  wire[511:0] T119;
  wire[511:0] outer_read_data;
  wire[511:0] outer_write_rel_data;
  wire[511:0] outer_write_acq_data;
  reg [511:0] xact_data;
  wire[511:0] T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire[1:0] T123;
  wire[1:0] outer_read_client_xact_id;
  wire[1:0] outer_write_rel_client_xact_id;
  wire[1:0] outer_write_acq_client_xact_id;
  wire[25:0] T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire[25:0] outer_read_addr;
  wire[25:0] outer_write_rel_addr;
  wire[25:0] outer_write_acq_addr;
  wire T127;
  wire T128;
  wire T129;
  wire[1:0] T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire[1:0] T135;
  wire[1:0] T136;
  wire[1:0] T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire[2:0] T145;
  wire[25:0] T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  reg [1:0] probe_flags;
  wire[1:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire[1:0] T155;
  wire T156;
  wire T157;
  wire T158;
  wire[3:0] T159;
  wire[2:0] T160;
  wire[1:0] T161;
  reg [1:0] xact_client_xact_id;
  wire[1:0] T162;
  wire[511:0] T163;
  wire[1:0] T164;
  reg  init_client_id;
  wire T165;
  wire[1:0] T166;
  wire[1:0] T167;
  wire[1:0] T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire[2:0] T173;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    state = {1{$random}};
    xact_a_type = {1{$random}};
    release_count = {1{$random}};
    init_sharer_cnt = {1{$random}};
    xact_addr = {1{$random}};
    xact_data = {16{$random}};
    probe_flags = {1{$random}};
    xact_client_xact_id = {1{$random}};
    init_client_id = {1{$random}};
  end
`endif

  assign io_has_release_conflict = T0;
  assign T0 = T100 & T1;
  assign T1 = state != 3'h0;
  assign T2 = reset ? 3'h0 : T3;
  assign T3 = T96 ? 3'h0 : T4;
  assign T4 = T94 ? T92 : T5;
  assign T5 = T90 ? T89 : T6;
  assign T6 = T87 ? T66 : T7;
  assign T7 = T64 ? T62 : T8;
  assign T8 = T32 ? T24 : T9;
  assign T9 = T22 ? T10 : state;
  assign T10 = T19 ? 3'h1 : T11;
  assign T11 = T14 ? 3'h3 : T12;
  assign T12 = T13 ? 3'h2 : 3'h4;
  assign T13 = io_inner_acquire_bits_payload_a_type != 3'h3;
  assign T14 = T16 | T15;
  assign T15 = 3'h6 == io_inner_acquire_bits_payload_a_type;
  assign T16 = T18 | T17;
  assign T17 = 3'h5 == io_inner_acquire_bits_payload_a_type;
  assign T18 = 3'h3 == io_inner_acquire_bits_payload_a_type;
  assign T19 = probe_initial_flags != 2'h0;
  assign probe_initial_flags = T20;
  assign T20 = ~ T21;
  assign T21 = io_tile_incoherent | 2'h0;
  assign T22 = T23 & io_inner_acquire_valid;
  assign T23 = 3'h0 == state;
  assign T24 = pending_outer_write ? 3'h3 : T25;
  assign T25 = T26 ? 3'h2 : 3'h4;
  assign T26 = xact_a_type != 3'h3;
  assign T27 = T22 ? io_inner_acquire_bits_payload_a_type : xact_a_type;
  assign pending_outer_write = T29 | T28;
  assign T28 = 3'h6 == xact_a_type;
  assign T29 = T31 | T30;
  assign T30 = 3'h5 == xact_a_type;
  assign T31 = 3'h3 == xact_a_type;
  assign T32 = T47 & T33;
  assign T33 = release_count == 1'h1;
  assign T34 = T35[1'h0:1'h0];
  assign T35 = reset ? 2'h0 : T36;
  assign T36 = T60 ? T58 : T37;
  assign T37 = T47 ? T45 : T38;
  assign T38 = T22 ? T40 : T39;
  assign T39 = {1'h0, release_count};
  assign T40 = T43 + T41;
  assign T41 = {1'h0, T42};
  assign T42 = probe_initial_flags[1'h1:1'h1];
  assign T43 = {1'h0, T44};
  assign T44 = probe_initial_flags[1'h0:1'h0];
  assign T45 = {1'h0, T46};
  assign T46 = release_count - 1'h1;
  assign T47 = T48 & io_outer_acquire_ready;
  assign T48 = T56 & T49;
  assign T49 = T51 | T50;
  assign T50 = 3'h3 == io_inner_release_bits_payload_r_type;
  assign T51 = T53 | T52;
  assign T52 = 3'h2 == io_inner_release_bits_payload_r_type;
  assign T53 = T55 | T54;
  assign T54 = 3'h1 == io_inner_release_bits_payload_r_type;
  assign T55 = 3'h0 == io_inner_release_bits_payload_r_type;
  assign T56 = T57 & io_inner_release_valid;
  assign T57 = 3'h1 == state;
  assign T58 = {1'h0, T59};
  assign T59 = release_count - 1'h1;
  assign T60 = T56 & T61;
  assign T61 = T49 ^ 1'h1;
  assign T62 = pending_outer_write ? 3'h3 : T63;
  assign T63 = T26 ? 3'h2 : 3'h4;
  assign T64 = T60 & T65;
  assign T65 = release_count == 1'h1;
  assign T66 = T67 ? 3'h5 : 3'h0;
  assign T67 = grant_type != 4'h0;
  assign grant_type = T86 ? T80 : T68;
  assign T68 = T79 ? 4'h2 : T69;
  assign T69 = T78 ? 4'h3 : T70;
  assign T70 = T77 ? 4'h4 : T71;
  assign T71 = T76 ? 4'h6 : T72;
  assign T72 = T75 ? 4'h7 : T73;
  assign T73 = T74 ? 4'h8 : 4'h3;
  assign T74 = xact_a_type == 3'h6;
  assign T75 = xact_a_type == 3'h5;
  assign T76 = xact_a_type == 3'h4;
  assign T77 = xact_a_type == 3'h3;
  assign T78 = xact_a_type == 3'h2;
  assign T79 = xact_a_type == 3'h1;
  assign T80 = T81 ? 4'h1 : 4'h2;
  assign T81 = 1'h0 < init_sharer_cnt;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = reset ? 2'h0 : T84;
  assign T84 = T22 ? 2'h2 : T85;
  assign T85 = {1'h0, init_sharer_cnt};
  assign T86 = xact_a_type == 3'h0;
  assign T87 = T88 & io_outer_acquire_ready;
  assign T88 = 3'h2 == state;
  assign T89 = T26 ? 3'h2 : 3'h4;
  assign T90 = T91 & io_outer_acquire_ready;
  assign T91 = 3'h3 == state;
  assign T92 = T93 ? 3'h5 : 3'h0;
  assign T93 = grant_type != 4'h0;
  assign T94 = T95 & io_inner_grant_ready;
  assign T95 = 3'h4 == state;
  assign T96 = T99 & T97;
  assign T97 = io_inner_finish_valid & T98;
  assign T98 = io_inner_finish_bits_payload_master_xact_id == 3'h7;
  assign T99 = 3'h5 == state;
  assign T100 = xact_addr == io_inner_release_bits_payload_addr;
  assign T101 = T22 ? io_inner_acquire_bits_payload_addr : xact_addr;
  assign io_has_acquire_conflict = T102;
  assign T102 = T104 & T103;
  assign T103 = state != 3'h0;
  assign T104 = xact_addr == io_inner_acquire_bits_payload_addr;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = T105;
  assign T105 = T91 ? outer_write_acq_atomic_opcode : T106;
  assign T106 = T88 ? outer_read_atomic_opcode : T107;
  assign T107 = T48 ? outer_write_rel_atomic_opcode : outer_read_atomic_opcode;
  assign outer_read_atomic_opcode = 4'h0;
  assign outer_write_rel_atomic_opcode = 4'h0;
  assign outer_write_acq_atomic_opcode = 4'h0;
  assign io_outer_acquire_bits_payload_subword_addr = T108;
  assign T108 = T91 ? outer_write_acq_subword_addr : T109;
  assign T109 = T88 ? outer_read_subword_addr : T110;
  assign T110 = T48 ? outer_write_rel_subword_addr : outer_read_subword_addr;
  assign outer_read_subword_addr = 3'h0;
  assign outer_write_rel_subword_addr = 3'h0;
  assign outer_write_acq_subword_addr = 3'h0;
  assign io_outer_acquire_bits_payload_write_mask = T111;
  assign T111 = T91 ? outer_write_acq_write_mask : T112;
  assign T112 = T88 ? outer_read_write_mask : T113;
  assign T113 = T48 ? outer_write_rel_write_mask : outer_read_write_mask;
  assign outer_read_write_mask = 6'h0;
  assign outer_write_rel_write_mask = 6'h0;
  assign outer_write_acq_write_mask = 6'h0;
  assign io_outer_acquire_bits_payload_a_type = T114;
  assign T114 = T91 ? outer_write_acq_a_type : T115;
  assign T115 = T88 ? outer_read_a_type : T116;
  assign T116 = T48 ? outer_write_rel_a_type : outer_read_a_type;
  assign outer_read_a_type = 3'h2;
  assign outer_write_rel_a_type = 3'h3;
  assign outer_write_acq_a_type = 3'h3;
  assign io_outer_acquire_bits_payload_data = T117;
  assign T117 = T91 ? outer_write_acq_data : T118;
  assign T118 = T88 ? outer_read_data : T119;
  assign T119 = T48 ? outer_write_rel_data : outer_read_data;
  assign outer_read_data = 512'h0;
  assign outer_write_rel_data = io_inner_release_bits_payload_data;
  assign outer_write_acq_data = xact_data;
  assign T120 = T22 ? io_inner_acquire_bits_payload_data : xact_data;
  assign io_outer_acquire_bits_payload_client_xact_id = T121;
  assign T121 = T91 ? outer_write_acq_client_xact_id : T122;
  assign T122 = T88 ? outer_read_client_xact_id : T123;
  assign T123 = T48 ? outer_write_rel_client_xact_id : outer_read_client_xact_id;
  assign outer_read_client_xact_id = 2'h3;
  assign outer_write_rel_client_xact_id = 2'h3;
  assign outer_write_acq_client_xact_id = 2'h3;
  assign io_outer_acquire_bits_payload_addr = T124;
  assign T124 = T91 ? outer_write_acq_addr : T125;
  assign T125 = T88 ? outer_read_addr : T126;
  assign T126 = T48 ? outer_write_rel_addr : outer_read_addr;
  assign outer_read_addr = xact_addr;
  assign outer_write_rel_addr = xact_addr;
  assign outer_write_acq_addr = xact_addr;
  assign io_outer_acquire_bits_header_src = 2'h0;
  assign io_outer_acquire_valid = T127;
  assign T127 = T91 ? 1'h1 : T128;
  assign T128 = T88 ? 1'h1 : T48;
  assign io_inner_release_ready = T129;
  assign T129 = T60 ? 1'h1 : T47;
  assign io_inner_probe_bits_payload_p_type = T130;
  assign T130 = T131;
  assign T131 = T144 ? 2'h1 : T132;
  assign T132 = T143 ? 2'h0 : T133;
  assign T133 = T142 ? 2'h2 : T134;
  assign T134 = T141 ? 2'h0 : T135;
  assign T135 = T140 ? 2'h2 : T136;
  assign T136 = T139 ? 2'h0 : T137;
  assign T137 = T138 ? 2'h0 : 2'h2;
  assign T138 = xact_a_type == 3'h6;
  assign T139 = xact_a_type == 3'h5;
  assign T140 = xact_a_type == 3'h4;
  assign T141 = xact_a_type == 3'h3;
  assign T142 = xact_a_type == 3'h2;
  assign T143 = xact_a_type == 3'h1;
  assign T144 = xact_a_type == 3'h0;
  assign io_inner_probe_bits_payload_master_xact_id = T145;
  assign T145 = 3'h7;
  assign io_inner_probe_bits_payload_addr = T146;
  assign T146 = xact_addr;
  assign io_inner_probe_bits_header_dst = T147;
  assign T147 = {1'h0, T148};
  assign T148 = T149 == 1'h0;
  assign T149 = probe_flags[1'h0:1'h0];
  assign T150 = reset ? 2'h0 : T151;
  assign T151 = T156 ? T153 : T152;
  assign T152 = T22 ? probe_initial_flags : probe_flags;
  assign T153 = probe_flags & T154;
  assign T154 = ~ T155;
  assign T155 = 1'h1 << T148;
  assign T156 = T57 & io_inner_probe_ready;
  assign io_inner_probe_bits_header_src = 2'h0;
  assign io_inner_probe_valid = T157;
  assign T157 = T57 ? T158 : 1'h0;
  assign T158 = probe_flags != 2'h0;
  assign io_inner_grant_bits_payload_g_type = T159;
  assign T159 = grant_type;
  assign io_inner_grant_bits_payload_master_xact_id = T160;
  assign T160 = 3'h7;
  assign io_inner_grant_bits_payload_client_xact_id = T161;
  assign T161 = xact_client_xact_id;
  assign T162 = T22 ? io_inner_acquire_bits_payload_client_xact_id : xact_client_xact_id;
  assign io_inner_grant_bits_payload_data = T163;
  assign T163 = io_outer_grant_bits_payload_data;
  assign io_inner_grant_bits_header_dst = T164;
  assign T164 = {1'h0, init_client_id};
  assign T165 = T166[1'h0:1'h0];
  assign T166 = reset ? 2'h0 : T167;
  assign T167 = T22 ? io_inner_acquire_bits_header_src : T168;
  assign T168 = {1'h0, init_client_id};
  assign io_inner_grant_bits_header_src = 2'h0;
  assign io_inner_grant_valid = T169;
  assign T169 = T170 ? 1'h1 : T95;
  assign T170 = T99 & T171;
  assign T171 = io_outer_grant_valid & T172;
  assign T172 = T173 == 3'h7;
  assign T173 = {1'h0, io_outer_grant_bits_payload_client_xact_id};
  assign io_inner_acquire_ready = T23;

  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else if(T96) begin
      state <= 3'h0;
    end else if(T94) begin
      state <= T92;
    end else if(T90) begin
      state <= T89;
    end else if(T87) begin
      state <= T66;
    end else if(T64) begin
      state <= T62;
    end else if(T32) begin
      state <= T24;
    end else if(T22) begin
      state <= T10;
    end
    if(T22) begin
      xact_a_type <= io_inner_acquire_bits_payload_a_type;
    end
    release_count <= T34;
    init_sharer_cnt <= T82;
    if(T22) begin
      xact_addr <= io_inner_acquire_bits_payload_addr;
    end
    if(T22) begin
      xact_data <= io_inner_acquire_bits_payload_data;
    end
    if(reset) begin
      probe_flags <= 2'h0;
    end else if(T156) begin
      probe_flags <= T153;
    end else if(T22) begin
      probe_flags <= probe_initial_flags;
    end
    if(T22) begin
      xact_client_xact_id <= io_inner_acquire_bits_payload_client_xact_id;
    end
    init_client_id <= T165;
  end
endmodule

module Arbiter_11(
    output io_in_7_ready,
    input  io_in_7_valid,
    input  io_in_7_bits,
    output io_in_6_ready,
    input  io_in_6_valid,
    input  io_in_6_bits,
    output io_in_5_ready,
    input  io_in_5_valid,
    input  io_in_5_bits,
    output io_in_4_ready,
    input  io_in_4_valid,
    input  io_in_4_bits,
    output io_in_3_ready,
    input  io_in_3_valid,
    input  io_in_3_bits,
    output io_in_2_ready,
    input  io_in_2_valid,
    input  io_in_2_bits,
    output io_in_1_ready,
    input  io_in_1_valid,
    input  io_in_1_bits,
    output io_in_0_ready,
    input  io_in_0_valid,
    input  io_in_0_bits,
    input  io_out_ready,
    output io_out_valid,
    output io_out_bits,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits : io_in_0_bits;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits : io_in_2_bits;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits : io_in_4_bits;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits : io_in_6_bits;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_valid = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_valid : io_in_0_valid;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_valid : io_in_2_valid;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_valid : io_in_4_valid;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_valid : io_in_6_valid;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T37;
  assign T37 = T38 & io_out_ready;
  assign T38 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T39;
  assign T39 = T40 & io_out_ready;
  assign T40 = T41 ^ 1'h1;
  assign T41 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T42;
  assign T42 = T43 & io_out_ready;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T45 | io_in_2_valid;
  assign T45 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T46;
  assign T46 = T47 & io_out_ready;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T49 | io_in_3_valid;
  assign T49 = T50 | io_in_2_valid;
  assign T50 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T51;
  assign T51 = T52 & io_out_ready;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T54 | io_in_4_valid;
  assign T54 = T55 | io_in_3_valid;
  assign T55 = T56 | io_in_2_valid;
  assign T56 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T57;
  assign T57 = T58 & io_out_ready;
  assign T58 = T59 ^ 1'h1;
  assign T59 = T60 | io_in_5_valid;
  assign T60 = T61 | io_in_4_valid;
  assign T61 = T62 | io_in_3_valid;
  assign T62 = T63 | io_in_2_valid;
  assign T63 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T64;
  assign T64 = T65 & io_out_ready;
  assign T65 = T66 ^ 1'h1;
  assign T66 = T67 | io_in_6_valid;
  assign T67 = T68 | io_in_5_valid;
  assign T68 = T69 | io_in_4_valid;
  assign T69 = T70 | io_in_3_valid;
  assign T70 = T71 | io_in_2_valid;
  assign T71 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_12(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [1:0] io_in_7_bits_payload_p_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [1:0] io_in_6_bits_payload_p_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [1:0] io_in_5_bits_payload_p_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [1:0] io_in_4_bits_payload_p_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [1:0] io_in_3_bits_payload_p_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [1:0] io_in_2_bits_payload_p_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [1:0] io_in_1_bits_payload_p_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [1:0] io_in_0_bits_payload_p_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[1:0] io_out_bits_payload_p_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire T18;
  wire[1:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[25:0] T37;
  wire[25:0] T38;
  wire[25:0] T39;
  wire T40;
  wire[25:0] T41;
  wire T42;
  wire T43;
  wire[25:0] T44;
  wire[25:0] T45;
  wire T46;
  wire[25:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire[1:0] T53;
  wire T54;
  wire[1:0] T55;
  wire T56;
  wire T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire T60;
  wire[1:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_p_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_p_type : io_in_2_bits_payload_p_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_p_type : io_in_4_bits_payload_p_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_p_type : io_in_6_bits_payload_p_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_addr = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_valid = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_valid : io_in_0_valid;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_valid : io_in_2_valid;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_valid : io_in_4_valid;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_valid : io_in_6_valid;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T93;
  assign T93 = T94 & io_out_ready;
  assign T94 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T95;
  assign T95 = T96 & io_out_ready;
  assign T96 = T97 ^ 1'h1;
  assign T97 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T98;
  assign T98 = T99 & io_out_ready;
  assign T99 = T100 ^ 1'h1;
  assign T100 = T101 | io_in_2_valid;
  assign T101 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T102;
  assign T102 = T103 & io_out_ready;
  assign T103 = T104 ^ 1'h1;
  assign T104 = T105 | io_in_3_valid;
  assign T105 = T106 | io_in_2_valid;
  assign T106 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = T109 ^ 1'h1;
  assign T109 = T110 | io_in_4_valid;
  assign T110 = T111 | io_in_3_valid;
  assign T111 = T112 | io_in_2_valid;
  assign T112 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T113;
  assign T113 = T114 & io_out_ready;
  assign T114 = T115 ^ 1'h1;
  assign T115 = T116 | io_in_5_valid;
  assign T116 = T117 | io_in_4_valid;
  assign T117 = T118 | io_in_3_valid;
  assign T118 = T119 | io_in_2_valid;
  assign T119 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T120;
  assign T120 = T121 & io_out_ready;
  assign T121 = T122 ^ 1'h1;
  assign T122 = T123 | io_in_6_valid;
  assign T123 = T124 | io_in_5_valid;
  assign T124 = T125 | io_in_4_valid;
  assign T125 = T126 | io_in_3_valid;
  assign T126 = T127 | io_in_2_valid;
  assign T127 = io_in_0_valid | io_in_1_valid;
endmodule

module Arbiter_13(
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [511:0] io_in_7_bits_payload_data,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    input [3:0] io_in_7_bits_payload_g_type,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [511:0] io_in_6_bits_payload_data,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    input [3:0] io_in_6_bits_payload_g_type,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [511:0] io_in_5_bits_payload_data,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    input [3:0] io_in_5_bits_payload_g_type,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [511:0] io_in_4_bits_payload_data,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    input [3:0] io_in_4_bits_payload_g_type,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [511:0] io_in_3_bits_payload_data,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    input [3:0] io_in_3_bits_payload_g_type,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [511:0] io_in_2_bits_payload_data,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    input [3:0] io_in_2_bits_payload_g_type,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [511:0] io_in_1_bits_payload_data,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    input [3:0] io_in_1_bits_payload_g_type,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [511:0] io_in_0_bits_payload_data,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input [3:0] io_in_0_bits_payload_g_type,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[511:0] io_out_bits_payload_data,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[3:0] io_out_bits_payload_g_type,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[3:0] T10;
  wire T11;
  wire[2:0] T12;
  wire[3:0] T13;
  wire T14;
  wire T15;
  wire[3:0] T16;
  wire[3:0] T17;
  wire T18;
  wire[3:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire[2:0] T23;
  wire[2:0] T24;
  wire[2:0] T25;
  wire T26;
  wire[2:0] T27;
  wire T28;
  wire T29;
  wire[2:0] T30;
  wire[2:0] T31;
  wire T32;
  wire[2:0] T33;
  wire T34;
  wire T35;
  wire T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[1:0] T44;
  wire[1:0] T45;
  wire T46;
  wire[1:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire[511:0] T51;
  wire[511:0] T52;
  wire[511:0] T53;
  wire T54;
  wire[511:0] T55;
  wire T56;
  wire T57;
  wire[511:0] T58;
  wire[511:0] T59;
  wire T60;
  wire[511:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire[1:0] T69;
  wire T70;
  wire T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire T82;
  wire[1:0] T83;
  wire T84;
  wire T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire T88;
  wire[1:0] T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;


  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = io_in_0_valid ? 3'h0 : T2;
  assign T2 = io_in_1_valid ? 3'h1 : T3;
  assign T3 = io_in_2_valid ? 3'h2 : T4;
  assign T4 = io_in_3_valid ? 3'h3 : T5;
  assign T5 = io_in_4_valid ? 3'h4 : T6;
  assign T6 = io_in_5_valid ? 3'h5 : T7;
  assign T7 = io_in_6_valid ? 3'h6 : 3'h7;
  assign io_out_bits_payload_g_type = T8;
  assign T8 = T22 ? T16 : T9;
  assign T9 = T15 ? T13 : T10;
  assign T10 = T11 ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign T11 = T12[1'h0:1'h0];
  assign T12 = T0;
  assign T13 = T14 ? io_in_3_bits_payload_g_type : io_in_2_bits_payload_g_type;
  assign T14 = T12[1'h0:1'h0];
  assign T15 = T12[1'h1:1'h1];
  assign T16 = T21 ? T19 : T17;
  assign T17 = T18 ? io_in_5_bits_payload_g_type : io_in_4_bits_payload_g_type;
  assign T18 = T12[1'h0:1'h0];
  assign T19 = T20 ? io_in_7_bits_payload_g_type : io_in_6_bits_payload_g_type;
  assign T20 = T12[1'h0:1'h0];
  assign T21 = T12[1'h1:1'h1];
  assign T22 = T12[2'h2:2'h2];
  assign io_out_bits_payload_master_xact_id = T23;
  assign T23 = T36 ? T30 : T24;
  assign T24 = T29 ? T27 : T25;
  assign T25 = T26 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T26 = T12[1'h0:1'h0];
  assign T27 = T28 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T28 = T12[1'h0:1'h0];
  assign T29 = T12[1'h1:1'h1];
  assign T30 = T35 ? T33 : T31;
  assign T31 = T32 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T32 = T12[1'h0:1'h0];
  assign T33 = T34 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T34 = T12[1'h0:1'h0];
  assign T35 = T12[1'h1:1'h1];
  assign T36 = T12[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T37;
  assign T37 = T50 ? T44 : T38;
  assign T38 = T43 ? T41 : T39;
  assign T39 = T40 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T40 = T12[1'h0:1'h0];
  assign T41 = T42 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T42 = T12[1'h0:1'h0];
  assign T43 = T12[1'h1:1'h1];
  assign T44 = T49 ? T47 : T45;
  assign T45 = T46 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T46 = T12[1'h0:1'h0];
  assign T47 = T48 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T48 = T12[1'h0:1'h0];
  assign T49 = T12[1'h1:1'h1];
  assign T50 = T12[2'h2:2'h2];
  assign io_out_bits_payload_data = T51;
  assign T51 = T64 ? T58 : T52;
  assign T52 = T57 ? T55 : T53;
  assign T53 = T54 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T54 = T12[1'h0:1'h0];
  assign T55 = T56 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T56 = T12[1'h0:1'h0];
  assign T57 = T12[1'h1:1'h1];
  assign T58 = T63 ? T61 : T59;
  assign T59 = T60 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T60 = T12[1'h0:1'h0];
  assign T61 = T62 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T62 = T12[1'h0:1'h0];
  assign T63 = T12[1'h1:1'h1];
  assign T64 = T12[2'h2:2'h2];
  assign io_out_bits_header_dst = T65;
  assign T65 = T78 ? T72 : T66;
  assign T66 = T71 ? T69 : T67;
  assign T67 = T68 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T68 = T12[1'h0:1'h0];
  assign T69 = T70 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T70 = T12[1'h0:1'h0];
  assign T71 = T12[1'h1:1'h1];
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T74 = T12[1'h0:1'h0];
  assign T75 = T76 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T76 = T12[1'h0:1'h0];
  assign T77 = T12[1'h1:1'h1];
  assign T78 = T12[2'h2:2'h2];
  assign io_out_bits_header_src = T79;
  assign T79 = T92 ? T86 : T80;
  assign T80 = T85 ? T83 : T81;
  assign T81 = T82 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T82 = T12[1'h0:1'h0];
  assign T83 = T84 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T84 = T12[1'h0:1'h0];
  assign T85 = T12[1'h1:1'h1];
  assign T86 = T91 ? T89 : T87;
  assign T87 = T88 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T88 = T12[1'h0:1'h0];
  assign T89 = T90 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T90 = T12[1'h0:1'h0];
  assign T91 = T12[1'h1:1'h1];
  assign T92 = T12[2'h2:2'h2];
  assign io_out_valid = T93;
  assign T93 = T106 ? T100 : T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96 ? io_in_1_valid : io_in_0_valid;
  assign T96 = T12[1'h0:1'h0];
  assign T97 = T98 ? io_in_3_valid : io_in_2_valid;
  assign T98 = T12[1'h0:1'h0];
  assign T99 = T12[1'h1:1'h1];
  assign T100 = T105 ? T103 : T101;
  assign T101 = T102 ? io_in_5_valid : io_in_4_valid;
  assign T102 = T12[1'h0:1'h0];
  assign T103 = T104 ? io_in_7_valid : io_in_6_valid;
  assign T104 = T12[1'h0:1'h0];
  assign T105 = T12[1'h1:1'h1];
  assign T106 = T12[2'h2:2'h2];
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T107;
  assign T107 = T108 & io_out_ready;
  assign T108 = io_in_0_valid ^ 1'h1;
  assign io_in_2_ready = T109;
  assign T109 = T110 & io_out_ready;
  assign T110 = T111 ^ 1'h1;
  assign T111 = io_in_0_valid | io_in_1_valid;
  assign io_in_3_ready = T112;
  assign T112 = T113 & io_out_ready;
  assign T113 = T114 ^ 1'h1;
  assign T114 = T115 | io_in_2_valid;
  assign T115 = io_in_0_valid | io_in_1_valid;
  assign io_in_4_ready = T116;
  assign T116 = T117 & io_out_ready;
  assign T117 = T118 ^ 1'h1;
  assign T118 = T119 | io_in_3_valid;
  assign T119 = T120 | io_in_2_valid;
  assign T120 = io_in_0_valid | io_in_1_valid;
  assign io_in_5_ready = T121;
  assign T121 = T122 & io_out_ready;
  assign T122 = T123 ^ 1'h1;
  assign T123 = T124 | io_in_4_valid;
  assign T124 = T125 | io_in_3_valid;
  assign T125 = T126 | io_in_2_valid;
  assign T126 = io_in_0_valid | io_in_1_valid;
  assign io_in_6_ready = T127;
  assign T127 = T128 & io_out_ready;
  assign T128 = T129 ^ 1'h1;
  assign T129 = T130 | io_in_5_valid;
  assign T130 = T131 | io_in_4_valid;
  assign T131 = T132 | io_in_3_valid;
  assign T132 = T133 | io_in_2_valid;
  assign T133 = io_in_0_valid | io_in_1_valid;
  assign io_in_7_ready = T134;
  assign T134 = T135 & io_out_ready;
  assign T135 = T136 ^ 1'h1;
  assign T136 = T137 | io_in_6_valid;
  assign T137 = T138 | io_in_5_valid;
  assign T138 = T139 | io_in_4_valid;
  assign T139 = T140 | io_in_3_valid;
  assign T140 = T141 | io_in_2_valid;
  assign T141 = io_in_0_valid | io_in_1_valid;
endmodule

module RRArbiter_3(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [25:0] io_in_7_bits_payload_addr,
    input [1:0] io_in_7_bits_payload_client_xact_id,
    input [511:0] io_in_7_bits_payload_data,
    input [2:0] io_in_7_bits_payload_a_type,
    input [5:0] io_in_7_bits_payload_write_mask,
    input [2:0] io_in_7_bits_payload_subword_addr,
    input [3:0] io_in_7_bits_payload_atomic_opcode,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [25:0] io_in_6_bits_payload_addr,
    input [1:0] io_in_6_bits_payload_client_xact_id,
    input [511:0] io_in_6_bits_payload_data,
    input [2:0] io_in_6_bits_payload_a_type,
    input [5:0] io_in_6_bits_payload_write_mask,
    input [2:0] io_in_6_bits_payload_subword_addr,
    input [3:0] io_in_6_bits_payload_atomic_opcode,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [25:0] io_in_5_bits_payload_addr,
    input [1:0] io_in_5_bits_payload_client_xact_id,
    input [511:0] io_in_5_bits_payload_data,
    input [2:0] io_in_5_bits_payload_a_type,
    input [5:0] io_in_5_bits_payload_write_mask,
    input [2:0] io_in_5_bits_payload_subword_addr,
    input [3:0] io_in_5_bits_payload_atomic_opcode,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [25:0] io_in_4_bits_payload_addr,
    input [1:0] io_in_4_bits_payload_client_xact_id,
    input [511:0] io_in_4_bits_payload_data,
    input [2:0] io_in_4_bits_payload_a_type,
    input [5:0] io_in_4_bits_payload_write_mask,
    input [2:0] io_in_4_bits_payload_subword_addr,
    input [3:0] io_in_4_bits_payload_atomic_opcode,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [25:0] io_in_3_bits_payload_addr,
    input [1:0] io_in_3_bits_payload_client_xact_id,
    input [511:0] io_in_3_bits_payload_data,
    input [2:0] io_in_3_bits_payload_a_type,
    input [5:0] io_in_3_bits_payload_write_mask,
    input [2:0] io_in_3_bits_payload_subword_addr,
    input [3:0] io_in_3_bits_payload_atomic_opcode,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [25:0] io_in_2_bits_payload_addr,
    input [1:0] io_in_2_bits_payload_client_xact_id,
    input [511:0] io_in_2_bits_payload_data,
    input [2:0] io_in_2_bits_payload_a_type,
    input [5:0] io_in_2_bits_payload_write_mask,
    input [2:0] io_in_2_bits_payload_subword_addr,
    input [3:0] io_in_2_bits_payload_atomic_opcode,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [25:0] io_in_1_bits_payload_addr,
    input [1:0] io_in_1_bits_payload_client_xact_id,
    input [511:0] io_in_1_bits_payload_data,
    input [2:0] io_in_1_bits_payload_a_type,
    input [5:0] io_in_1_bits_payload_write_mask,
    input [2:0] io_in_1_bits_payload_subword_addr,
    input [3:0] io_in_1_bits_payload_atomic_opcode,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [25:0] io_in_0_bits_payload_addr,
    input [1:0] io_in_0_bits_payload_client_xact_id,
    input [511:0] io_in_0_bits_payload_data,
    input [2:0] io_in_0_bits_payload_a_type,
    input [5:0] io_in_0_bits_payload_write_mask,
    input [2:0] io_in_0_bits_payload_subword_addr,
    input [3:0] io_in_0_bits_payload_atomic_opcode,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[25:0] io_out_bits_payload_addr,
    output[1:0] io_out_bits_payload_client_xact_id,
    output[511:0] io_out_bits_payload_data,
    output[2:0] io_out_bits_payload_a_type,
    output[5:0] io_out_bits_payload_write_mask,
    output[2:0] io_out_bits_payload_subword_addr,
    output[3:0] io_out_bits_payload_atomic_opcode,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[3:0] T33;
  wire[3:0] T34;
  wire[3:0] T35;
  wire T36;
  wire[2:0] T37;
  wire[3:0] T38;
  wire T39;
  wire T40;
  wire[3:0] T41;
  wire[3:0] T42;
  wire T43;
  wire[3:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[2:0] T48;
  wire[2:0] T49;
  wire[2:0] T50;
  wire T51;
  wire[2:0] T52;
  wire T53;
  wire T54;
  wire[2:0] T55;
  wire[2:0] T56;
  wire T57;
  wire[2:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[5:0] T62;
  wire[5:0] T63;
  wire[5:0] T64;
  wire T65;
  wire[5:0] T66;
  wire T67;
  wire T68;
  wire[5:0] T69;
  wire[5:0] T70;
  wire T71;
  wire[5:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire[2:0] T76;
  wire[2:0] T77;
  wire[2:0] T78;
  wire T79;
  wire[2:0] T80;
  wire T81;
  wire T82;
  wire[2:0] T83;
  wire[2:0] T84;
  wire T85;
  wire[2:0] T86;
  wire T87;
  wire T88;
  wire T89;
  wire[511:0] T90;
  wire[511:0] T91;
  wire[511:0] T92;
  wire T93;
  wire[511:0] T94;
  wire T95;
  wire T96;
  wire[511:0] T97;
  wire[511:0] T98;
  wire T99;
  wire[511:0] T100;
  wire T101;
  wire T102;
  wire T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire[1:0] T106;
  wire T107;
  wire[1:0] T108;
  wire T109;
  wire T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire T113;
  wire[1:0] T114;
  wire T115;
  wire T116;
  wire T117;
  wire[25:0] T118;
  wire[25:0] T119;
  wire[25:0] T120;
  wire T121;
  wire[25:0] T122;
  wire T123;
  wire T124;
  wire[25:0] T125;
  wire[25:0] T126;
  wire T127;
  wire[25:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[1:0] T132;
  wire[1:0] T133;
  wire[1:0] T134;
  wire T135;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire[1:0] T139;
  wire[1:0] T140;
  wire T141;
  wire[1:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire[1:0] T146;
  wire[1:0] T147;
  wire[1:0] T148;
  wire T149;
  wire[1:0] T150;
  wire T151;
  wire T152;
  wire[1:0] T153;
  wire[1:0] T154;
  wire T155;
  wire[1:0] T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T31 ? 3'h1 : T2;
  assign T2 = T29 ? 3'h2 : T3;
  assign T3 = T27 ? 3'h3 : T4;
  assign T4 = T25 ? 3'h4 : T5;
  assign T5 = T23 ? 3'h5 : T6;
  assign T6 = T21 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T18 = reset ? 3'h0 : T19;
  assign T19 = T20 ? T0 : R17;
  assign T20 = io_out_ready & io_out_valid;
  assign T21 = io_in_6_valid & T22;
  assign T22 = R17 < 3'h6;
  assign T23 = io_in_5_valid & T24;
  assign T24 = R17 < 3'h5;
  assign T25 = io_in_4_valid & T26;
  assign T26 = R17 < 3'h4;
  assign T27 = io_in_3_valid & T28;
  assign T28 = R17 < 3'h3;
  assign T29 = io_in_2_valid & T30;
  assign T30 = R17 < 3'h2;
  assign T31 = io_in_1_valid & T32;
  assign T32 = R17 < 3'h1;
  assign io_out_bits_payload_atomic_opcode = T33;
  assign T33 = T47 ? T41 : T34;
  assign T34 = T40 ? T38 : T35;
  assign T35 = T36 ? io_in_1_bits_payload_atomic_opcode : io_in_0_bits_payload_atomic_opcode;
  assign T36 = T37[1'h0:1'h0];
  assign T37 = T0;
  assign T38 = T39 ? io_in_3_bits_payload_atomic_opcode : io_in_2_bits_payload_atomic_opcode;
  assign T39 = T37[1'h0:1'h0];
  assign T40 = T37[1'h1:1'h1];
  assign T41 = T46 ? T44 : T42;
  assign T42 = T43 ? io_in_5_bits_payload_atomic_opcode : io_in_4_bits_payload_atomic_opcode;
  assign T43 = T37[1'h0:1'h0];
  assign T44 = T45 ? io_in_7_bits_payload_atomic_opcode : io_in_6_bits_payload_atomic_opcode;
  assign T45 = T37[1'h0:1'h0];
  assign T46 = T37[1'h1:1'h1];
  assign T47 = T37[2'h2:2'h2];
  assign io_out_bits_payload_subword_addr = T48;
  assign T48 = T61 ? T55 : T49;
  assign T49 = T54 ? T52 : T50;
  assign T50 = T51 ? io_in_1_bits_payload_subword_addr : io_in_0_bits_payload_subword_addr;
  assign T51 = T37[1'h0:1'h0];
  assign T52 = T53 ? io_in_3_bits_payload_subword_addr : io_in_2_bits_payload_subword_addr;
  assign T53 = T37[1'h0:1'h0];
  assign T54 = T37[1'h1:1'h1];
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_5_bits_payload_subword_addr : io_in_4_bits_payload_subword_addr;
  assign T57 = T37[1'h0:1'h0];
  assign T58 = T59 ? io_in_7_bits_payload_subword_addr : io_in_6_bits_payload_subword_addr;
  assign T59 = T37[1'h0:1'h0];
  assign T60 = T37[1'h1:1'h1];
  assign T61 = T37[2'h2:2'h2];
  assign io_out_bits_payload_write_mask = T62;
  assign T62 = T75 ? T69 : T63;
  assign T63 = T68 ? T66 : T64;
  assign T64 = T65 ? io_in_1_bits_payload_write_mask : io_in_0_bits_payload_write_mask;
  assign T65 = T37[1'h0:1'h0];
  assign T66 = T67 ? io_in_3_bits_payload_write_mask : io_in_2_bits_payload_write_mask;
  assign T67 = T37[1'h0:1'h0];
  assign T68 = T37[1'h1:1'h1];
  assign T69 = T74 ? T72 : T70;
  assign T70 = T71 ? io_in_5_bits_payload_write_mask : io_in_4_bits_payload_write_mask;
  assign T71 = T37[1'h0:1'h0];
  assign T72 = T73 ? io_in_7_bits_payload_write_mask : io_in_6_bits_payload_write_mask;
  assign T73 = T37[1'h0:1'h0];
  assign T74 = T37[1'h1:1'h1];
  assign T75 = T37[2'h2:2'h2];
  assign io_out_bits_payload_a_type = T76;
  assign T76 = T89 ? T83 : T77;
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign T79 = T37[1'h0:1'h0];
  assign T80 = T81 ? io_in_3_bits_payload_a_type : io_in_2_bits_payload_a_type;
  assign T81 = T37[1'h0:1'h0];
  assign T82 = T37[1'h1:1'h1];
  assign T83 = T88 ? T86 : T84;
  assign T84 = T85 ? io_in_5_bits_payload_a_type : io_in_4_bits_payload_a_type;
  assign T85 = T37[1'h0:1'h0];
  assign T86 = T87 ? io_in_7_bits_payload_a_type : io_in_6_bits_payload_a_type;
  assign T87 = T37[1'h0:1'h0];
  assign T88 = T37[1'h1:1'h1];
  assign T89 = T37[2'h2:2'h2];
  assign io_out_bits_payload_data = T90;
  assign T90 = T103 ? T97 : T91;
  assign T91 = T96 ? T94 : T92;
  assign T92 = T93 ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign T93 = T37[1'h0:1'h0];
  assign T94 = T95 ? io_in_3_bits_payload_data : io_in_2_bits_payload_data;
  assign T95 = T37[1'h0:1'h0];
  assign T96 = T37[1'h1:1'h1];
  assign T97 = T102 ? T100 : T98;
  assign T98 = T99 ? io_in_5_bits_payload_data : io_in_4_bits_payload_data;
  assign T99 = T37[1'h0:1'h0];
  assign T100 = T101 ? io_in_7_bits_payload_data : io_in_6_bits_payload_data;
  assign T101 = T37[1'h0:1'h0];
  assign T102 = T37[1'h1:1'h1];
  assign T103 = T37[2'h2:2'h2];
  assign io_out_bits_payload_client_xact_id = T104;
  assign T104 = T117 ? T111 : T105;
  assign T105 = T110 ? T108 : T106;
  assign T106 = T107 ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign T107 = T37[1'h0:1'h0];
  assign T108 = T109 ? io_in_3_bits_payload_client_xact_id : io_in_2_bits_payload_client_xact_id;
  assign T109 = T37[1'h0:1'h0];
  assign T110 = T37[1'h1:1'h1];
  assign T111 = T116 ? T114 : T112;
  assign T112 = T113 ? io_in_5_bits_payload_client_xact_id : io_in_4_bits_payload_client_xact_id;
  assign T113 = T37[1'h0:1'h0];
  assign T114 = T115 ? io_in_7_bits_payload_client_xact_id : io_in_6_bits_payload_client_xact_id;
  assign T115 = T37[1'h0:1'h0];
  assign T116 = T37[1'h1:1'h1];
  assign T117 = T37[2'h2:2'h2];
  assign io_out_bits_payload_addr = T118;
  assign T118 = T131 ? T125 : T119;
  assign T119 = T124 ? T122 : T120;
  assign T120 = T121 ? io_in_1_bits_payload_addr : io_in_0_bits_payload_addr;
  assign T121 = T37[1'h0:1'h0];
  assign T122 = T123 ? io_in_3_bits_payload_addr : io_in_2_bits_payload_addr;
  assign T123 = T37[1'h0:1'h0];
  assign T124 = T37[1'h1:1'h1];
  assign T125 = T130 ? T128 : T126;
  assign T126 = T127 ? io_in_5_bits_payload_addr : io_in_4_bits_payload_addr;
  assign T127 = T37[1'h0:1'h0];
  assign T128 = T129 ? io_in_7_bits_payload_addr : io_in_6_bits_payload_addr;
  assign T129 = T37[1'h0:1'h0];
  assign T130 = T37[1'h1:1'h1];
  assign T131 = T37[2'h2:2'h2];
  assign io_out_bits_header_dst = T132;
  assign T132 = T145 ? T139 : T133;
  assign T133 = T138 ? T136 : T134;
  assign T134 = T135 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T135 = T37[1'h0:1'h0];
  assign T136 = T137 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T137 = T37[1'h0:1'h0];
  assign T138 = T37[1'h1:1'h1];
  assign T139 = T144 ? T142 : T140;
  assign T140 = T141 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T141 = T37[1'h0:1'h0];
  assign T142 = T143 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T143 = T37[1'h0:1'h0];
  assign T144 = T37[1'h1:1'h1];
  assign T145 = T37[2'h2:2'h2];
  assign io_out_bits_header_src = T146;
  assign T146 = T159 ? T153 : T147;
  assign T147 = T152 ? T150 : T148;
  assign T148 = T149 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T149 = T37[1'h0:1'h0];
  assign T150 = T151 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T151 = T37[1'h0:1'h0];
  assign T152 = T37[1'h1:1'h1];
  assign T153 = T158 ? T156 : T154;
  assign T154 = T155 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T155 = T37[1'h0:1'h0];
  assign T156 = T157 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T157 = T37[1'h0:1'h0];
  assign T158 = T37[1'h1:1'h1];
  assign T159 = T37[2'h2:2'h2];
  assign io_out_valid = T160;
  assign T160 = T173 ? T167 : T161;
  assign T161 = T166 ? T164 : T162;
  assign T162 = T163 ? io_in_1_valid : io_in_0_valid;
  assign T163 = T37[1'h0:1'h0];
  assign T164 = T165 ? io_in_3_valid : io_in_2_valid;
  assign T165 = T37[1'h0:1'h0];
  assign T166 = T37[1'h1:1'h1];
  assign T167 = T172 ? T170 : T168;
  assign T168 = T169 ? io_in_5_valid : io_in_4_valid;
  assign T169 = T37[1'h0:1'h0];
  assign T170 = T171 ? io_in_7_valid : io_in_6_valid;
  assign T171 = T37[1'h0:1'h0];
  assign T172 = T37[1'h1:1'h1];
  assign T173 = T37[2'h2:2'h2];
  assign io_in_0_ready = T174;
  assign T174 = T175 & io_out_ready;
  assign T175 = T200 | T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = T180 | T178;
  assign T178 = io_in_7_valid & T179;
  assign T179 = R17 < 3'h7;
  assign T180 = T183 | T181;
  assign T181 = io_in_6_valid & T182;
  assign T182 = R17 < 3'h6;
  assign T183 = T186 | T184;
  assign T184 = io_in_5_valid & T185;
  assign T185 = R17 < 3'h5;
  assign T186 = T189 | T187;
  assign T187 = io_in_4_valid & T188;
  assign T188 = R17 < 3'h4;
  assign T189 = T192 | T190;
  assign T190 = io_in_3_valid & T191;
  assign T191 = R17 < 3'h3;
  assign T192 = T195 | T193;
  assign T193 = io_in_2_valid & T194;
  assign T194 = R17 < 3'h2;
  assign T195 = T198 | T196;
  assign T196 = io_in_1_valid & T197;
  assign T197 = R17 < 3'h1;
  assign T198 = io_in_0_valid & T199;
  assign T199 = R17 < 3'h0;
  assign T200 = R17 < 3'h0;
  assign io_in_1_ready = T201;
  assign T201 = T202 & io_out_ready;
  assign T202 = T212 | T203;
  assign T203 = T204 ^ 1'h1;
  assign T204 = T205 | io_in_0_valid;
  assign T205 = T206 | T178;
  assign T206 = T207 | T181;
  assign T207 = T208 | T184;
  assign T208 = T209 | T187;
  assign T209 = T210 | T190;
  assign T210 = T211 | T193;
  assign T211 = T198 | T196;
  assign T212 = T214 & T213;
  assign T213 = R17 < 3'h1;
  assign T214 = T198 ^ 1'h1;
  assign io_in_2_ready = T215;
  assign T215 = T216 & io_out_ready;
  assign T216 = T227 | T217;
  assign T217 = T218 ^ 1'h1;
  assign T218 = T219 | io_in_1_valid;
  assign T219 = T220 | io_in_0_valid;
  assign T220 = T221 | T178;
  assign T221 = T222 | T181;
  assign T222 = T223 | T184;
  assign T223 = T224 | T187;
  assign T224 = T225 | T190;
  assign T225 = T226 | T193;
  assign T226 = T198 | T196;
  assign T227 = T229 & T228;
  assign T228 = R17 < 3'h2;
  assign T229 = T230 ^ 1'h1;
  assign T230 = T198 | T196;
  assign io_in_3_ready = T231;
  assign T231 = T232 & io_out_ready;
  assign T232 = T244 | T233;
  assign T233 = T234 ^ 1'h1;
  assign T234 = T235 | io_in_2_valid;
  assign T235 = T236 | io_in_1_valid;
  assign T236 = T237 | io_in_0_valid;
  assign T237 = T238 | T178;
  assign T238 = T239 | T181;
  assign T239 = T240 | T184;
  assign T240 = T241 | T187;
  assign T241 = T242 | T190;
  assign T242 = T243 | T193;
  assign T243 = T198 | T196;
  assign T244 = T246 & T245;
  assign T245 = R17 < 3'h3;
  assign T246 = T247 ^ 1'h1;
  assign T247 = T248 | T193;
  assign T248 = T198 | T196;
  assign io_in_4_ready = T249;
  assign T249 = T250 & io_out_ready;
  assign T250 = T263 | T251;
  assign T251 = T252 ^ 1'h1;
  assign T252 = T253 | io_in_3_valid;
  assign T253 = T254 | io_in_2_valid;
  assign T254 = T255 | io_in_1_valid;
  assign T255 = T256 | io_in_0_valid;
  assign T256 = T257 | T178;
  assign T257 = T258 | T181;
  assign T258 = T259 | T184;
  assign T259 = T260 | T187;
  assign T260 = T261 | T190;
  assign T261 = T262 | T193;
  assign T262 = T198 | T196;
  assign T263 = T265 & T264;
  assign T264 = R17 < 3'h4;
  assign T265 = T266 ^ 1'h1;
  assign T266 = T267 | T190;
  assign T267 = T268 | T193;
  assign T268 = T198 | T196;
  assign io_in_5_ready = T269;
  assign T269 = T270 & io_out_ready;
  assign T270 = T284 | T271;
  assign T271 = T272 ^ 1'h1;
  assign T272 = T273 | io_in_4_valid;
  assign T273 = T274 | io_in_3_valid;
  assign T274 = T275 | io_in_2_valid;
  assign T275 = T276 | io_in_1_valid;
  assign T276 = T277 | io_in_0_valid;
  assign T277 = T278 | T178;
  assign T278 = T279 | T181;
  assign T279 = T280 | T184;
  assign T280 = T281 | T187;
  assign T281 = T282 | T190;
  assign T282 = T283 | T193;
  assign T283 = T198 | T196;
  assign T284 = T286 & T285;
  assign T285 = R17 < 3'h5;
  assign T286 = T287 ^ 1'h1;
  assign T287 = T288 | T187;
  assign T288 = T289 | T190;
  assign T289 = T290 | T193;
  assign T290 = T198 | T196;
  assign io_in_6_ready = T291;
  assign T291 = T292 & io_out_ready;
  assign T292 = T307 | T293;
  assign T293 = T294 ^ 1'h1;
  assign T294 = T295 | io_in_5_valid;
  assign T295 = T296 | io_in_4_valid;
  assign T296 = T297 | io_in_3_valid;
  assign T297 = T298 | io_in_2_valid;
  assign T298 = T299 | io_in_1_valid;
  assign T299 = T300 | io_in_0_valid;
  assign T300 = T301 | T178;
  assign T301 = T302 | T181;
  assign T302 = T303 | T184;
  assign T303 = T304 | T187;
  assign T304 = T305 | T190;
  assign T305 = T306 | T193;
  assign T306 = T198 | T196;
  assign T307 = T309 & T308;
  assign T308 = R17 < 3'h6;
  assign T309 = T310 ^ 1'h1;
  assign T310 = T311 | T184;
  assign T311 = T312 | T187;
  assign T312 = T313 | T190;
  assign T313 = T314 | T193;
  assign T314 = T198 | T196;
  assign io_in_7_ready = T315;
  assign T315 = T316 & io_out_ready;
  assign T316 = T332 | T317;
  assign T317 = T318 ^ 1'h1;
  assign T318 = T319 | io_in_6_valid;
  assign T319 = T320 | io_in_5_valid;
  assign T320 = T321 | io_in_4_valid;
  assign T321 = T322 | io_in_3_valid;
  assign T322 = T323 | io_in_2_valid;
  assign T323 = T324 | io_in_1_valid;
  assign T324 = T325 | io_in_0_valid;
  assign T325 = T326 | T178;
  assign T326 = T327 | T181;
  assign T327 = T328 | T184;
  assign T328 = T329 | T187;
  assign T329 = T330 | T190;
  assign T330 = T331 | T193;
  assign T331 = T198 | T196;
  assign T332 = T334 & T333;
  assign T333 = R17 < 3'h7;
  assign T334 = T335 ^ 1'h1;
  assign T335 = T336 | T181;
  assign T336 = T337 | T184;
  assign T337 = T338 | T187;
  assign T338 = T339 | T190;
  assign T339 = T340 | T193;
  assign T340 = T198 | T196;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T20) begin
      R17 <= T0;
    end
  end
endmodule

module RRArbiter_4(input clk, input reset,
    output io_in_7_ready,
    input  io_in_7_valid,
    input [1:0] io_in_7_bits_header_src,
    input [1:0] io_in_7_bits_header_dst,
    input [2:0] io_in_7_bits_payload_master_xact_id,
    output io_in_6_ready,
    input  io_in_6_valid,
    input [1:0] io_in_6_bits_header_src,
    input [1:0] io_in_6_bits_header_dst,
    input [2:0] io_in_6_bits_payload_master_xact_id,
    output io_in_5_ready,
    input  io_in_5_valid,
    input [1:0] io_in_5_bits_header_src,
    input [1:0] io_in_5_bits_header_dst,
    input [2:0] io_in_5_bits_payload_master_xact_id,
    output io_in_4_ready,
    input  io_in_4_valid,
    input [1:0] io_in_4_bits_header_src,
    input [1:0] io_in_4_bits_header_dst,
    input [2:0] io_in_4_bits_payload_master_xact_id,
    output io_in_3_ready,
    input  io_in_3_valid,
    input [1:0] io_in_3_bits_header_src,
    input [1:0] io_in_3_bits_header_dst,
    input [2:0] io_in_3_bits_payload_master_xact_id,
    output io_in_2_ready,
    input  io_in_2_valid,
    input [1:0] io_in_2_bits_header_src,
    input [1:0] io_in_2_bits_header_dst,
    input [2:0] io_in_2_bits_payload_master_xact_id,
    output io_in_1_ready,
    input  io_in_1_valid,
    input [1:0] io_in_1_bits_header_src,
    input [1:0] io_in_1_bits_header_dst,
    input [2:0] io_in_1_bits_payload_master_xact_id,
    output io_in_0_ready,
    input  io_in_0_valid,
    input [1:0] io_in_0_bits_header_src,
    input [1:0] io_in_0_bits_header_dst,
    input [2:0] io_in_0_bits_payload_master_xact_id,
    input  io_out_ready,
    output io_out_valid,
    output[1:0] io_out_bits_header_src,
    output[1:0] io_out_bits_header_dst,
    output[2:0] io_out_bits_payload_master_xact_id,
    output[2:0] io_chosen
);

  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  reg [2:0] R17;
  wire[2:0] T18;
  wire[2:0] T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire[2:0] T33;
  wire[2:0] T34;
  wire[2:0] T35;
  wire T36;
  wire[2:0] T37;
  wire[2:0] T38;
  wire T39;
  wire T40;
  wire[2:0] T41;
  wire[2:0] T42;
  wire T43;
  wire[2:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  wire[1:0] T55;
  wire[1:0] T56;
  wire T57;
  wire[1:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[1:0] T62;
  wire[1:0] T63;
  wire[1:0] T64;
  wire T65;
  wire[1:0] T66;
  wire T67;
  wire T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R17 = {1{$random}};
  end
`endif

  assign io_chosen = T0;
  assign T0 = T1;
  assign T1 = T31 ? 3'h1 : T2;
  assign T2 = T29 ? 3'h2 : T3;
  assign T3 = T27 ? 3'h3 : T4;
  assign T4 = T25 ? 3'h4 : T5;
  assign T5 = T23 ? 3'h5 : T6;
  assign T6 = T21 ? 3'h6 : T7;
  assign T7 = T15 ? 3'h7 : T8;
  assign T8 = io_in_0_valid ? 3'h0 : T9;
  assign T9 = io_in_1_valid ? 3'h1 : T10;
  assign T10 = io_in_2_valid ? 3'h2 : T11;
  assign T11 = io_in_3_valid ? 3'h3 : T12;
  assign T12 = io_in_4_valid ? 3'h4 : T13;
  assign T13 = io_in_5_valid ? 3'h5 : T14;
  assign T14 = io_in_6_valid ? 3'h6 : 3'h7;
  assign T15 = io_in_7_valid & T16;
  assign T16 = R17 < 3'h7;
  assign T18 = reset ? 3'h0 : T19;
  assign T19 = T20 ? T0 : R17;
  assign T20 = io_out_ready & io_out_valid;
  assign T21 = io_in_6_valid & T22;
  assign T22 = R17 < 3'h6;
  assign T23 = io_in_5_valid & T24;
  assign T24 = R17 < 3'h5;
  assign T25 = io_in_4_valid & T26;
  assign T26 = R17 < 3'h4;
  assign T27 = io_in_3_valid & T28;
  assign T28 = R17 < 3'h3;
  assign T29 = io_in_2_valid & T30;
  assign T30 = R17 < 3'h2;
  assign T31 = io_in_1_valid & T32;
  assign T32 = R17 < 3'h1;
  assign io_out_bits_payload_master_xact_id = T33;
  assign T33 = T47 ? T41 : T34;
  assign T34 = T40 ? T38 : T35;
  assign T35 = T36 ? io_in_1_bits_payload_master_xact_id : io_in_0_bits_payload_master_xact_id;
  assign T36 = T37[1'h0:1'h0];
  assign T37 = T0;
  assign T38 = T39 ? io_in_3_bits_payload_master_xact_id : io_in_2_bits_payload_master_xact_id;
  assign T39 = T37[1'h0:1'h0];
  assign T40 = T37[1'h1:1'h1];
  assign T41 = T46 ? T44 : T42;
  assign T42 = T43 ? io_in_5_bits_payload_master_xact_id : io_in_4_bits_payload_master_xact_id;
  assign T43 = T37[1'h0:1'h0];
  assign T44 = T45 ? io_in_7_bits_payload_master_xact_id : io_in_6_bits_payload_master_xact_id;
  assign T45 = T37[1'h0:1'h0];
  assign T46 = T37[1'h1:1'h1];
  assign T47 = T37[2'h2:2'h2];
  assign io_out_bits_header_dst = T48;
  assign T48 = T61 ? T55 : T49;
  assign T49 = T54 ? T52 : T50;
  assign T50 = T51 ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign T51 = T37[1'h0:1'h0];
  assign T52 = T53 ? io_in_3_bits_header_dst : io_in_2_bits_header_dst;
  assign T53 = T37[1'h0:1'h0];
  assign T54 = T37[1'h1:1'h1];
  assign T55 = T60 ? T58 : T56;
  assign T56 = T57 ? io_in_5_bits_header_dst : io_in_4_bits_header_dst;
  assign T57 = T37[1'h0:1'h0];
  assign T58 = T59 ? io_in_7_bits_header_dst : io_in_6_bits_header_dst;
  assign T59 = T37[1'h0:1'h0];
  assign T60 = T37[1'h1:1'h1];
  assign T61 = T37[2'h2:2'h2];
  assign io_out_bits_header_src = T62;
  assign T62 = T75 ? T69 : T63;
  assign T63 = T68 ? T66 : T64;
  assign T64 = T65 ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign T65 = T37[1'h0:1'h0];
  assign T66 = T67 ? io_in_3_bits_header_src : io_in_2_bits_header_src;
  assign T67 = T37[1'h0:1'h0];
  assign T68 = T37[1'h1:1'h1];
  assign T69 = T74 ? T72 : T70;
  assign T70 = T71 ? io_in_5_bits_header_src : io_in_4_bits_header_src;
  assign T71 = T37[1'h0:1'h0];
  assign T72 = T73 ? io_in_7_bits_header_src : io_in_6_bits_header_src;
  assign T73 = T37[1'h0:1'h0];
  assign T74 = T37[1'h1:1'h1];
  assign T75 = T37[2'h2:2'h2];
  assign io_out_valid = T76;
  assign T76 = T89 ? T83 : T77;
  assign T77 = T82 ? T80 : T78;
  assign T78 = T79 ? io_in_1_valid : io_in_0_valid;
  assign T79 = T37[1'h0:1'h0];
  assign T80 = T81 ? io_in_3_valid : io_in_2_valid;
  assign T81 = T37[1'h0:1'h0];
  assign T82 = T37[1'h1:1'h1];
  assign T83 = T88 ? T86 : T84;
  assign T84 = T85 ? io_in_5_valid : io_in_4_valid;
  assign T85 = T37[1'h0:1'h0];
  assign T86 = T87 ? io_in_7_valid : io_in_6_valid;
  assign T87 = T37[1'h0:1'h0];
  assign T88 = T37[1'h1:1'h1];
  assign T89 = T37[2'h2:2'h2];
  assign io_in_0_ready = T90;
  assign T90 = T91 & io_out_ready;
  assign T91 = T116 | T92;
  assign T92 = T93 ^ 1'h1;
  assign T93 = T96 | T94;
  assign T94 = io_in_7_valid & T95;
  assign T95 = R17 < 3'h7;
  assign T96 = T99 | T97;
  assign T97 = io_in_6_valid & T98;
  assign T98 = R17 < 3'h6;
  assign T99 = T102 | T100;
  assign T100 = io_in_5_valid & T101;
  assign T101 = R17 < 3'h5;
  assign T102 = T105 | T103;
  assign T103 = io_in_4_valid & T104;
  assign T104 = R17 < 3'h4;
  assign T105 = T108 | T106;
  assign T106 = io_in_3_valid & T107;
  assign T107 = R17 < 3'h3;
  assign T108 = T111 | T109;
  assign T109 = io_in_2_valid & T110;
  assign T110 = R17 < 3'h2;
  assign T111 = T114 | T112;
  assign T112 = io_in_1_valid & T113;
  assign T113 = R17 < 3'h1;
  assign T114 = io_in_0_valid & T115;
  assign T115 = R17 < 3'h0;
  assign T116 = R17 < 3'h0;
  assign io_in_1_ready = T117;
  assign T117 = T118 & io_out_ready;
  assign T118 = T128 | T119;
  assign T119 = T120 ^ 1'h1;
  assign T120 = T121 | io_in_0_valid;
  assign T121 = T122 | T94;
  assign T122 = T123 | T97;
  assign T123 = T124 | T100;
  assign T124 = T125 | T103;
  assign T125 = T126 | T106;
  assign T126 = T127 | T109;
  assign T127 = T114 | T112;
  assign T128 = T130 & T129;
  assign T129 = R17 < 3'h1;
  assign T130 = T114 ^ 1'h1;
  assign io_in_2_ready = T131;
  assign T131 = T132 & io_out_ready;
  assign T132 = T143 | T133;
  assign T133 = T134 ^ 1'h1;
  assign T134 = T135 | io_in_1_valid;
  assign T135 = T136 | io_in_0_valid;
  assign T136 = T137 | T94;
  assign T137 = T138 | T97;
  assign T138 = T139 | T100;
  assign T139 = T140 | T103;
  assign T140 = T141 | T106;
  assign T141 = T142 | T109;
  assign T142 = T114 | T112;
  assign T143 = T145 & T144;
  assign T144 = R17 < 3'h2;
  assign T145 = T146 ^ 1'h1;
  assign T146 = T114 | T112;
  assign io_in_3_ready = T147;
  assign T147 = T148 & io_out_ready;
  assign T148 = T160 | T149;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T151 | io_in_2_valid;
  assign T151 = T152 | io_in_1_valid;
  assign T152 = T153 | io_in_0_valid;
  assign T153 = T154 | T94;
  assign T154 = T155 | T97;
  assign T155 = T156 | T100;
  assign T156 = T157 | T103;
  assign T157 = T158 | T106;
  assign T158 = T159 | T109;
  assign T159 = T114 | T112;
  assign T160 = T162 & T161;
  assign T161 = R17 < 3'h3;
  assign T162 = T163 ^ 1'h1;
  assign T163 = T164 | T109;
  assign T164 = T114 | T112;
  assign io_in_4_ready = T165;
  assign T165 = T166 & io_out_ready;
  assign T166 = T179 | T167;
  assign T167 = T168 ^ 1'h1;
  assign T168 = T169 | io_in_3_valid;
  assign T169 = T170 | io_in_2_valid;
  assign T170 = T171 | io_in_1_valid;
  assign T171 = T172 | io_in_0_valid;
  assign T172 = T173 | T94;
  assign T173 = T174 | T97;
  assign T174 = T175 | T100;
  assign T175 = T176 | T103;
  assign T176 = T177 | T106;
  assign T177 = T178 | T109;
  assign T178 = T114 | T112;
  assign T179 = T181 & T180;
  assign T180 = R17 < 3'h4;
  assign T181 = T182 ^ 1'h1;
  assign T182 = T183 | T106;
  assign T183 = T184 | T109;
  assign T184 = T114 | T112;
  assign io_in_5_ready = T185;
  assign T185 = T186 & io_out_ready;
  assign T186 = T200 | T187;
  assign T187 = T188 ^ 1'h1;
  assign T188 = T189 | io_in_4_valid;
  assign T189 = T190 | io_in_3_valid;
  assign T190 = T191 | io_in_2_valid;
  assign T191 = T192 | io_in_1_valid;
  assign T192 = T193 | io_in_0_valid;
  assign T193 = T194 | T94;
  assign T194 = T195 | T97;
  assign T195 = T196 | T100;
  assign T196 = T197 | T103;
  assign T197 = T198 | T106;
  assign T198 = T199 | T109;
  assign T199 = T114 | T112;
  assign T200 = T202 & T201;
  assign T201 = R17 < 3'h5;
  assign T202 = T203 ^ 1'h1;
  assign T203 = T204 | T103;
  assign T204 = T205 | T106;
  assign T205 = T206 | T109;
  assign T206 = T114 | T112;
  assign io_in_6_ready = T207;
  assign T207 = T208 & io_out_ready;
  assign T208 = T223 | T209;
  assign T209 = T210 ^ 1'h1;
  assign T210 = T211 | io_in_5_valid;
  assign T211 = T212 | io_in_4_valid;
  assign T212 = T213 | io_in_3_valid;
  assign T213 = T214 | io_in_2_valid;
  assign T214 = T215 | io_in_1_valid;
  assign T215 = T216 | io_in_0_valid;
  assign T216 = T217 | T94;
  assign T217 = T218 | T97;
  assign T218 = T219 | T100;
  assign T219 = T220 | T103;
  assign T220 = T221 | T106;
  assign T221 = T222 | T109;
  assign T222 = T114 | T112;
  assign T223 = T225 & T224;
  assign T224 = R17 < 3'h6;
  assign T225 = T226 ^ 1'h1;
  assign T226 = T227 | T100;
  assign T227 = T228 | T103;
  assign T228 = T229 | T106;
  assign T229 = T230 | T109;
  assign T230 = T114 | T112;
  assign io_in_7_ready = T231;
  assign T231 = T232 & io_out_ready;
  assign T232 = T248 | T233;
  assign T233 = T234 ^ 1'h1;
  assign T234 = T235 | io_in_6_valid;
  assign T235 = T236 | io_in_5_valid;
  assign T236 = T237 | io_in_4_valid;
  assign T237 = T238 | io_in_3_valid;
  assign T238 = T239 | io_in_2_valid;
  assign T239 = T240 | io_in_1_valid;
  assign T240 = T241 | io_in_0_valid;
  assign T241 = T242 | T94;
  assign T242 = T243 | T97;
  assign T243 = T244 | T100;
  assign T244 = T245 | T103;
  assign T245 = T246 | T106;
  assign T246 = T247 | T109;
  assign T247 = T114 | T112;
  assign T248 = T250 & T249;
  assign T249 = R17 < 3'h7;
  assign T250 = T251 ^ 1'h1;
  assign T251 = T252 | T97;
  assign T252 = T253 | T100;
  assign T253 = T254 | T103;
  assign T254 = T255 | T106;
  assign T255 = T256 | T109;
  assign T256 = T114 | T112;

  always @(posedge clk) begin
    if(reset) begin
      R17 <= 3'h0;
    end else if(T20) begin
      R17 <= T0;
    end
  end
endmodule

module UncachedTileLinkIOArbiterThatPassesId(input clk, input reset,
    output io_in_7_acquire_ready,
    input  io_in_7_acquire_valid,
    input [1:0] io_in_7_acquire_bits_header_src,
    input [1:0] io_in_7_acquire_bits_header_dst,
    input [25:0] io_in_7_acquire_bits_payload_addr,
    input [1:0] io_in_7_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_7_acquire_bits_payload_data,
    input [2:0] io_in_7_acquire_bits_payload_a_type,
    input [5:0] io_in_7_acquire_bits_payload_write_mask,
    input [2:0] io_in_7_acquire_bits_payload_subword_addr,
    input [3:0] io_in_7_acquire_bits_payload_atomic_opcode,
    input  io_in_7_grant_ready,
    output io_in_7_grant_valid,
    output[1:0] io_in_7_grant_bits_header_src,
    output[1:0] io_in_7_grant_bits_header_dst,
    output[511:0] io_in_7_grant_bits_payload_data,
    output[1:0] io_in_7_grant_bits_payload_client_xact_id,
    output[2:0] io_in_7_grant_bits_payload_master_xact_id,
    output[3:0] io_in_7_grant_bits_payload_g_type,
    output io_in_7_finish_ready,
    input  io_in_7_finish_valid,
    input [1:0] io_in_7_finish_bits_header_src,
    input [1:0] io_in_7_finish_bits_header_dst,
    input [2:0] io_in_7_finish_bits_payload_master_xact_id,
    output io_in_6_acquire_ready,
    input  io_in_6_acquire_valid,
    input [1:0] io_in_6_acquire_bits_header_src,
    input [1:0] io_in_6_acquire_bits_header_dst,
    input [25:0] io_in_6_acquire_bits_payload_addr,
    input [1:0] io_in_6_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_6_acquire_bits_payload_data,
    input [2:0] io_in_6_acquire_bits_payload_a_type,
    input [5:0] io_in_6_acquire_bits_payload_write_mask,
    input [2:0] io_in_6_acquire_bits_payload_subword_addr,
    input [3:0] io_in_6_acquire_bits_payload_atomic_opcode,
    input  io_in_6_grant_ready,
    output io_in_6_grant_valid,
    output[1:0] io_in_6_grant_bits_header_src,
    output[1:0] io_in_6_grant_bits_header_dst,
    output[511:0] io_in_6_grant_bits_payload_data,
    output[1:0] io_in_6_grant_bits_payload_client_xact_id,
    output[2:0] io_in_6_grant_bits_payload_master_xact_id,
    output[3:0] io_in_6_grant_bits_payload_g_type,
    output io_in_6_finish_ready,
    input  io_in_6_finish_valid,
    input [1:0] io_in_6_finish_bits_header_src,
    input [1:0] io_in_6_finish_bits_header_dst,
    input [2:0] io_in_6_finish_bits_payload_master_xact_id,
    output io_in_5_acquire_ready,
    input  io_in_5_acquire_valid,
    input [1:0] io_in_5_acquire_bits_header_src,
    input [1:0] io_in_5_acquire_bits_header_dst,
    input [25:0] io_in_5_acquire_bits_payload_addr,
    input [1:0] io_in_5_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_5_acquire_bits_payload_data,
    input [2:0] io_in_5_acquire_bits_payload_a_type,
    input [5:0] io_in_5_acquire_bits_payload_write_mask,
    input [2:0] io_in_5_acquire_bits_payload_subword_addr,
    input [3:0] io_in_5_acquire_bits_payload_atomic_opcode,
    input  io_in_5_grant_ready,
    output io_in_5_grant_valid,
    output[1:0] io_in_5_grant_bits_header_src,
    output[1:0] io_in_5_grant_bits_header_dst,
    output[511:0] io_in_5_grant_bits_payload_data,
    output[1:0] io_in_5_grant_bits_payload_client_xact_id,
    output[2:0] io_in_5_grant_bits_payload_master_xact_id,
    output[3:0] io_in_5_grant_bits_payload_g_type,
    output io_in_5_finish_ready,
    input  io_in_5_finish_valid,
    input [1:0] io_in_5_finish_bits_header_src,
    input [1:0] io_in_5_finish_bits_header_dst,
    input [2:0] io_in_5_finish_bits_payload_master_xact_id,
    output io_in_4_acquire_ready,
    input  io_in_4_acquire_valid,
    input [1:0] io_in_4_acquire_bits_header_src,
    input [1:0] io_in_4_acquire_bits_header_dst,
    input [25:0] io_in_4_acquire_bits_payload_addr,
    input [1:0] io_in_4_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_4_acquire_bits_payload_data,
    input [2:0] io_in_4_acquire_bits_payload_a_type,
    input [5:0] io_in_4_acquire_bits_payload_write_mask,
    input [2:0] io_in_4_acquire_bits_payload_subword_addr,
    input [3:0] io_in_4_acquire_bits_payload_atomic_opcode,
    input  io_in_4_grant_ready,
    output io_in_4_grant_valid,
    output[1:0] io_in_4_grant_bits_header_src,
    output[1:0] io_in_4_grant_bits_header_dst,
    output[511:0] io_in_4_grant_bits_payload_data,
    output[1:0] io_in_4_grant_bits_payload_client_xact_id,
    output[2:0] io_in_4_grant_bits_payload_master_xact_id,
    output[3:0] io_in_4_grant_bits_payload_g_type,
    output io_in_4_finish_ready,
    input  io_in_4_finish_valid,
    input [1:0] io_in_4_finish_bits_header_src,
    input [1:0] io_in_4_finish_bits_header_dst,
    input [2:0] io_in_4_finish_bits_payload_master_xact_id,
    output io_in_3_acquire_ready,
    input  io_in_3_acquire_valid,
    input [1:0] io_in_3_acquire_bits_header_src,
    input [1:0] io_in_3_acquire_bits_header_dst,
    input [25:0] io_in_3_acquire_bits_payload_addr,
    input [1:0] io_in_3_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_3_acquire_bits_payload_data,
    input [2:0] io_in_3_acquire_bits_payload_a_type,
    input [5:0] io_in_3_acquire_bits_payload_write_mask,
    input [2:0] io_in_3_acquire_bits_payload_subword_addr,
    input [3:0] io_in_3_acquire_bits_payload_atomic_opcode,
    input  io_in_3_grant_ready,
    output io_in_3_grant_valid,
    output[1:0] io_in_3_grant_bits_header_src,
    output[1:0] io_in_3_grant_bits_header_dst,
    output[511:0] io_in_3_grant_bits_payload_data,
    output[1:0] io_in_3_grant_bits_payload_client_xact_id,
    output[2:0] io_in_3_grant_bits_payload_master_xact_id,
    output[3:0] io_in_3_grant_bits_payload_g_type,
    output io_in_3_finish_ready,
    input  io_in_3_finish_valid,
    input [1:0] io_in_3_finish_bits_header_src,
    input [1:0] io_in_3_finish_bits_header_dst,
    input [2:0] io_in_3_finish_bits_payload_master_xact_id,
    output io_in_2_acquire_ready,
    input  io_in_2_acquire_valid,
    input [1:0] io_in_2_acquire_bits_header_src,
    input [1:0] io_in_2_acquire_bits_header_dst,
    input [25:0] io_in_2_acquire_bits_payload_addr,
    input [1:0] io_in_2_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_2_acquire_bits_payload_data,
    input [2:0] io_in_2_acquire_bits_payload_a_type,
    input [5:0] io_in_2_acquire_bits_payload_write_mask,
    input [2:0] io_in_2_acquire_bits_payload_subword_addr,
    input [3:0] io_in_2_acquire_bits_payload_atomic_opcode,
    input  io_in_2_grant_ready,
    output io_in_2_grant_valid,
    output[1:0] io_in_2_grant_bits_header_src,
    output[1:0] io_in_2_grant_bits_header_dst,
    output[511:0] io_in_2_grant_bits_payload_data,
    output[1:0] io_in_2_grant_bits_payload_client_xact_id,
    output[2:0] io_in_2_grant_bits_payload_master_xact_id,
    output[3:0] io_in_2_grant_bits_payload_g_type,
    output io_in_2_finish_ready,
    input  io_in_2_finish_valid,
    input [1:0] io_in_2_finish_bits_header_src,
    input [1:0] io_in_2_finish_bits_header_dst,
    input [2:0] io_in_2_finish_bits_payload_master_xact_id,
    output io_in_1_acquire_ready,
    input  io_in_1_acquire_valid,
    input [1:0] io_in_1_acquire_bits_header_src,
    input [1:0] io_in_1_acquire_bits_header_dst,
    input [25:0] io_in_1_acquire_bits_payload_addr,
    input [1:0] io_in_1_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_1_acquire_bits_payload_data,
    input [2:0] io_in_1_acquire_bits_payload_a_type,
    input [5:0] io_in_1_acquire_bits_payload_write_mask,
    input [2:0] io_in_1_acquire_bits_payload_subword_addr,
    input [3:0] io_in_1_acquire_bits_payload_atomic_opcode,
    input  io_in_1_grant_ready,
    output io_in_1_grant_valid,
    output[1:0] io_in_1_grant_bits_header_src,
    output[1:0] io_in_1_grant_bits_header_dst,
    output[511:0] io_in_1_grant_bits_payload_data,
    output[1:0] io_in_1_grant_bits_payload_client_xact_id,
    output[2:0] io_in_1_grant_bits_payload_master_xact_id,
    output[3:0] io_in_1_grant_bits_payload_g_type,
    output io_in_1_finish_ready,
    input  io_in_1_finish_valid,
    input [1:0] io_in_1_finish_bits_header_src,
    input [1:0] io_in_1_finish_bits_header_dst,
    input [2:0] io_in_1_finish_bits_payload_master_xact_id,
    output io_in_0_acquire_ready,
    input  io_in_0_acquire_valid,
    input [1:0] io_in_0_acquire_bits_header_src,
    input [1:0] io_in_0_acquire_bits_header_dst,
    input [25:0] io_in_0_acquire_bits_payload_addr,
    input [1:0] io_in_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_in_0_acquire_bits_payload_data,
    input [2:0] io_in_0_acquire_bits_payload_a_type,
    input [5:0] io_in_0_acquire_bits_payload_write_mask,
    input [2:0] io_in_0_acquire_bits_payload_subword_addr,
    input [3:0] io_in_0_acquire_bits_payload_atomic_opcode,
    input  io_in_0_grant_ready,
    output io_in_0_grant_valid,
    output[1:0] io_in_0_grant_bits_header_src,
    output[1:0] io_in_0_grant_bits_header_dst,
    output[511:0] io_in_0_grant_bits_payload_data,
    output[1:0] io_in_0_grant_bits_payload_client_xact_id,
    output[2:0] io_in_0_grant_bits_payload_master_xact_id,
    output[3:0] io_in_0_grant_bits_payload_g_type,
    output io_in_0_finish_ready,
    input  io_in_0_finish_valid,
    input [1:0] io_in_0_finish_bits_header_src,
    input [1:0] io_in_0_finish_bits_header_dst,
    input [2:0] io_in_0_finish_bits_payload_master_xact_id,
    input  io_out_acquire_ready,
    output io_out_acquire_valid,
    output[1:0] io_out_acquire_bits_header_src,
    output[1:0] io_out_acquire_bits_header_dst,
    output[25:0] io_out_acquire_bits_payload_addr,
    output[1:0] io_out_acquire_bits_payload_client_xact_id,
    output[511:0] io_out_acquire_bits_payload_data,
    output[2:0] io_out_acquire_bits_payload_a_type,
    output[5:0] io_out_acquire_bits_payload_write_mask,
    output[2:0] io_out_acquire_bits_payload_subword_addr,
    output[3:0] io_out_acquire_bits_payload_atomic_opcode,
    output io_out_grant_ready,
    input  io_out_grant_valid,
    input [1:0] io_out_grant_bits_header_src,
    input [1:0] io_out_grant_bits_header_dst,
    input [511:0] io_out_grant_bits_payload_data,
    input [1:0] io_out_grant_bits_payload_client_xact_id,
    input [2:0] io_out_grant_bits_payload_master_xact_id,
    input [3:0] io_out_grant_bits_payload_g_type,
    input  io_out_finish_ready,
    output io_out_finish_valid,
    output[1:0] io_out_finish_bits_header_src,
    output[1:0] io_out_finish_bits_header_dst,
    output[2:0] io_out_finish_bits_payload_master_xact_id
);

  wire[2:0] RRArbiter_1_io_out_bits_payload_master_xact_id;
  wire[1:0] RRArbiter_1_io_out_bits_header_dst;
  wire[1:0] RRArbiter_1_io_out_bits_header_src;
  wire RRArbiter_1_io_out_valid;
  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[2:0] T13;
  wire T14;
  wire[2:0] T15;
  wire T16;
  wire[2:0] T17;
  wire T18;
  wire[2:0] T19;
  wire[3:0] RRArbiter_0_io_out_bits_payload_atomic_opcode;
  wire[2:0] RRArbiter_0_io_out_bits_payload_subword_addr;
  wire[5:0] RRArbiter_0_io_out_bits_payload_write_mask;
  wire[2:0] RRArbiter_0_io_out_bits_payload_a_type;
  wire[511:0] RRArbiter_0_io_out_bits_payload_data;
  wire[1:0] RRArbiter_0_io_out_bits_payload_client_xact_id;
  wire[25:0] RRArbiter_0_io_out_bits_payload_addr;
  wire[1:0] RRArbiter_0_io_out_bits_header_dst;
  wire[1:0] RRArbiter_0_io_out_bits_header_src;
  wire RRArbiter_0_io_out_valid;
  wire RRArbiter_1_io_in_0_ready;
  wire T20;
  wire RRArbiter_0_io_in_0_ready;
  wire RRArbiter_1_io_in_1_ready;
  wire T21;
  wire RRArbiter_0_io_in_1_ready;
  wire RRArbiter_1_io_in_2_ready;
  wire T22;
  wire RRArbiter_0_io_in_2_ready;
  wire RRArbiter_1_io_in_3_ready;
  wire T23;
  wire RRArbiter_0_io_in_3_ready;
  wire RRArbiter_1_io_in_4_ready;
  wire T24;
  wire RRArbiter_0_io_in_4_ready;
  wire RRArbiter_1_io_in_5_ready;
  wire T25;
  wire RRArbiter_0_io_in_5_ready;
  wire RRArbiter_1_io_in_6_ready;
  wire T26;
  wire RRArbiter_0_io_in_6_ready;
  wire RRArbiter_1_io_in_7_ready;
  wire T27;
  wire RRArbiter_0_io_in_7_ready;


  assign io_out_finish_bits_payload_master_xact_id = RRArbiter_1_io_out_bits_payload_master_xact_id;
  assign io_out_finish_bits_header_dst = RRArbiter_1_io_out_bits_header_dst;
  assign io_out_finish_bits_header_src = RRArbiter_1_io_out_bits_header_src;
  assign io_out_finish_valid = RRArbiter_1_io_out_valid;
  assign io_out_grant_ready = T0;
  assign T0 = T18 ? io_in_7_grant_ready : T1;
  assign T1 = T16 ? io_in_6_grant_ready : T2;
  assign T2 = T14 ? io_in_5_grant_ready : T3;
  assign T3 = T12 ? io_in_4_grant_ready : T4;
  assign T4 = T11 ? io_in_3_grant_ready : T5;
  assign T5 = T10 ? io_in_2_grant_ready : T6;
  assign T6 = T9 ? io_in_1_grant_ready : T7;
  assign T7 = T8 ? io_in_0_grant_ready : 1'h0;
  assign T8 = io_out_grant_bits_payload_client_xact_id == 2'h0;
  assign T9 = io_out_grant_bits_payload_client_xact_id == 2'h1;
  assign T10 = io_out_grant_bits_payload_client_xact_id == 2'h2;
  assign T11 = io_out_grant_bits_payload_client_xact_id == 2'h3;
  assign T12 = T13 == 3'h4;
  assign T13 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T14 = T15 == 3'h5;
  assign T15 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T16 = T17 == 3'h6;
  assign T17 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign T18 = T19 == 3'h7;
  assign T19 = {1'h0, io_out_grant_bits_payload_client_xact_id};
  assign io_out_acquire_bits_payload_atomic_opcode = RRArbiter_0_io_out_bits_payload_atomic_opcode;
  assign io_out_acquire_bits_payload_subword_addr = RRArbiter_0_io_out_bits_payload_subword_addr;
  assign io_out_acquire_bits_payload_write_mask = RRArbiter_0_io_out_bits_payload_write_mask;
  assign io_out_acquire_bits_payload_a_type = RRArbiter_0_io_out_bits_payload_a_type;
  assign io_out_acquire_bits_payload_data = RRArbiter_0_io_out_bits_payload_data;
  assign io_out_acquire_bits_payload_client_xact_id = RRArbiter_0_io_out_bits_payload_client_xact_id;
  assign io_out_acquire_bits_payload_addr = RRArbiter_0_io_out_bits_payload_addr;
  assign io_out_acquire_bits_header_dst = RRArbiter_0_io_out_bits_header_dst;
  assign io_out_acquire_bits_header_src = RRArbiter_0_io_out_bits_header_src;
  assign io_out_acquire_valid = RRArbiter_0_io_out_valid;
  assign io_in_0_finish_ready = RRArbiter_1_io_in_0_ready;
  assign io_in_0_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_0_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_0_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_0_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_0_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_0_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_0_grant_valid = T20;
  assign T20 = T8 ? io_out_grant_valid : 1'h0;
  assign io_in_0_acquire_ready = RRArbiter_0_io_in_0_ready;
  assign io_in_1_finish_ready = RRArbiter_1_io_in_1_ready;
  assign io_in_1_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_1_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_1_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_1_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_1_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_1_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_1_grant_valid = T21;
  assign T21 = T9 ? io_out_grant_valid : 1'h0;
  assign io_in_1_acquire_ready = RRArbiter_0_io_in_1_ready;
  assign io_in_2_finish_ready = RRArbiter_1_io_in_2_ready;
  assign io_in_2_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_2_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_2_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_2_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_2_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_2_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_2_grant_valid = T22;
  assign T22 = T10 ? io_out_grant_valid : 1'h0;
  assign io_in_2_acquire_ready = RRArbiter_0_io_in_2_ready;
  assign io_in_3_finish_ready = RRArbiter_1_io_in_3_ready;
  assign io_in_3_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_3_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_3_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_3_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_3_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_3_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_3_grant_valid = T23;
  assign T23 = T11 ? io_out_grant_valid : 1'h0;
  assign io_in_3_acquire_ready = RRArbiter_0_io_in_3_ready;
  assign io_in_4_finish_ready = RRArbiter_1_io_in_4_ready;
  assign io_in_4_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_4_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_4_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_4_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_4_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_4_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_4_grant_valid = T24;
  assign T24 = T12 ? io_out_grant_valid : 1'h0;
  assign io_in_4_acquire_ready = RRArbiter_0_io_in_4_ready;
  assign io_in_5_finish_ready = RRArbiter_1_io_in_5_ready;
  assign io_in_5_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_5_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_5_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_5_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_5_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_5_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_5_grant_valid = T25;
  assign T25 = T14 ? io_out_grant_valid : 1'h0;
  assign io_in_5_acquire_ready = RRArbiter_0_io_in_5_ready;
  assign io_in_6_finish_ready = RRArbiter_1_io_in_6_ready;
  assign io_in_6_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_6_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_6_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_6_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_6_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_6_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_6_grant_valid = T26;
  assign T26 = T16 ? io_out_grant_valid : 1'h0;
  assign io_in_6_acquire_ready = RRArbiter_0_io_in_6_ready;
  assign io_in_7_finish_ready = RRArbiter_1_io_in_7_ready;
  assign io_in_7_grant_bits_payload_g_type = io_out_grant_bits_payload_g_type;
  assign io_in_7_grant_bits_payload_master_xact_id = io_out_grant_bits_payload_master_xact_id;
  assign io_in_7_grant_bits_payload_client_xact_id = io_out_grant_bits_payload_client_xact_id;
  assign io_in_7_grant_bits_payload_data = io_out_grant_bits_payload_data;
  assign io_in_7_grant_bits_header_dst = io_out_grant_bits_header_dst;
  assign io_in_7_grant_bits_header_src = io_out_grant_bits_header_src;
  assign io_in_7_grant_valid = T27;
  assign T27 = T18 ? io_out_grant_valid : 1'h0;
  assign io_in_7_acquire_ready = RRArbiter_0_io_in_7_ready;
  RRArbiter_3 RRArbiter_0(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_0_io_in_7_ready ),
       .io_in_7_valid( io_in_7_acquire_valid ),
       .io_in_7_bits_header_src( io_in_7_acquire_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_acquire_bits_header_dst ),
       .io_in_7_bits_payload_addr( io_in_7_acquire_bits_payload_addr ),
       .io_in_7_bits_payload_client_xact_id( io_in_7_acquire_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_data( io_in_7_acquire_bits_payload_data ),
       .io_in_7_bits_payload_a_type( io_in_7_acquire_bits_payload_a_type ),
       .io_in_7_bits_payload_write_mask( io_in_7_acquire_bits_payload_write_mask ),
       .io_in_7_bits_payload_subword_addr( io_in_7_acquire_bits_payload_subword_addr ),
       .io_in_7_bits_payload_atomic_opcode( io_in_7_acquire_bits_payload_atomic_opcode ),
       .io_in_6_ready( RRArbiter_0_io_in_6_ready ),
       .io_in_6_valid( io_in_6_acquire_valid ),
       .io_in_6_bits_header_src( io_in_6_acquire_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_acquire_bits_header_dst ),
       .io_in_6_bits_payload_addr( io_in_6_acquire_bits_payload_addr ),
       .io_in_6_bits_payload_client_xact_id( io_in_6_acquire_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_data( io_in_6_acquire_bits_payload_data ),
       .io_in_6_bits_payload_a_type( io_in_6_acquire_bits_payload_a_type ),
       .io_in_6_bits_payload_write_mask( io_in_6_acquire_bits_payload_write_mask ),
       .io_in_6_bits_payload_subword_addr( io_in_6_acquire_bits_payload_subword_addr ),
       .io_in_6_bits_payload_atomic_opcode( io_in_6_acquire_bits_payload_atomic_opcode ),
       .io_in_5_ready( RRArbiter_0_io_in_5_ready ),
       .io_in_5_valid( io_in_5_acquire_valid ),
       .io_in_5_bits_header_src( io_in_5_acquire_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_acquire_bits_header_dst ),
       .io_in_5_bits_payload_addr( io_in_5_acquire_bits_payload_addr ),
       .io_in_5_bits_payload_client_xact_id( io_in_5_acquire_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_data( io_in_5_acquire_bits_payload_data ),
       .io_in_5_bits_payload_a_type( io_in_5_acquire_bits_payload_a_type ),
       .io_in_5_bits_payload_write_mask( io_in_5_acquire_bits_payload_write_mask ),
       .io_in_5_bits_payload_subword_addr( io_in_5_acquire_bits_payload_subword_addr ),
       .io_in_5_bits_payload_atomic_opcode( io_in_5_acquire_bits_payload_atomic_opcode ),
       .io_in_4_ready( RRArbiter_0_io_in_4_ready ),
       .io_in_4_valid( io_in_4_acquire_valid ),
       .io_in_4_bits_header_src( io_in_4_acquire_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_acquire_bits_header_dst ),
       .io_in_4_bits_payload_addr( io_in_4_acquire_bits_payload_addr ),
       .io_in_4_bits_payload_client_xact_id( io_in_4_acquire_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_data( io_in_4_acquire_bits_payload_data ),
       .io_in_4_bits_payload_a_type( io_in_4_acquire_bits_payload_a_type ),
       .io_in_4_bits_payload_write_mask( io_in_4_acquire_bits_payload_write_mask ),
       .io_in_4_bits_payload_subword_addr( io_in_4_acquire_bits_payload_subword_addr ),
       .io_in_4_bits_payload_atomic_opcode( io_in_4_acquire_bits_payload_atomic_opcode ),
       .io_in_3_ready( RRArbiter_0_io_in_3_ready ),
       .io_in_3_valid( io_in_3_acquire_valid ),
       .io_in_3_bits_header_src( io_in_3_acquire_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_acquire_bits_header_dst ),
       .io_in_3_bits_payload_addr( io_in_3_acquire_bits_payload_addr ),
       .io_in_3_bits_payload_client_xact_id( io_in_3_acquire_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_data( io_in_3_acquire_bits_payload_data ),
       .io_in_3_bits_payload_a_type( io_in_3_acquire_bits_payload_a_type ),
       .io_in_3_bits_payload_write_mask( io_in_3_acquire_bits_payload_write_mask ),
       .io_in_3_bits_payload_subword_addr( io_in_3_acquire_bits_payload_subword_addr ),
       .io_in_3_bits_payload_atomic_opcode( io_in_3_acquire_bits_payload_atomic_opcode ),
       .io_in_2_ready( RRArbiter_0_io_in_2_ready ),
       .io_in_2_valid( io_in_2_acquire_valid ),
       .io_in_2_bits_header_src( io_in_2_acquire_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_acquire_bits_header_dst ),
       .io_in_2_bits_payload_addr( io_in_2_acquire_bits_payload_addr ),
       .io_in_2_bits_payload_client_xact_id( io_in_2_acquire_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_data( io_in_2_acquire_bits_payload_data ),
       .io_in_2_bits_payload_a_type( io_in_2_acquire_bits_payload_a_type ),
       .io_in_2_bits_payload_write_mask( io_in_2_acquire_bits_payload_write_mask ),
       .io_in_2_bits_payload_subword_addr( io_in_2_acquire_bits_payload_subword_addr ),
       .io_in_2_bits_payload_atomic_opcode( io_in_2_acquire_bits_payload_atomic_opcode ),
       .io_in_1_ready( RRArbiter_0_io_in_1_ready ),
       .io_in_1_valid( io_in_1_acquire_valid ),
       .io_in_1_bits_header_src( io_in_1_acquire_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_acquire_bits_header_dst ),
       .io_in_1_bits_payload_addr( io_in_1_acquire_bits_payload_addr ),
       .io_in_1_bits_payload_client_xact_id( io_in_1_acquire_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_data( io_in_1_acquire_bits_payload_data ),
       .io_in_1_bits_payload_a_type( io_in_1_acquire_bits_payload_a_type ),
       .io_in_1_bits_payload_write_mask( io_in_1_acquire_bits_payload_write_mask ),
       .io_in_1_bits_payload_subword_addr( io_in_1_acquire_bits_payload_subword_addr ),
       .io_in_1_bits_payload_atomic_opcode( io_in_1_acquire_bits_payload_atomic_opcode ),
       .io_in_0_ready( RRArbiter_0_io_in_0_ready ),
       .io_in_0_valid( io_in_0_acquire_valid ),
       .io_in_0_bits_header_src( io_in_0_acquire_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_acquire_bits_header_dst ),
       .io_in_0_bits_payload_addr( io_in_0_acquire_bits_payload_addr ),
       .io_in_0_bits_payload_client_xact_id( io_in_0_acquire_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_data( io_in_0_acquire_bits_payload_data ),
       .io_in_0_bits_payload_a_type( io_in_0_acquire_bits_payload_a_type ),
       .io_in_0_bits_payload_write_mask( io_in_0_acquire_bits_payload_write_mask ),
       .io_in_0_bits_payload_subword_addr( io_in_0_acquire_bits_payload_subword_addr ),
       .io_in_0_bits_payload_atomic_opcode( io_in_0_acquire_bits_payload_atomic_opcode ),
       .io_out_ready( io_out_acquire_ready ),
       .io_out_valid( RRArbiter_0_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_0_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_0_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( RRArbiter_0_io_out_bits_payload_addr ),
       .io_out_bits_payload_client_xact_id( RRArbiter_0_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_data( RRArbiter_0_io_out_bits_payload_data ),
       .io_out_bits_payload_a_type( RRArbiter_0_io_out_bits_payload_a_type ),
       .io_out_bits_payload_write_mask( RRArbiter_0_io_out_bits_payload_write_mask ),
       .io_out_bits_payload_subword_addr( RRArbiter_0_io_out_bits_payload_subword_addr ),
       .io_out_bits_payload_atomic_opcode( RRArbiter_0_io_out_bits_payload_atomic_opcode )
       //.io_chosen(  )
  );
  RRArbiter_4 RRArbiter_1(.clk(clk), .reset(reset),
       .io_in_7_ready( RRArbiter_1_io_in_7_ready ),
       .io_in_7_valid( io_in_7_finish_valid ),
       .io_in_7_bits_header_src( io_in_7_finish_bits_header_src ),
       .io_in_7_bits_header_dst( io_in_7_finish_bits_header_dst ),
       .io_in_7_bits_payload_master_xact_id( io_in_7_finish_bits_payload_master_xact_id ),
       .io_in_6_ready( RRArbiter_1_io_in_6_ready ),
       .io_in_6_valid( io_in_6_finish_valid ),
       .io_in_6_bits_header_src( io_in_6_finish_bits_header_src ),
       .io_in_6_bits_header_dst( io_in_6_finish_bits_header_dst ),
       .io_in_6_bits_payload_master_xact_id( io_in_6_finish_bits_payload_master_xact_id ),
       .io_in_5_ready( RRArbiter_1_io_in_5_ready ),
       .io_in_5_valid( io_in_5_finish_valid ),
       .io_in_5_bits_header_src( io_in_5_finish_bits_header_src ),
       .io_in_5_bits_header_dst( io_in_5_finish_bits_header_dst ),
       .io_in_5_bits_payload_master_xact_id( io_in_5_finish_bits_payload_master_xact_id ),
       .io_in_4_ready( RRArbiter_1_io_in_4_ready ),
       .io_in_4_valid( io_in_4_finish_valid ),
       .io_in_4_bits_header_src( io_in_4_finish_bits_header_src ),
       .io_in_4_bits_header_dst( io_in_4_finish_bits_header_dst ),
       .io_in_4_bits_payload_master_xact_id( io_in_4_finish_bits_payload_master_xact_id ),
       .io_in_3_ready( RRArbiter_1_io_in_3_ready ),
       .io_in_3_valid( io_in_3_finish_valid ),
       .io_in_3_bits_header_src( io_in_3_finish_bits_header_src ),
       .io_in_3_bits_header_dst( io_in_3_finish_bits_header_dst ),
       .io_in_3_bits_payload_master_xact_id( io_in_3_finish_bits_payload_master_xact_id ),
       .io_in_2_ready( RRArbiter_1_io_in_2_ready ),
       .io_in_2_valid( io_in_2_finish_valid ),
       .io_in_2_bits_header_src( io_in_2_finish_bits_header_src ),
       .io_in_2_bits_header_dst( io_in_2_finish_bits_header_dst ),
       .io_in_2_bits_payload_master_xact_id( io_in_2_finish_bits_payload_master_xact_id ),
       .io_in_1_ready( RRArbiter_1_io_in_1_ready ),
       .io_in_1_valid( io_in_1_finish_valid ),
       .io_in_1_bits_header_src( io_in_1_finish_bits_header_src ),
       .io_in_1_bits_header_dst( io_in_1_finish_bits_header_dst ),
       .io_in_1_bits_payload_master_xact_id( io_in_1_finish_bits_payload_master_xact_id ),
       .io_in_0_ready( RRArbiter_1_io_in_0_ready ),
       .io_in_0_valid( io_in_0_finish_valid ),
       .io_in_0_bits_header_src( io_in_0_finish_bits_header_src ),
       .io_in_0_bits_header_dst( io_in_0_finish_bits_header_dst ),
       .io_in_0_bits_payload_master_xact_id( io_in_0_finish_bits_payload_master_xact_id ),
       .io_out_ready( io_out_finish_ready ),
       .io_out_valid( RRArbiter_1_io_out_valid ),
       .io_out_bits_header_src( RRArbiter_1_io_out_bits_header_src ),
       .io_out_bits_header_dst( RRArbiter_1_io_out_bits_header_dst ),
       .io_out_bits_payload_master_xact_id( RRArbiter_1_io_out_bits_payload_master_xact_id )
       //.io_chosen(  )
  );
endmodule

module L2CoherenceAgent(input clk, input reset,
    output io_inner_acquire_ready,
    input  io_inner_acquire_valid,
    input [1:0] io_inner_acquire_bits_header_src,
    input [1:0] io_inner_acquire_bits_header_dst,
    input [25:0] io_inner_acquire_bits_payload_addr,
    input [1:0] io_inner_acquire_bits_payload_client_xact_id,
    input [511:0] io_inner_acquire_bits_payload_data,
    input [2:0] io_inner_acquire_bits_payload_a_type,
    input [5:0] io_inner_acquire_bits_payload_write_mask,
    input [2:0] io_inner_acquire_bits_payload_subword_addr,
    input [3:0] io_inner_acquire_bits_payload_atomic_opcode,
    input  io_inner_grant_ready,
    output io_inner_grant_valid,
    output[1:0] io_inner_grant_bits_header_src,
    output[1:0] io_inner_grant_bits_header_dst,
    output[511:0] io_inner_grant_bits_payload_data,
    output[1:0] io_inner_grant_bits_payload_client_xact_id,
    output[2:0] io_inner_grant_bits_payload_master_xact_id,
    output[3:0] io_inner_grant_bits_payload_g_type,
    output io_inner_finish_ready,
    input  io_inner_finish_valid,
    input [1:0] io_inner_finish_bits_header_src,
    input [1:0] io_inner_finish_bits_header_dst,
    input [2:0] io_inner_finish_bits_payload_master_xact_id,
    input  io_inner_probe_ready,
    output io_inner_probe_valid,
    output[1:0] io_inner_probe_bits_header_src,
    output[1:0] io_inner_probe_bits_header_dst,
    output[25:0] io_inner_probe_bits_payload_addr,
    output[2:0] io_inner_probe_bits_payload_master_xact_id,
    output[1:0] io_inner_probe_bits_payload_p_type,
    output io_inner_release_ready,
    input  io_inner_release_valid,
    input [1:0] io_inner_release_bits_header_src,
    input [1:0] io_inner_release_bits_header_dst,
    input [25:0] io_inner_release_bits_payload_addr,
    input [1:0] io_inner_release_bits_payload_client_xact_id,
    input [2:0] io_inner_release_bits_payload_master_xact_id,
    input [511:0] io_inner_release_bits_payload_data,
    input [2:0] io_inner_release_bits_payload_r_type,
    input  io_outer_acquire_ready,
    output io_outer_acquire_valid,
    output[1:0] io_outer_acquire_bits_header_src,
    output[1:0] io_outer_acquire_bits_header_dst,
    output[25:0] io_outer_acquire_bits_payload_addr,
    output[1:0] io_outer_acquire_bits_payload_client_xact_id,
    output[511:0] io_outer_acquire_bits_payload_data,
    output[2:0] io_outer_acquire_bits_payload_a_type,
    output[5:0] io_outer_acquire_bits_payload_write_mask,
    output[2:0] io_outer_acquire_bits_payload_subword_addr,
    output[3:0] io_outer_acquire_bits_payload_atomic_opcode,
    output io_outer_grant_ready,
    input  io_outer_grant_valid,
    input [1:0] io_outer_grant_bits_header_src,
    input [1:0] io_outer_grant_bits_header_dst,
    input [511:0] io_outer_grant_bits_payload_data,
    input [1:0] io_outer_grant_bits_payload_client_xact_id,
    input [2:0] io_outer_grant_bits_payload_master_xact_id,
    input [3:0] io_outer_grant_bits_payload_g_type,
    input  io_outer_finish_ready,
    output io_outer_finish_valid,
    output[1:0] io_outer_finish_bits_header_src,
    output[1:0] io_outer_finish_bits_header_dst,
    output[2:0] io_outer_finish_bits_payload_master_xact_id,
    input  io_incoherent_1,
    input  io_incoherent_0
);

  wire VoluntaryReleaseTracker_io_outer_grant_ready;
  wire[3:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type;
  wire[511:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr;
  wire[1:0] VoluntaryReleaseTracker_io_outer_acquire_bits_header_src;
  wire VoluntaryReleaseTracker_io_outer_acquire_valid;
  wire AcquireTracker_0_io_outer_grant_ready;
  wire[3:0] AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_0_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_0_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_0_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_0_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_outer_acquire_bits_header_src;
  wire AcquireTracker_0_io_outer_acquire_valid;
  wire AcquireTracker_1_io_outer_grant_ready;
  wire[3:0] AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_1_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_1_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_1_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_1_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_outer_acquire_bits_header_src;
  wire AcquireTracker_1_io_outer_acquire_valid;
  wire AcquireTracker_2_io_outer_grant_ready;
  wire[3:0] AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_2_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_2_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_2_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_2_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_outer_acquire_bits_header_src;
  wire AcquireTracker_2_io_outer_acquire_valid;
  wire AcquireTracker_3_io_outer_grant_ready;
  wire[3:0] AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_3_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_3_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_3_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_3_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_outer_acquire_bits_header_src;
  wire AcquireTracker_3_io_outer_acquire_valid;
  wire AcquireTracker_4_io_outer_grant_ready;
  wire[3:0] AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_4_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_4_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_4_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_4_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_4_io_outer_acquire_bits_header_src;
  wire AcquireTracker_4_io_outer_acquire_valid;
  wire AcquireTracker_5_io_outer_grant_ready;
  wire[3:0] AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_5_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_5_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_5_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_5_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_5_io_outer_acquire_bits_header_src;
  wire AcquireTracker_5_io_outer_acquire_valid;
  wire AcquireTracker_6_io_outer_grant_ready;
  wire[3:0] AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] AcquireTracker_6_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] AcquireTracker_6_io_outer_acquire_bits_payload_a_type;
  wire[511:0] AcquireTracker_6_io_outer_acquire_bits_payload_data;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] AcquireTracker_6_io_outer_acquire_bits_payload_addr;
  wire[1:0] AcquireTracker_6_io_outer_acquire_bits_header_src;
  wire AcquireTracker_6_io_outer_acquire_valid;
  wire[3:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type;
  wire[2:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] VoluntaryReleaseTracker_io_inner_grant_bits_payload_data;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_dst;
  wire[1:0] VoluntaryReleaseTracker_io_inner_grant_bits_header_src;
  wire VoluntaryReleaseTracker_io_inner_grant_valid;
  wire[3:0] AcquireTracker_0_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_0_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_0_io_inner_grant_bits_header_src;
  wire AcquireTracker_0_io_inner_grant_valid;
  wire[3:0] AcquireTracker_1_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_1_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_1_io_inner_grant_bits_header_src;
  wire AcquireTracker_1_io_inner_grant_valid;
  wire[3:0] AcquireTracker_2_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_2_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_2_io_inner_grant_bits_header_src;
  wire AcquireTracker_2_io_inner_grant_valid;
  wire[3:0] AcquireTracker_3_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_3_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_3_io_inner_grant_bits_header_src;
  wire AcquireTracker_3_io_inner_grant_valid;
  wire[3:0] AcquireTracker_4_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_4_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_4_io_inner_grant_bits_header_src;
  wire AcquireTracker_4_io_inner_grant_valid;
  wire[3:0] AcquireTracker_5_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_5_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_5_io_inner_grant_bits_header_src;
  wire AcquireTracker_5_io_inner_grant_valid;
  wire[3:0] AcquireTracker_6_io_inner_grant_bits_payload_g_type;
  wire[2:0] AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] AcquireTracker_6_io_inner_grant_bits_payload_data;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_dst;
  wire[1:0] AcquireTracker_6_io_inner_grant_bits_header_src;
  wire AcquireTracker_6_io_inner_grant_valid;
  wire VoluntaryReleaseTracker_io_inner_probe_valid;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_0_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_0_io_inner_probe_bits_header_src;
  wire AcquireTracker_0_io_inner_probe_valid;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_1_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_1_io_inner_probe_bits_header_src;
  wire AcquireTracker_1_io_inner_probe_valid;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_2_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_2_io_inner_probe_bits_header_src;
  wire AcquireTracker_2_io_inner_probe_valid;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_3_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_3_io_inner_probe_bits_header_src;
  wire AcquireTracker_3_io_inner_probe_valid;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_4_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_4_io_inner_probe_bits_header_src;
  wire AcquireTracker_4_io_inner_probe_valid;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_5_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_5_io_inner_probe_bits_header_src;
  wire AcquireTracker_5_io_inner_probe_valid;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_payload_p_type;
  wire[2:0] AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] AcquireTracker_6_io_inner_probe_bits_payload_addr;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_dst;
  wire[1:0] AcquireTracker_6_io_inner_probe_bits_header_src;
  wire AcquireTracker_6_io_inner_probe_valid;
  wire T0;
  wire T1;
  wire block_acquires;
  wire AcquireTracker_6_io_has_acquire_conflict;
  wire T2;
  wire AcquireTracker_5_io_has_acquire_conflict;
  wire T3;
  wire AcquireTracker_4_io_has_acquire_conflict;
  wire T4;
  wire AcquireTracker_3_io_has_acquire_conflict;
  wire T5;
  wire AcquireTracker_2_io_has_acquire_conflict;
  wire T6;
  wire AcquireTracker_1_io_has_acquire_conflict;
  wire T7;
  wire AcquireTracker_0_io_has_acquire_conflict;
  wire VoluntaryReleaseTracker_io_has_acquire_conflict;
  wire VoluntaryReleaseTracker_io_inner_acquire_ready;
  wire AcquireTracker_0_io_inner_acquire_ready;
  wire AcquireTracker_1_io_inner_acquire_ready;
  wire AcquireTracker_2_io_inner_acquire_ready;
  wire AcquireTracker_3_io_inner_acquire_ready;
  wire AcquireTracker_4_io_inner_acquire_ready;
  wire AcquireTracker_5_io_inner_acquire_ready;
  wire AcquireTracker_6_io_inner_acquire_ready;
  wire[1:0] T8;
  wire[1:0] T9;
  wire outer_arb_io_in_7_finish_ready;
  wire[3:0] outer_arb_io_in_7_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_7_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_7_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_7_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_7_grant_bits_header_src;
  wire outer_arb_io_in_7_grant_valid;
  wire outer_arb_io_in_7_acquire_ready;
  wire T10;
  wire T11;
  wire[2:0] release_idx;
  wire voluntary;
  wire probe_arb_io_in_7_ready;
  wire grant_arb_io_in_7_ready;
  wire alloc_arb_io_in_7_ready;
  wire[1:0] T12;
  wire outer_arb_io_in_6_finish_ready;
  wire[3:0] outer_arb_io_in_6_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_6_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_6_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_6_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_6_grant_bits_header_src;
  wire outer_arb_io_in_6_grant_valid;
  wire outer_arb_io_in_6_acquire_ready;
  wire T13;
  wire T14;
  wire probe_arb_io_in_6_ready;
  wire grant_arb_io_in_6_ready;
  wire alloc_arb_io_in_6_ready;
  wire[1:0] T15;
  wire outer_arb_io_in_5_finish_ready;
  wire[3:0] outer_arb_io_in_5_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_5_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_5_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_5_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_5_grant_bits_header_src;
  wire outer_arb_io_in_5_grant_valid;
  wire outer_arb_io_in_5_acquire_ready;
  wire T16;
  wire T17;
  wire probe_arb_io_in_5_ready;
  wire grant_arb_io_in_5_ready;
  wire alloc_arb_io_in_5_ready;
  wire[1:0] T18;
  wire outer_arb_io_in_4_finish_ready;
  wire[3:0] outer_arb_io_in_4_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_4_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_4_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_4_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_4_grant_bits_header_src;
  wire outer_arb_io_in_4_grant_valid;
  wire outer_arb_io_in_4_acquire_ready;
  wire T19;
  wire T20;
  wire probe_arb_io_in_4_ready;
  wire grant_arb_io_in_4_ready;
  wire alloc_arb_io_in_4_ready;
  wire[1:0] T21;
  wire outer_arb_io_in_3_finish_ready;
  wire[3:0] outer_arb_io_in_3_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_3_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_3_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_3_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_3_grant_bits_header_src;
  wire outer_arb_io_in_3_grant_valid;
  wire outer_arb_io_in_3_acquire_ready;
  wire T22;
  wire T23;
  wire probe_arb_io_in_3_ready;
  wire grant_arb_io_in_3_ready;
  wire alloc_arb_io_in_3_ready;
  wire[1:0] T24;
  wire outer_arb_io_in_2_finish_ready;
  wire[3:0] outer_arb_io_in_2_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_2_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_2_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_2_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_2_grant_bits_header_src;
  wire outer_arb_io_in_2_grant_valid;
  wire outer_arb_io_in_2_acquire_ready;
  wire T25;
  wire T26;
  wire probe_arb_io_in_2_ready;
  wire grant_arb_io_in_2_ready;
  wire alloc_arb_io_in_2_ready;
  wire[1:0] T27;
  wire outer_arb_io_in_1_finish_ready;
  wire[3:0] outer_arb_io_in_1_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_1_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_1_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_1_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_1_grant_bits_header_src;
  wire outer_arb_io_in_1_grant_valid;
  wire outer_arb_io_in_1_acquire_ready;
  wire T28;
  wire T29;
  wire probe_arb_io_in_1_ready;
  wire grant_arb_io_in_1_ready;
  wire alloc_arb_io_in_1_ready;
  wire[1:0] T30;
  wire outer_arb_io_in_0_finish_ready;
  wire[3:0] outer_arb_io_in_0_grant_bits_payload_g_type;
  wire[2:0] outer_arb_io_in_0_grant_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_in_0_grant_bits_payload_client_xact_id;
  wire[511:0] outer_arb_io_in_0_grant_bits_payload_data;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_dst;
  wire[1:0] outer_arb_io_in_0_grant_bits_header_src;
  wire outer_arb_io_in_0_grant_valid;
  wire outer_arb_io_in_0_acquire_ready;
  wire T31;
  wire T32;
  wire probe_arb_io_in_0_ready;
  wire grant_arb_io_in_0_ready;
  wire alloc_arb_io_in_0_ready;
  wire[2:0] outer_arb_io_out_finish_bits_payload_master_xact_id;
  wire[1:0] outer_arb_io_out_finish_bits_header_dst;
  wire[1:0] outer_arb_io_out_finish_bits_header_src;
  wire outer_arb_io_out_finish_valid;
  wire outer_arb_io_out_grant_ready;
  wire[3:0] outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_subword_addr;
  wire[5:0] outer_arb_io_out_acquire_bits_payload_write_mask;
  wire[2:0] outer_arb_io_out_acquire_bits_payload_a_type;
  wire[511:0] outer_arb_io_out_acquire_bits_payload_data;
  wire[1:0] outer_arb_io_out_acquire_bits_payload_client_xact_id;
  wire[25:0] outer_arb_io_out_acquire_bits_payload_addr;
  wire[1:0] outer_arb_io_out_acquire_bits_header_dst;
  wire[1:0] outer_arb_io_out_acquire_bits_header_src;
  wire outer_arb_io_out_acquire_valid;
  wire T33;
  wire T34;
  wire T35;
  wire VoluntaryReleaseTracker_io_inner_release_ready;
  wire AcquireTracker_0_io_inner_release_ready;
  wire T36;
  wire[2:0] T37;
  wire T38;
  wire AcquireTracker_1_io_inner_release_ready;
  wire AcquireTracker_2_io_inner_release_ready;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire AcquireTracker_3_io_inner_release_ready;
  wire AcquireTracker_4_io_inner_release_ready;
  wire T43;
  wire T44;
  wire AcquireTracker_5_io_inner_release_ready;
  wire AcquireTracker_6_io_inner_release_ready;
  wire T45;
  wire T46;
  wire T47;
  wire[1:0] probe_arb_io_out_bits_payload_p_type;
  wire[2:0] probe_arb_io_out_bits_payload_master_xact_id;
  wire[25:0] probe_arb_io_out_bits_payload_addr;
  wire[1:0] probe_arb_io_out_bits_header_dst;
  wire[1:0] probe_arb_io_out_bits_header_src;
  wire probe_arb_io_out_valid;
  wire[3:0] grant_arb_io_out_bits_payload_g_type;
  wire[2:0] grant_arb_io_out_bits_payload_master_xact_id;
  wire[1:0] grant_arb_io_out_bits_payload_client_xact_id;
  wire[511:0] grant_arb_io_out_bits_payload_data;
  wire[1:0] grant_arb_io_out_bits_header_dst;
  wire[1:0] grant_arb_io_out_bits_header_src;
  wire grant_arb_io_out_valid;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;


  assign T0 = io_inner_acquire_valid & T1;
  assign T1 = block_acquires ^ 1'h1;
  assign block_acquires = T2 | AcquireTracker_6_io_has_acquire_conflict;
  assign T2 = T3 | AcquireTracker_5_io_has_acquire_conflict;
  assign T3 = T4 | AcquireTracker_4_io_has_acquire_conflict;
  assign T4 = T5 | AcquireTracker_3_io_has_acquire_conflict;
  assign T5 = T6 | AcquireTracker_2_io_has_acquire_conflict;
  assign T6 = T7 | AcquireTracker_1_io_has_acquire_conflict;
  assign T7 = VoluntaryReleaseTracker_io_has_acquire_conflict | AcquireTracker_0_io_has_acquire_conflict;
  assign T8 = T9;
  assign T9 = {io_incoherent_1, io_incoherent_0};
  assign T10 = io_inner_release_valid & T11;
  assign T11 = release_idx == 3'h7;
  assign release_idx = voluntary ? 3'h0 : io_inner_release_bits_payload_master_xact_id;
  assign voluntary = io_inner_release_bits_payload_r_type == 3'h0;
  assign T12 = T9;
  assign T13 = io_inner_release_valid & T14;
  assign T14 = release_idx == 3'h6;
  assign T15 = T9;
  assign T16 = io_inner_release_valid & T17;
  assign T17 = release_idx == 3'h5;
  assign T18 = T9;
  assign T19 = io_inner_release_valid & T20;
  assign T20 = release_idx == 3'h4;
  assign T21 = T9;
  assign T22 = io_inner_release_valid & T23;
  assign T23 = release_idx == 3'h3;
  assign T24 = T9;
  assign T25 = io_inner_release_valid & T26;
  assign T26 = release_idx == 3'h2;
  assign T27 = T9;
  assign T28 = io_inner_release_valid & T29;
  assign T29 = release_idx == 3'h1;
  assign T30 = T9;
  assign T31 = io_inner_release_valid & T32;
  assign T32 = release_idx == 3'h0;
  assign io_outer_finish_bits_payload_master_xact_id = outer_arb_io_out_finish_bits_payload_master_xact_id;
  assign io_outer_finish_bits_header_dst = outer_arb_io_out_finish_bits_header_dst;
  assign io_outer_finish_bits_header_src = outer_arb_io_out_finish_bits_header_src;
  assign io_outer_finish_valid = outer_arb_io_out_finish_valid;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign io_outer_acquire_bits_payload_atomic_opcode = outer_arb_io_out_acquire_bits_payload_atomic_opcode;
  assign io_outer_acquire_bits_payload_subword_addr = outer_arb_io_out_acquire_bits_payload_subword_addr;
  assign io_outer_acquire_bits_payload_write_mask = outer_arb_io_out_acquire_bits_payload_write_mask;
  assign io_outer_acquire_bits_payload_a_type = outer_arb_io_out_acquire_bits_payload_a_type;
  assign io_outer_acquire_bits_payload_data = outer_arb_io_out_acquire_bits_payload_data;
  assign io_outer_acquire_bits_payload_client_xact_id = outer_arb_io_out_acquire_bits_payload_client_xact_id;
  assign io_outer_acquire_bits_payload_addr = outer_arb_io_out_acquire_bits_payload_addr;
  assign io_outer_acquire_bits_header_dst = outer_arb_io_out_acquire_bits_header_dst;
  assign io_outer_acquire_bits_header_src = outer_arb_io_out_acquire_bits_header_src;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_inner_release_ready = T33;
  assign T33 = T47 ? T41 : T34;
  assign T34 = T40 ? T38 : T35;
  assign T35 = T36 ? AcquireTracker_0_io_inner_release_ready : VoluntaryReleaseTracker_io_inner_release_ready;
  assign T36 = T37[1'h0:1'h0];
  assign T37 = release_idx;
  assign T38 = T39 ? AcquireTracker_2_io_inner_release_ready : AcquireTracker_1_io_inner_release_ready;
  assign T39 = T37[1'h0:1'h0];
  assign T40 = T37[1'h1:1'h1];
  assign T41 = T46 ? T44 : T42;
  assign T42 = T43 ? AcquireTracker_4_io_inner_release_ready : AcquireTracker_3_io_inner_release_ready;
  assign T43 = T37[1'h0:1'h0];
  assign T44 = T45 ? AcquireTracker_6_io_inner_release_ready : AcquireTracker_5_io_inner_release_ready;
  assign T45 = T37[1'h0:1'h0];
  assign T46 = T37[1'h1:1'h1];
  assign T47 = T37[2'h2:2'h2];
  assign io_inner_probe_bits_payload_p_type = probe_arb_io_out_bits_payload_p_type;
  assign io_inner_probe_bits_payload_master_xact_id = probe_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_probe_bits_payload_addr = probe_arb_io_out_bits_payload_addr;
  assign io_inner_probe_bits_header_dst = probe_arb_io_out_bits_header_dst;
  assign io_inner_probe_bits_header_src = probe_arb_io_out_bits_header_src;
  assign io_inner_probe_valid = probe_arb_io_out_valid;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_grant_bits_payload_g_type = grant_arb_io_out_bits_payload_g_type;
  assign io_inner_grant_bits_payload_master_xact_id = grant_arb_io_out_bits_payload_master_xact_id;
  assign io_inner_grant_bits_payload_client_xact_id = grant_arb_io_out_bits_payload_client_xact_id;
  assign io_inner_grant_bits_payload_data = grant_arb_io_out_bits_payload_data;
  assign io_inner_grant_bits_header_dst = grant_arb_io_out_bits_header_dst;
  assign io_inner_grant_bits_header_src = grant_arb_io_out_bits_header_src;
  assign io_inner_grant_valid = grant_arb_io_out_valid;
  assign io_inner_acquire_ready = T48;
  assign T48 = T50 & T49;
  assign T49 = block_acquires ^ 1'h1;
  assign T50 = T51 | AcquireTracker_6_io_inner_acquire_ready;
  assign T51 = T52 | AcquireTracker_5_io_inner_acquire_ready;
  assign T52 = T53 | AcquireTracker_4_io_inner_acquire_ready;
  assign T53 = T54 | AcquireTracker_3_io_inner_acquire_ready;
  assign T54 = T55 | AcquireTracker_2_io_inner_acquire_ready;
  assign T55 = T56 | AcquireTracker_1_io_inner_acquire_ready;
  assign T56 = VoluntaryReleaseTracker_io_inner_acquire_ready | AcquireTracker_0_io_inner_acquire_ready;
  VoluntaryReleaseTracker VoluntaryReleaseTracker(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_0_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_0_ready ),
       .io_inner_grant_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_0_ready ),
       .io_inner_probe_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_inner_probe_bits_header_src(  )
       //.io_inner_probe_bits_header_dst(  )
       //.io_inner_probe_bits_payload_addr(  )
       //.io_inner_probe_bits_payload_master_xact_id(  )
       //.io_inner_probe_bits_payload_p_type(  )
       .io_inner_release_ready( VoluntaryReleaseTracker_io_inner_release_ready ),
       .io_inner_release_valid( T31 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_outer_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T30 ),
       .io_has_acquire_conflict( VoluntaryReleaseTracker_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_0 AcquireTracker_0(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_0_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_1_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_1_ready ),
       .io_inner_grant_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_1_ready ),
       .io_inner_probe_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_0_io_inner_release_ready ),
       .io_inner_release_valid( T28 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T27 ),
       .io_has_acquire_conflict( AcquireTracker_0_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_1 AcquireTracker_1(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_1_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_2_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_2_ready ),
       .io_inner_grant_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_2_ready ),
       .io_inner_probe_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_1_io_inner_release_ready ),
       .io_inner_release_valid( T25 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T24 ),
       .io_has_acquire_conflict( AcquireTracker_1_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_2 AcquireTracker_2(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_2_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_3_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_3_ready ),
       .io_inner_grant_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_3_ready ),
       .io_inner_probe_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_2_io_inner_release_ready ),
       .io_inner_release_valid( T22 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T21 ),
       .io_has_acquire_conflict( AcquireTracker_2_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_3 AcquireTracker_3(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_3_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_4_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_4_ready ),
       .io_inner_grant_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_4_ready ),
       .io_inner_probe_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_3_io_inner_release_ready ),
       .io_inner_release_valid( T19 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T18 ),
       .io_has_acquire_conflict( AcquireTracker_3_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_4 AcquireTracker_4(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_4_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_5_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_5_ready ),
       .io_inner_grant_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_5_ready ),
       .io_inner_probe_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_4_io_inner_release_ready ),
       .io_inner_release_valid( T16 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T15 ),
       .io_has_acquire_conflict( AcquireTracker_4_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_5 AcquireTracker_5(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_5_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_6_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_6_ready ),
       .io_inner_grant_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_6_ready ),
       .io_inner_probe_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_5_io_inner_release_ready ),
       .io_inner_release_valid( T13 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T12 ),
       .io_has_acquire_conflict( AcquireTracker_5_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  AcquireTracker_6 AcquireTracker_6(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( AcquireTracker_6_io_inner_acquire_ready ),
       .io_inner_acquire_valid( alloc_arb_io_in_7_ready ),
       .io_inner_acquire_bits_header_src( io_inner_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( io_inner_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( io_inner_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( io_inner_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( io_inner_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( io_inner_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( io_inner_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( io_inner_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( io_inner_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( grant_arb_io_in_7_ready ),
       .io_inner_grant_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       //.io_inner_finish_ready(  )
       .io_inner_finish_valid( io_inner_finish_valid ),
       .io_inner_finish_bits_header_src( io_inner_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( io_inner_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( io_inner_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( probe_arb_io_in_7_ready ),
       .io_inner_probe_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( AcquireTracker_6_io_inner_release_ready ),
       .io_inner_release_valid( T10 ),
       .io_inner_release_bits_header_src( io_inner_release_bits_header_src ),
       .io_inner_release_bits_header_dst( io_inner_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( io_inner_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( io_inner_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( io_inner_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( io_inner_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( io_inner_release_bits_payload_r_type ),
       .io_outer_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_outer_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_outer_acquire_bits_header_dst(  )
       .io_outer_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_outer_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_outer_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_outer_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_outer_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_outer_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_outer_finish_valid(  )
       //.io_outer_finish_bits_header_src(  )
       //.io_outer_finish_bits_header_dst(  )
       //.io_outer_finish_bits_payload_master_xact_id(  )
       .io_tile_incoherent( T8 ),
       .io_has_acquire_conflict( AcquireTracker_6_io_has_acquire_conflict )
       //.io_has_release_conflict(  )
  );
  Arbiter_11 alloc_arb(
       .io_in_7_ready( alloc_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_acquire_ready ),
       //.io_in_7_bits(  )
       .io_in_6_ready( alloc_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_acquire_ready ),
       //.io_in_6_bits(  )
       .io_in_5_ready( alloc_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_acquire_ready ),
       //.io_in_5_bits(  )
       .io_in_4_ready( alloc_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_acquire_ready ),
       //.io_in_4_bits(  )
       .io_in_3_ready( alloc_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_acquire_ready ),
       //.io_in_3_bits(  )
       .io_in_2_ready( alloc_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_acquire_ready ),
       //.io_in_2_bits(  )
       .io_in_1_ready( alloc_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_acquire_ready ),
       //.io_in_1_bits(  )
       .io_in_0_ready( alloc_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_acquire_ready ),
       //.io_in_0_bits(  )
       .io_out_ready( T0 )
       //.io_out_valid(  )
       //.io_out_bits(  )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign alloc_arb.io_in_7_bits = {1{$random}};
    assign alloc_arb.io_in_6_bits = {1{$random}};
    assign alloc_arb.io_in_5_bits = {1{$random}};
    assign alloc_arb.io_in_4_bits = {1{$random}};
    assign alloc_arb.io_in_3_bits = {1{$random}};
    assign alloc_arb.io_in_2_bits = {1{$random}};
    assign alloc_arb.io_in_1_bits = {1{$random}};
    assign alloc_arb.io_in_0_bits = {1{$random}};
  `endif
  Arbiter_12 probe_arb(
       .io_in_7_ready( probe_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_probe_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_probe_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_probe_bits_header_dst ),
       .io_in_7_bits_payload_addr( AcquireTracker_6_io_inner_probe_bits_payload_addr ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_p_type( AcquireTracker_6_io_inner_probe_bits_payload_p_type ),
       .io_in_6_ready( probe_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_probe_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_probe_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_probe_bits_header_dst ),
       .io_in_6_bits_payload_addr( AcquireTracker_5_io_inner_probe_bits_payload_addr ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_p_type( AcquireTracker_5_io_inner_probe_bits_payload_p_type ),
       .io_in_5_ready( probe_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_probe_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_probe_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_probe_bits_header_dst ),
       .io_in_5_bits_payload_addr( AcquireTracker_4_io_inner_probe_bits_payload_addr ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_p_type( AcquireTracker_4_io_inner_probe_bits_payload_p_type ),
       .io_in_4_ready( probe_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_probe_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_probe_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_probe_bits_header_dst ),
       .io_in_4_bits_payload_addr( AcquireTracker_3_io_inner_probe_bits_payload_addr ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_p_type( AcquireTracker_3_io_inner_probe_bits_payload_p_type ),
       .io_in_3_ready( probe_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_probe_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_probe_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_probe_bits_header_dst ),
       .io_in_3_bits_payload_addr( AcquireTracker_2_io_inner_probe_bits_payload_addr ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_p_type( AcquireTracker_2_io_inner_probe_bits_payload_p_type ),
       .io_in_2_ready( probe_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_probe_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_probe_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_probe_bits_header_dst ),
       .io_in_2_bits_payload_addr( AcquireTracker_1_io_inner_probe_bits_payload_addr ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_p_type( AcquireTracker_1_io_inner_probe_bits_payload_p_type ),
       .io_in_1_ready( probe_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_probe_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_probe_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_probe_bits_header_dst ),
       .io_in_1_bits_payload_addr( AcquireTracker_0_io_inner_probe_bits_payload_addr ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_probe_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_p_type( AcquireTracker_0_io_inner_probe_bits_payload_p_type ),
       .io_in_0_ready( probe_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_probe_valid ),
       //.io_in_0_bits_header_src(  )
       //.io_in_0_bits_header_dst(  )
       //.io_in_0_bits_payload_addr(  )
       //.io_in_0_bits_payload_master_xact_id(  )
       //.io_in_0_bits_payload_p_type(  )
       .io_out_ready( io_inner_probe_ready ),
       .io_out_valid( probe_arb_io_out_valid ),
       .io_out_bits_header_src( probe_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( probe_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_addr( probe_arb_io_out_bits_payload_addr ),
       .io_out_bits_payload_master_xact_id( probe_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_p_type( probe_arb_io_out_bits_payload_p_type )
       //.io_chosen(  )
  );
  `ifndef SYNTHESIS
    assign probe_arb.io_in_0_bits_header_src = {1{$random}};
    assign probe_arb.io_in_0_bits_header_dst = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_addr = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_master_xact_id = {1{$random}};
    assign probe_arb.io_in_0_bits_payload_p_type = {1{$random}};
  `endif
  Arbiter_13 grant_arb(
       .io_in_7_ready( grant_arb_io_in_7_ready ),
       .io_in_7_valid( AcquireTracker_6_io_inner_grant_valid ),
       .io_in_7_bits_header_src( AcquireTracker_6_io_inner_grant_bits_header_src ),
       .io_in_7_bits_header_dst( AcquireTracker_6_io_inner_grant_bits_header_dst ),
       .io_in_7_bits_payload_data( AcquireTracker_6_io_inner_grant_bits_payload_data ),
       .io_in_7_bits_payload_client_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_7_bits_payload_master_xact_id( AcquireTracker_6_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_7_bits_payload_g_type( AcquireTracker_6_io_inner_grant_bits_payload_g_type ),
       .io_in_6_ready( grant_arb_io_in_6_ready ),
       .io_in_6_valid( AcquireTracker_5_io_inner_grant_valid ),
       .io_in_6_bits_header_src( AcquireTracker_5_io_inner_grant_bits_header_src ),
       .io_in_6_bits_header_dst( AcquireTracker_5_io_inner_grant_bits_header_dst ),
       .io_in_6_bits_payload_data( AcquireTracker_5_io_inner_grant_bits_payload_data ),
       .io_in_6_bits_payload_client_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_6_bits_payload_master_xact_id( AcquireTracker_5_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_6_bits_payload_g_type( AcquireTracker_5_io_inner_grant_bits_payload_g_type ),
       .io_in_5_ready( grant_arb_io_in_5_ready ),
       .io_in_5_valid( AcquireTracker_4_io_inner_grant_valid ),
       .io_in_5_bits_header_src( AcquireTracker_4_io_inner_grant_bits_header_src ),
       .io_in_5_bits_header_dst( AcquireTracker_4_io_inner_grant_bits_header_dst ),
       .io_in_5_bits_payload_data( AcquireTracker_4_io_inner_grant_bits_payload_data ),
       .io_in_5_bits_payload_client_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_5_bits_payload_master_xact_id( AcquireTracker_4_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_5_bits_payload_g_type( AcquireTracker_4_io_inner_grant_bits_payload_g_type ),
       .io_in_4_ready( grant_arb_io_in_4_ready ),
       .io_in_4_valid( AcquireTracker_3_io_inner_grant_valid ),
       .io_in_4_bits_header_src( AcquireTracker_3_io_inner_grant_bits_header_src ),
       .io_in_4_bits_header_dst( AcquireTracker_3_io_inner_grant_bits_header_dst ),
       .io_in_4_bits_payload_data( AcquireTracker_3_io_inner_grant_bits_payload_data ),
       .io_in_4_bits_payload_client_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_4_bits_payload_master_xact_id( AcquireTracker_3_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_4_bits_payload_g_type( AcquireTracker_3_io_inner_grant_bits_payload_g_type ),
       .io_in_3_ready( grant_arb_io_in_3_ready ),
       .io_in_3_valid( AcquireTracker_2_io_inner_grant_valid ),
       .io_in_3_bits_header_src( AcquireTracker_2_io_inner_grant_bits_header_src ),
       .io_in_3_bits_header_dst( AcquireTracker_2_io_inner_grant_bits_header_dst ),
       .io_in_3_bits_payload_data( AcquireTracker_2_io_inner_grant_bits_payload_data ),
       .io_in_3_bits_payload_client_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_3_bits_payload_master_xact_id( AcquireTracker_2_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_3_bits_payload_g_type( AcquireTracker_2_io_inner_grant_bits_payload_g_type ),
       .io_in_2_ready( grant_arb_io_in_2_ready ),
       .io_in_2_valid( AcquireTracker_1_io_inner_grant_valid ),
       .io_in_2_bits_header_src( AcquireTracker_1_io_inner_grant_bits_header_src ),
       .io_in_2_bits_header_dst( AcquireTracker_1_io_inner_grant_bits_header_dst ),
       .io_in_2_bits_payload_data( AcquireTracker_1_io_inner_grant_bits_payload_data ),
       .io_in_2_bits_payload_client_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_2_bits_payload_master_xact_id( AcquireTracker_1_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_2_bits_payload_g_type( AcquireTracker_1_io_inner_grant_bits_payload_g_type ),
       .io_in_1_ready( grant_arb_io_in_1_ready ),
       .io_in_1_valid( AcquireTracker_0_io_inner_grant_valid ),
       .io_in_1_bits_header_src( AcquireTracker_0_io_inner_grant_bits_header_src ),
       .io_in_1_bits_header_dst( AcquireTracker_0_io_inner_grant_bits_header_dst ),
       .io_in_1_bits_payload_data( AcquireTracker_0_io_inner_grant_bits_payload_data ),
       .io_in_1_bits_payload_client_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_1_bits_payload_master_xact_id( AcquireTracker_0_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_1_bits_payload_g_type( AcquireTracker_0_io_inner_grant_bits_payload_g_type ),
       .io_in_0_ready( grant_arb_io_in_0_ready ),
       .io_in_0_valid( VoluntaryReleaseTracker_io_inner_grant_valid ),
       .io_in_0_bits_header_src( VoluntaryReleaseTracker_io_inner_grant_bits_header_src ),
       .io_in_0_bits_header_dst( VoluntaryReleaseTracker_io_inner_grant_bits_header_dst ),
       .io_in_0_bits_payload_data( VoluntaryReleaseTracker_io_inner_grant_bits_payload_data ),
       .io_in_0_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_client_xact_id ),
       .io_in_0_bits_payload_master_xact_id( VoluntaryReleaseTracker_io_inner_grant_bits_payload_master_xact_id ),
       .io_in_0_bits_payload_g_type( VoluntaryReleaseTracker_io_inner_grant_bits_payload_g_type ),
       .io_out_ready( io_inner_grant_ready ),
       .io_out_valid( grant_arb_io_out_valid ),
       .io_out_bits_header_src( grant_arb_io_out_bits_header_src ),
       .io_out_bits_header_dst( grant_arb_io_out_bits_header_dst ),
       .io_out_bits_payload_data( grant_arb_io_out_bits_payload_data ),
       .io_out_bits_payload_client_xact_id( grant_arb_io_out_bits_payload_client_xact_id ),
       .io_out_bits_payload_master_xact_id( grant_arb_io_out_bits_payload_master_xact_id ),
       .io_out_bits_payload_g_type( grant_arb_io_out_bits_payload_g_type )
       //.io_chosen(  )
  );
  UncachedTileLinkIOArbiterThatPassesId outer_arb(.clk(clk), .reset(reset),
       .io_in_7_acquire_ready( outer_arb_io_in_7_acquire_ready ),
       .io_in_7_acquire_valid( AcquireTracker_6_io_outer_acquire_valid ),
       .io_in_7_acquire_bits_header_src( AcquireTracker_6_io_outer_acquire_bits_header_src ),
       //.io_in_7_acquire_bits_header_dst(  )
       .io_in_7_acquire_bits_payload_addr( AcquireTracker_6_io_outer_acquire_bits_payload_addr ),
       .io_in_7_acquire_bits_payload_client_xact_id( AcquireTracker_6_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_7_acquire_bits_payload_data( AcquireTracker_6_io_outer_acquire_bits_payload_data ),
       .io_in_7_acquire_bits_payload_a_type( AcquireTracker_6_io_outer_acquire_bits_payload_a_type ),
       .io_in_7_acquire_bits_payload_write_mask( AcquireTracker_6_io_outer_acquire_bits_payload_write_mask ),
       .io_in_7_acquire_bits_payload_subword_addr( AcquireTracker_6_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_7_acquire_bits_payload_atomic_opcode( AcquireTracker_6_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_7_grant_ready( AcquireTracker_6_io_outer_grant_ready ),
       .io_in_7_grant_valid( outer_arb_io_in_7_grant_valid ),
       .io_in_7_grant_bits_header_src( outer_arb_io_in_7_grant_bits_header_src ),
       .io_in_7_grant_bits_header_dst( outer_arb_io_in_7_grant_bits_header_dst ),
       .io_in_7_grant_bits_payload_data( outer_arb_io_in_7_grant_bits_payload_data ),
       .io_in_7_grant_bits_payload_client_xact_id( outer_arb_io_in_7_grant_bits_payload_client_xact_id ),
       .io_in_7_grant_bits_payload_master_xact_id( outer_arb_io_in_7_grant_bits_payload_master_xact_id ),
       .io_in_7_grant_bits_payload_g_type( outer_arb_io_in_7_grant_bits_payload_g_type ),
       .io_in_7_finish_ready( outer_arb_io_in_7_finish_ready ),
       //.io_in_7_finish_valid(  )
       //.io_in_7_finish_bits_header_src(  )
       //.io_in_7_finish_bits_header_dst(  )
       //.io_in_7_finish_bits_payload_master_xact_id(  )
       .io_in_6_acquire_ready( outer_arb_io_in_6_acquire_ready ),
       .io_in_6_acquire_valid( AcquireTracker_5_io_outer_acquire_valid ),
       .io_in_6_acquire_bits_header_src( AcquireTracker_5_io_outer_acquire_bits_header_src ),
       //.io_in_6_acquire_bits_header_dst(  )
       .io_in_6_acquire_bits_payload_addr( AcquireTracker_5_io_outer_acquire_bits_payload_addr ),
       .io_in_6_acquire_bits_payload_client_xact_id( AcquireTracker_5_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_6_acquire_bits_payload_data( AcquireTracker_5_io_outer_acquire_bits_payload_data ),
       .io_in_6_acquire_bits_payload_a_type( AcquireTracker_5_io_outer_acquire_bits_payload_a_type ),
       .io_in_6_acquire_bits_payload_write_mask( AcquireTracker_5_io_outer_acquire_bits_payload_write_mask ),
       .io_in_6_acquire_bits_payload_subword_addr( AcquireTracker_5_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_6_acquire_bits_payload_atomic_opcode( AcquireTracker_5_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_6_grant_ready( AcquireTracker_5_io_outer_grant_ready ),
       .io_in_6_grant_valid( outer_arb_io_in_6_grant_valid ),
       .io_in_6_grant_bits_header_src( outer_arb_io_in_6_grant_bits_header_src ),
       .io_in_6_grant_bits_header_dst( outer_arb_io_in_6_grant_bits_header_dst ),
       .io_in_6_grant_bits_payload_data( outer_arb_io_in_6_grant_bits_payload_data ),
       .io_in_6_grant_bits_payload_client_xact_id( outer_arb_io_in_6_grant_bits_payload_client_xact_id ),
       .io_in_6_grant_bits_payload_master_xact_id( outer_arb_io_in_6_grant_bits_payload_master_xact_id ),
       .io_in_6_grant_bits_payload_g_type( outer_arb_io_in_6_grant_bits_payload_g_type ),
       .io_in_6_finish_ready( outer_arb_io_in_6_finish_ready ),
       //.io_in_6_finish_valid(  )
       //.io_in_6_finish_bits_header_src(  )
       //.io_in_6_finish_bits_header_dst(  )
       //.io_in_6_finish_bits_payload_master_xact_id(  )
       .io_in_5_acquire_ready( outer_arb_io_in_5_acquire_ready ),
       .io_in_5_acquire_valid( AcquireTracker_4_io_outer_acquire_valid ),
       .io_in_5_acquire_bits_header_src( AcquireTracker_4_io_outer_acquire_bits_header_src ),
       //.io_in_5_acquire_bits_header_dst(  )
       .io_in_5_acquire_bits_payload_addr( AcquireTracker_4_io_outer_acquire_bits_payload_addr ),
       .io_in_5_acquire_bits_payload_client_xact_id( AcquireTracker_4_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_5_acquire_bits_payload_data( AcquireTracker_4_io_outer_acquire_bits_payload_data ),
       .io_in_5_acquire_bits_payload_a_type( AcquireTracker_4_io_outer_acquire_bits_payload_a_type ),
       .io_in_5_acquire_bits_payload_write_mask( AcquireTracker_4_io_outer_acquire_bits_payload_write_mask ),
       .io_in_5_acquire_bits_payload_subword_addr( AcquireTracker_4_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_5_acquire_bits_payload_atomic_opcode( AcquireTracker_4_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_5_grant_ready( AcquireTracker_4_io_outer_grant_ready ),
       .io_in_5_grant_valid( outer_arb_io_in_5_grant_valid ),
       .io_in_5_grant_bits_header_src( outer_arb_io_in_5_grant_bits_header_src ),
       .io_in_5_grant_bits_header_dst( outer_arb_io_in_5_grant_bits_header_dst ),
       .io_in_5_grant_bits_payload_data( outer_arb_io_in_5_grant_bits_payload_data ),
       .io_in_5_grant_bits_payload_client_xact_id( outer_arb_io_in_5_grant_bits_payload_client_xact_id ),
       .io_in_5_grant_bits_payload_master_xact_id( outer_arb_io_in_5_grant_bits_payload_master_xact_id ),
       .io_in_5_grant_bits_payload_g_type( outer_arb_io_in_5_grant_bits_payload_g_type ),
       .io_in_5_finish_ready( outer_arb_io_in_5_finish_ready ),
       //.io_in_5_finish_valid(  )
       //.io_in_5_finish_bits_header_src(  )
       //.io_in_5_finish_bits_header_dst(  )
       //.io_in_5_finish_bits_payload_master_xact_id(  )
       .io_in_4_acquire_ready( outer_arb_io_in_4_acquire_ready ),
       .io_in_4_acquire_valid( AcquireTracker_3_io_outer_acquire_valid ),
       .io_in_4_acquire_bits_header_src( AcquireTracker_3_io_outer_acquire_bits_header_src ),
       //.io_in_4_acquire_bits_header_dst(  )
       .io_in_4_acquire_bits_payload_addr( AcquireTracker_3_io_outer_acquire_bits_payload_addr ),
       .io_in_4_acquire_bits_payload_client_xact_id( AcquireTracker_3_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_4_acquire_bits_payload_data( AcquireTracker_3_io_outer_acquire_bits_payload_data ),
       .io_in_4_acquire_bits_payload_a_type( AcquireTracker_3_io_outer_acquire_bits_payload_a_type ),
       .io_in_4_acquire_bits_payload_write_mask( AcquireTracker_3_io_outer_acquire_bits_payload_write_mask ),
       .io_in_4_acquire_bits_payload_subword_addr( AcquireTracker_3_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_4_acquire_bits_payload_atomic_opcode( AcquireTracker_3_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_4_grant_ready( AcquireTracker_3_io_outer_grant_ready ),
       .io_in_4_grant_valid( outer_arb_io_in_4_grant_valid ),
       .io_in_4_grant_bits_header_src( outer_arb_io_in_4_grant_bits_header_src ),
       .io_in_4_grant_bits_header_dst( outer_arb_io_in_4_grant_bits_header_dst ),
       .io_in_4_grant_bits_payload_data( outer_arb_io_in_4_grant_bits_payload_data ),
       .io_in_4_grant_bits_payload_client_xact_id( outer_arb_io_in_4_grant_bits_payload_client_xact_id ),
       .io_in_4_grant_bits_payload_master_xact_id( outer_arb_io_in_4_grant_bits_payload_master_xact_id ),
       .io_in_4_grant_bits_payload_g_type( outer_arb_io_in_4_grant_bits_payload_g_type ),
       .io_in_4_finish_ready( outer_arb_io_in_4_finish_ready ),
       //.io_in_4_finish_valid(  )
       //.io_in_4_finish_bits_header_src(  )
       //.io_in_4_finish_bits_header_dst(  )
       //.io_in_4_finish_bits_payload_master_xact_id(  )
       .io_in_3_acquire_ready( outer_arb_io_in_3_acquire_ready ),
       .io_in_3_acquire_valid( AcquireTracker_2_io_outer_acquire_valid ),
       .io_in_3_acquire_bits_header_src( AcquireTracker_2_io_outer_acquire_bits_header_src ),
       //.io_in_3_acquire_bits_header_dst(  )
       .io_in_3_acquire_bits_payload_addr( AcquireTracker_2_io_outer_acquire_bits_payload_addr ),
       .io_in_3_acquire_bits_payload_client_xact_id( AcquireTracker_2_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_3_acquire_bits_payload_data( AcquireTracker_2_io_outer_acquire_bits_payload_data ),
       .io_in_3_acquire_bits_payload_a_type( AcquireTracker_2_io_outer_acquire_bits_payload_a_type ),
       .io_in_3_acquire_bits_payload_write_mask( AcquireTracker_2_io_outer_acquire_bits_payload_write_mask ),
       .io_in_3_acquire_bits_payload_subword_addr( AcquireTracker_2_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_3_acquire_bits_payload_atomic_opcode( AcquireTracker_2_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_3_grant_ready( AcquireTracker_2_io_outer_grant_ready ),
       .io_in_3_grant_valid( outer_arb_io_in_3_grant_valid ),
       .io_in_3_grant_bits_header_src( outer_arb_io_in_3_grant_bits_header_src ),
       .io_in_3_grant_bits_header_dst( outer_arb_io_in_3_grant_bits_header_dst ),
       .io_in_3_grant_bits_payload_data( outer_arb_io_in_3_grant_bits_payload_data ),
       .io_in_3_grant_bits_payload_client_xact_id( outer_arb_io_in_3_grant_bits_payload_client_xact_id ),
       .io_in_3_grant_bits_payload_master_xact_id( outer_arb_io_in_3_grant_bits_payload_master_xact_id ),
       .io_in_3_grant_bits_payload_g_type( outer_arb_io_in_3_grant_bits_payload_g_type ),
       .io_in_3_finish_ready( outer_arb_io_in_3_finish_ready ),
       //.io_in_3_finish_valid(  )
       //.io_in_3_finish_bits_header_src(  )
       //.io_in_3_finish_bits_header_dst(  )
       //.io_in_3_finish_bits_payload_master_xact_id(  )
       .io_in_2_acquire_ready( outer_arb_io_in_2_acquire_ready ),
       .io_in_2_acquire_valid( AcquireTracker_1_io_outer_acquire_valid ),
       .io_in_2_acquire_bits_header_src( AcquireTracker_1_io_outer_acquire_bits_header_src ),
       //.io_in_2_acquire_bits_header_dst(  )
       .io_in_2_acquire_bits_payload_addr( AcquireTracker_1_io_outer_acquire_bits_payload_addr ),
       .io_in_2_acquire_bits_payload_client_xact_id( AcquireTracker_1_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_2_acquire_bits_payload_data( AcquireTracker_1_io_outer_acquire_bits_payload_data ),
       .io_in_2_acquire_bits_payload_a_type( AcquireTracker_1_io_outer_acquire_bits_payload_a_type ),
       .io_in_2_acquire_bits_payload_write_mask( AcquireTracker_1_io_outer_acquire_bits_payload_write_mask ),
       .io_in_2_acquire_bits_payload_subword_addr( AcquireTracker_1_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_2_acquire_bits_payload_atomic_opcode( AcquireTracker_1_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_2_grant_ready( AcquireTracker_1_io_outer_grant_ready ),
       .io_in_2_grant_valid( outer_arb_io_in_2_grant_valid ),
       .io_in_2_grant_bits_header_src( outer_arb_io_in_2_grant_bits_header_src ),
       .io_in_2_grant_bits_header_dst( outer_arb_io_in_2_grant_bits_header_dst ),
       .io_in_2_grant_bits_payload_data( outer_arb_io_in_2_grant_bits_payload_data ),
       .io_in_2_grant_bits_payload_client_xact_id( outer_arb_io_in_2_grant_bits_payload_client_xact_id ),
       .io_in_2_grant_bits_payload_master_xact_id( outer_arb_io_in_2_grant_bits_payload_master_xact_id ),
       .io_in_2_grant_bits_payload_g_type( outer_arb_io_in_2_grant_bits_payload_g_type ),
       .io_in_2_finish_ready( outer_arb_io_in_2_finish_ready ),
       //.io_in_2_finish_valid(  )
       //.io_in_2_finish_bits_header_src(  )
       //.io_in_2_finish_bits_header_dst(  )
       //.io_in_2_finish_bits_payload_master_xact_id(  )
       .io_in_1_acquire_ready( outer_arb_io_in_1_acquire_ready ),
       .io_in_1_acquire_valid( AcquireTracker_0_io_outer_acquire_valid ),
       .io_in_1_acquire_bits_header_src( AcquireTracker_0_io_outer_acquire_bits_header_src ),
       //.io_in_1_acquire_bits_header_dst(  )
       .io_in_1_acquire_bits_payload_addr( AcquireTracker_0_io_outer_acquire_bits_payload_addr ),
       .io_in_1_acquire_bits_payload_client_xact_id( AcquireTracker_0_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_1_acquire_bits_payload_data( AcquireTracker_0_io_outer_acquire_bits_payload_data ),
       .io_in_1_acquire_bits_payload_a_type( AcquireTracker_0_io_outer_acquire_bits_payload_a_type ),
       .io_in_1_acquire_bits_payload_write_mask( AcquireTracker_0_io_outer_acquire_bits_payload_write_mask ),
       .io_in_1_acquire_bits_payload_subword_addr( AcquireTracker_0_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_1_acquire_bits_payload_atomic_opcode( AcquireTracker_0_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_1_grant_ready( AcquireTracker_0_io_outer_grant_ready ),
       .io_in_1_grant_valid( outer_arb_io_in_1_grant_valid ),
       .io_in_1_grant_bits_header_src( outer_arb_io_in_1_grant_bits_header_src ),
       .io_in_1_grant_bits_header_dst( outer_arb_io_in_1_grant_bits_header_dst ),
       .io_in_1_grant_bits_payload_data( outer_arb_io_in_1_grant_bits_payload_data ),
       .io_in_1_grant_bits_payload_client_xact_id( outer_arb_io_in_1_grant_bits_payload_client_xact_id ),
       .io_in_1_grant_bits_payload_master_xact_id( outer_arb_io_in_1_grant_bits_payload_master_xact_id ),
       .io_in_1_grant_bits_payload_g_type( outer_arb_io_in_1_grant_bits_payload_g_type ),
       .io_in_1_finish_ready( outer_arb_io_in_1_finish_ready ),
       //.io_in_1_finish_valid(  )
       //.io_in_1_finish_bits_header_src(  )
       //.io_in_1_finish_bits_header_dst(  )
       //.io_in_1_finish_bits_payload_master_xact_id(  )
       .io_in_0_acquire_ready( outer_arb_io_in_0_acquire_ready ),
       .io_in_0_acquire_valid( VoluntaryReleaseTracker_io_outer_acquire_valid ),
       .io_in_0_acquire_bits_header_src( VoluntaryReleaseTracker_io_outer_acquire_bits_header_src ),
       //.io_in_0_acquire_bits_header_dst(  )
       .io_in_0_acquire_bits_payload_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_addr ),
       .io_in_0_acquire_bits_payload_client_xact_id( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_client_xact_id ),
       .io_in_0_acquire_bits_payload_data( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_data ),
       .io_in_0_acquire_bits_payload_a_type( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_a_type ),
       .io_in_0_acquire_bits_payload_write_mask( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_write_mask ),
       .io_in_0_acquire_bits_payload_subword_addr( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_subword_addr ),
       .io_in_0_acquire_bits_payload_atomic_opcode( VoluntaryReleaseTracker_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_in_0_grant_ready( VoluntaryReleaseTracker_io_outer_grant_ready ),
       .io_in_0_grant_valid( outer_arb_io_in_0_grant_valid ),
       .io_in_0_grant_bits_header_src( outer_arb_io_in_0_grant_bits_header_src ),
       .io_in_0_grant_bits_header_dst( outer_arb_io_in_0_grant_bits_header_dst ),
       .io_in_0_grant_bits_payload_data( outer_arb_io_in_0_grant_bits_payload_data ),
       .io_in_0_grant_bits_payload_client_xact_id( outer_arb_io_in_0_grant_bits_payload_client_xact_id ),
       .io_in_0_grant_bits_payload_master_xact_id( outer_arb_io_in_0_grant_bits_payload_master_xact_id ),
       .io_in_0_grant_bits_payload_g_type( outer_arb_io_in_0_grant_bits_payload_g_type ),
       .io_in_0_finish_ready( outer_arb_io_in_0_finish_ready ),
       //.io_in_0_finish_valid(  )
       //.io_in_0_finish_bits_header_src(  )
       //.io_in_0_finish_bits_header_dst(  )
       //.io_in_0_finish_bits_payload_master_xact_id(  )
       .io_out_acquire_ready( io_outer_acquire_ready ),
       .io_out_acquire_valid( outer_arb_io_out_acquire_valid ),
       .io_out_acquire_bits_header_src( outer_arb_io_out_acquire_bits_header_src ),
       .io_out_acquire_bits_header_dst( outer_arb_io_out_acquire_bits_header_dst ),
       .io_out_acquire_bits_payload_addr( outer_arb_io_out_acquire_bits_payload_addr ),
       .io_out_acquire_bits_payload_client_xact_id( outer_arb_io_out_acquire_bits_payload_client_xact_id ),
       .io_out_acquire_bits_payload_data( outer_arb_io_out_acquire_bits_payload_data ),
       .io_out_acquire_bits_payload_a_type( outer_arb_io_out_acquire_bits_payload_a_type ),
       .io_out_acquire_bits_payload_write_mask( outer_arb_io_out_acquire_bits_payload_write_mask ),
       .io_out_acquire_bits_payload_subword_addr( outer_arb_io_out_acquire_bits_payload_subword_addr ),
       .io_out_acquire_bits_payload_atomic_opcode( outer_arb_io_out_acquire_bits_payload_atomic_opcode ),
       .io_out_grant_ready( outer_arb_io_out_grant_ready ),
       .io_out_grant_valid( io_outer_grant_valid ),
       .io_out_grant_bits_header_src( io_outer_grant_bits_header_src ),
       .io_out_grant_bits_header_dst( io_outer_grant_bits_header_dst ),
       .io_out_grant_bits_payload_data( io_outer_grant_bits_payload_data ),
       .io_out_grant_bits_payload_client_xact_id( io_outer_grant_bits_payload_client_xact_id ),
       .io_out_grant_bits_payload_master_xact_id( io_outer_grant_bits_payload_master_xact_id ),
       .io_out_grant_bits_payload_g_type( io_outer_grant_bits_payload_g_type ),
       .io_out_finish_ready( io_outer_finish_ready ),
       .io_out_finish_valid( outer_arb_io_out_finish_valid ),
       .io_out_finish_bits_header_src( outer_arb_io_out_finish_bits_header_src ),
       .io_out_finish_bits_header_dst( outer_arb_io_out_finish_bits_header_dst ),
       .io_out_finish_bits_payload_master_xact_id( outer_arb_io_out_finish_bits_payload_master_xact_id )
  );
  `ifndef SYNTHESIS
    assign outer_arb.io_in_7_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_valid = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_7_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_6_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_valid = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_6_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_5_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_valid = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_5_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_4_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_valid = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_4_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_3_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_valid = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_3_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_2_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_valid = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_2_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_1_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_valid = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_1_finish_bits_payload_master_xact_id = {1{$random}};
    assign outer_arb.io_in_0_acquire_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_valid = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_src = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_header_dst = {1{$random}};
    assign outer_arb.io_in_0_finish_bits_payload_master_xact_id = {1{$random}};
  `endif
endmodule

module Queue_3(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T2;
  wire T3;
  wire T4;
  wire do_deq;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire do_enq;
  wire T9;
  wire ptr_match;
  reg  maybe_full;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire[31:0] T14;
  reg [31:0] ram [1:0];
  wire[31:0] T15;
  wire[31:0] T16;
  wire[31:0] T17;
  wire[5:0] T18;
  wire[4:0] T19;
  wire[25:0] T20;
  wire T21;
  wire empty;
  wire T22;
  wire T23;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T9, ptr_diff};
  assign ptr_diff = R5 - R1;
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = do_deq ? T4 : R1;
  assign T4 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R5;
  assign T8 = R5 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T9 = maybe_full & ptr_match;
  assign ptr_match = R5 == R1;
  assign T10 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign io_deq_bits_rw = T13;
  assign T13 = T14[1'h0:1'h0];
  assign T14 = ram[R1];
  assign T16 = T17;
  assign T17 = {io_enq_bits_addr, T18};
  assign T18 = {io_enq_bits_tag, io_enq_bits_rw};
  assign io_deq_bits_tag = T19;
  assign T19 = T14[3'h5:1'h1];
  assign io_deq_bits_addr = T20;
  assign T20 = T14[5'h1f:3'h6];
  assign io_deq_valid = T21;
  assign T21 = empty ^ 1'h1;
  assign empty = ptr_match & T22;
  assign T22 = maybe_full ^ 1'h1;
  assign io_enq_ready = T23;
  assign T23 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_enq) begin
      R5 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R5] <= T16;
  end
endmodule

module Queue_4(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[1:0] io_count
);

  wire[1:0] T0;
  wire ptr_diff;
  reg  R1;
  wire T2;
  wire T3;
  wire T4;
  wire do_deq;
  reg  R5;
  wire T6;
  wire T7;
  wire T8;
  wire do_enq;
  wire T9;
  wire ptr_match;
  reg  maybe_full;
  wire T10;
  wire T11;
  wire T12;
  wire[127:0] T13;
  wire[127:0] T14;
  reg [127:0] ram [1:0];
  wire[127:0] T15;
  wire T16;
  wire empty;
  wire T17;
  wire T18;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{$random}};
    R5 = {1{$random}};
    maybe_full = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {4{$random}};
  end
`endif

  assign io_count = T0;
  assign T0 = {T9, ptr_diff};
  assign ptr_diff = R5 - R1;
  assign T2 = reset ? 1'h0 : T3;
  assign T3 = do_deq ? T4 : R1;
  assign T4 = R1 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T6 = reset ? 1'h0 : T7;
  assign T7 = do_enq ? T8 : R5;
  assign T8 = R5 + 1'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T9 = maybe_full & ptr_match;
  assign ptr_match = R5 == R1;
  assign T10 = reset ? 1'h0 : T11;
  assign T11 = T12 ? do_enq : maybe_full;
  assign T12 = do_enq != do_deq;
  assign io_deq_bits_data = T13;
  assign T13 = T14[7'h7f:1'h0];
  assign T14 = ram[R1];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign io_enq_ready = T18;
  assign T18 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else if(do_deq) begin
      R1 <= T4;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else if(do_enq) begin
      R5 <= T8;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T12) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R5] <= io_enq_bits_data;
  end
endmodule

module MemIOUncachedTileLinkIOConverter(input clk, input reset,
    output io_uncached_acquire_ready,
    input  io_uncached_acquire_valid,
    input [1:0] io_uncached_acquire_bits_header_src,
    input [1:0] io_uncached_acquire_bits_header_dst,
    input [25:0] io_uncached_acquire_bits_payload_addr,
    input [1:0] io_uncached_acquire_bits_payload_client_xact_id,
    input [511:0] io_uncached_acquire_bits_payload_data,
    input [2:0] io_uncached_acquire_bits_payload_a_type,
    input [5:0] io_uncached_acquire_bits_payload_write_mask,
    input [2:0] io_uncached_acquire_bits_payload_subword_addr,
    input [3:0] io_uncached_acquire_bits_payload_atomic_opcode,
    input  io_uncached_grant_ready,
    output io_uncached_grant_valid,
    //output[1:0] io_uncached_grant_bits_header_src
    //output[1:0] io_uncached_grant_bits_header_dst
    output[511:0] io_uncached_grant_bits_payload_data,
    output[1:0] io_uncached_grant_bits_payload_client_xact_id,
    output[2:0] io_uncached_grant_bits_payload_master_xact_id,
    output[3:0] io_uncached_grant_bits_payload_g_type,
    //output io_uncached_finish_ready
    input  io_uncached_finish_valid,
    input [1:0] io_uncached_finish_bits_header_src,
    input [1:0] io_uncached_finish_bits_header_dst,
    input [2:0] io_uncached_finish_bits_payload_master_xact_id,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire[127:0] T0;
  reg [511:0] buf_out;
  wire[511:0] T1;
  wire[511:0] T2;
  wire T3;
  wire T4;
  reg  active_out;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  reg [2:0] cnt_out;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire T15;
  wire T16;
  wire mem_data_q_io_enq_ready;
  wire T17;
  reg  has_data;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  reg  cmd_sent_out;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire mem_cmd_q_io_enq_ready;
  wire[511:0] T30;
  wire[383:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire[4:0] T35;
  reg [1:0] tag_out;
  wire[1:0] T36;
  reg [25:0] addr_out;
  wire[25:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg [2:0] cnt_in;
  wire[2:0] T42;
  wire[2:0] T43;
  wire T44;
  wire T45;
  reg  active_in;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire[2:0] T51;
  wire T52;
  wire T53;
  wire T54;
  wire[127:0] mem_data_q_io_deq_bits_data;
  wire mem_data_q_io_deq_valid;
  wire mem_cmd_q_io_deq_bits_rw;
  wire[4:0] mem_cmd_q_io_deq_bits_tag;
  wire[25:0] mem_cmd_q_io_deq_bits_addr;
  wire mem_cmd_q_io_deq_valid;
  wire[3:0] T55;
  wire[2:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  reg [4:0] tag_in;
  wire[4:0] T59;
  wire[511:0] T60;
  reg [511:0] buf_in;
  wire[511:0] T61;
  wire[511:0] T62;
  wire[511:0] T63;
  wire[511:0] T64;
  wire[383:0] T65;
  wire T66;
  wire T67;
  wire T68;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    buf_out = {16{$random}};
    active_out = {1{$random}};
    cnt_out = {1{$random}};
    has_data = {1{$random}};
    cmd_sent_out = {1{$random}};
    tag_out = {1{$random}};
    addr_out = {1{$random}};
    cnt_in = {1{$random}};
    active_in = {1{$random}};
    tag_in = {1{$random}};
    buf_in = {16{$random}};
  end
`endif

  assign T0 = buf_out[7'h7f:1'h0];
  assign T1 = T15 ? T30 : T2;
  assign T2 = T3 ? io_uncached_acquire_bits_payload_data : buf_out;
  assign T3 = T4 & io_uncached_acquire_valid;
  assign T4 = active_out ^ 1'h1;
  assign T5 = reset ? 1'h0 : T6;
  assign T6 = T8 ? 1'h0 : T7;
  assign T7 = T3 ? 1'h1 : active_out;
  assign T8 = active_out & T9;
  assign T9 = cmd_sent_out & T10;
  assign T10 = T17 | T11;
  assign T11 = cnt_out == 3'h4;
  assign T12 = T15 ? T14 : T13;
  assign T13 = T3 ? 3'h0 : cnt_out;
  assign T14 = cnt_out + 3'h1;
  assign T15 = active_out & T16;
  assign T16 = mem_data_q_io_enq_ready & T32;
  assign T17 = has_data ^ 1'h1;
  assign T18 = reset ? 1'h0 : T19;
  assign T19 = T3 ? T20 : has_data;
  assign T20 = T22 | T21;
  assign T21 = 3'h6 == io_uncached_acquire_bits_payload_a_type;
  assign T22 = T24 | T23;
  assign T23 = 3'h5 == io_uncached_acquire_bits_payload_a_type;
  assign T24 = 3'h3 == io_uncached_acquire_bits_payload_a_type;
  assign T25 = reset ? 1'h0 : T26;
  assign T26 = T28 ? 1'h1 : T27;
  assign T27 = T3 ? 1'h0 : cmd_sent_out;
  assign T28 = active_out & T29;
  assign T29 = mem_cmd_q_io_enq_ready & T38;
  assign T30 = {128'h0, T31};
  assign T31 = buf_out >> 8'h80;
  assign T32 = T34 & T33;
  assign T33 = cnt_out < 3'h4;
  assign T34 = active_out & has_data;
  assign T35 = {3'h0, tag_out};
  assign T36 = T3 ? io_uncached_acquire_bits_payload_client_xact_id : tag_out;
  assign T37 = T3 ? io_uncached_acquire_bits_payload_addr : addr_out;
  assign T38 = active_out & T39;
  assign T39 = cmd_sent_out ^ 1'h1;
  assign io_mem_resp_ready = T40;
  assign T40 = T54 | T41;
  assign T41 = cnt_in < 3'h4;
  assign T42 = T52 ? T51 : T43;
  assign T43 = T44 ? 3'h1 : cnt_in;
  assign T44 = T45 & io_mem_resp_valid;
  assign T45 = active_in ^ 1'h1;
  assign T46 = reset ? 1'h0 : T47;
  assign T47 = T49 ? 1'h0 : T48;
  assign T48 = T44 ? 1'h1 : active_in;
  assign T49 = active_in & T50;
  assign T50 = io_uncached_grant_ready & io_uncached_grant_valid;
  assign T51 = cnt_in + 3'h1;
  assign T52 = active_in & T53;
  assign T53 = io_mem_resp_ready & io_mem_resp_valid;
  assign T54 = active_in ^ 1'h1;
  assign io_mem_req_data_bits_data = mem_data_q_io_deq_bits_data;
  assign io_mem_req_data_valid = mem_data_q_io_deq_valid;
  assign io_mem_req_cmd_bits_rw = mem_cmd_q_io_deq_bits_rw;
  assign io_mem_req_cmd_bits_tag = mem_cmd_q_io_deq_bits_tag;
  assign io_mem_req_cmd_bits_addr = mem_cmd_q_io_deq_bits_addr;
  assign io_mem_req_cmd_valid = mem_cmd_q_io_deq_valid;
  assign io_uncached_grant_bits_payload_g_type = T55;
  assign T55 = 4'h0;
  assign io_uncached_grant_bits_payload_master_xact_id = T56;
  assign T56 = 3'h0;
  assign io_uncached_grant_bits_payload_client_xact_id = T57;
  assign T57 = T58;
  assign T58 = tag_in[1'h1:1'h0];
  assign T59 = T44 ? io_mem_resp_bits_tag : tag_in;
  assign io_uncached_grant_bits_payload_data = T60;
  assign T60 = buf_in;
  assign T61 = T52 ? T64 : T62;
  assign T62 = T44 ? T63 : buf_in;
  assign T63 = io_mem_resp_bits_data << 9'h180;
  assign T64 = {io_mem_resp_bits_data, T65};
  assign T65 = buf_in[9'h1ff:8'h80];
  assign io_uncached_grant_valid = T66;
  assign T66 = active_in & T67;
  assign T67 = cnt_in == 3'h4;
  assign io_uncached_acquire_ready = T68;
  assign T68 = active_out ^ 1'h1;
  Queue_3 mem_cmd_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_cmd_q_io_enq_ready ),
       .io_enq_valid( T38 ),
       .io_enq_bits_addr( addr_out ),
       .io_enq_bits_tag( T35 ),
       .io_enq_bits_rw( has_data ),
       .io_deq_ready( io_mem_req_cmd_ready ),
       .io_deq_valid( mem_cmd_q_io_deq_valid ),
       .io_deq_bits_addr( mem_cmd_q_io_deq_bits_addr ),
       .io_deq_bits_tag( mem_cmd_q_io_deq_bits_tag ),
       .io_deq_bits_rw( mem_cmd_q_io_deq_bits_rw )
       //.io_count(  )
  );
  Queue_4 mem_data_q(.clk(clk), .reset(reset),
       .io_enq_ready( mem_data_q_io_enq_ready ),
       .io_enq_valid( T32 ),
       .io_enq_bits_data( T0 ),
       .io_deq_ready( io_mem_req_data_ready ),
       .io_deq_valid( mem_data_q_io_deq_valid ),
       .io_deq_bits_data( mem_data_q_io_deq_bits_data )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(T15) begin
      buf_out <= T30;
    end else if(T3) begin
      buf_out <= io_uncached_acquire_bits_payload_data;
    end
    if(reset) begin
      active_out <= 1'h0;
    end else if(T8) begin
      active_out <= 1'h0;
    end else if(T3) begin
      active_out <= 1'h1;
    end
    if(T15) begin
      cnt_out <= T14;
    end else if(T3) begin
      cnt_out <= 3'h0;
    end
    if(reset) begin
      has_data <= 1'h0;
    end else if(T3) begin
      has_data <= T20;
    end
    if(reset) begin
      cmd_sent_out <= 1'h0;
    end else if(T28) begin
      cmd_sent_out <= 1'h1;
    end else if(T3) begin
      cmd_sent_out <= 1'h0;
    end
    if(T3) begin
      tag_out <= io_uncached_acquire_bits_payload_client_xact_id;
    end
    if(T3) begin
      addr_out <= io_uncached_acquire_bits_payload_addr;
    end
    if(T52) begin
      cnt_in <= T51;
    end else if(T44) begin
      cnt_in <= 3'h1;
    end
    if(reset) begin
      active_in <= 1'h0;
    end else if(T49) begin
      active_in <= 1'h0;
    end else if(T44) begin
      active_in <= 1'h1;
    end
    if(T44) begin
      tag_in <= io_mem_resp_bits_tag;
    end
    if(T52) begin
      buf_in <= T64;
    end else if(T44) begin
      buf_in <= T63;
    end
  end
endmodule

module HellaFlowQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[5:0] io_count
);

  wire[4:0] T0;
  wire[4:0] T1;
  wire[132:0] T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire empty;
  wire T7;
  reg  maybe_full;
  wire T8;
  wire T9;
  wire do_enq;
  wire T10;
  wire do_flow;
  wire T11;
  wire T12;
  wire T13;
  wire do_deq;
  wire T14;
  wire T15;
  wire ptr_match;
  reg [4:0] deq_ptr;
  wire[4:0] T16;
  wire[4:0] T17;
  wire[4:0] T18;
  reg [4:0] enq_ptr;
  wire[4:0] T19;
  wire[4:0] T20;
  wire[4:0] T21;
  wire T22;
  wire atLeastTwo;
  wire T23;
  wire[4:0] T24;
  wire full;
  wire[4:0] T25;
  wire[4:0] T26;
  wire[132:0] T27;
  wire[132:0] T28;
  wire[132:0] T29;
  reg [4:0] ram_addr;
  wire[4:0] T30;
  wire[127:0] T31;
  wire[127:0] T32;
  wire T33;
  reg  ram_out_valid;
  wire T34;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    maybe_full = {1{$random}};
    deq_ptr = {1{$random}};
    enq_ptr = {1{$random}};
    ram_addr = {1{$random}};
    ram_out_valid = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = empty ? io_enq_bits_tag : T1;
  assign T1 = T2[3'h4:1'h0];
  assign T3 = io_deq_ready & T4;
  assign T4 = atLeastTwo | T5;
  assign T5 = T22 & T6;
  assign T6 = empty ^ 1'h1;
  assign empty = ptr_match & T7;
  assign T7 = maybe_full ^ 1'h1;
  assign T8 = reset ? 1'h0 : T9;
  assign T9 = T13 ? do_enq : maybe_full;
  assign do_enq = T12 & T10;
  assign T10 = do_flow ^ 1'h1;
  assign do_flow = T11;
  assign T11 = empty & io_deq_ready;
  assign T12 = io_enq_ready & io_enq_valid;
  assign T13 = do_enq != do_deq;
  assign do_deq = T15 & T14;
  assign T14 = do_flow ^ 1'h1;
  assign T15 = io_deq_ready & io_deq_valid;
  assign ptr_match = enq_ptr == deq_ptr;
  assign T16 = reset ? 5'h0 : T17;
  assign T17 = do_deq ? T18 : deq_ptr;
  assign T18 = deq_ptr + 5'h1;
  assign T19 = reset ? 5'h0 : T20;
  assign T20 = do_enq ? T21 : enq_ptr;
  assign T21 = enq_ptr + 5'h1;
  assign T22 = io_deq_valid ^ 1'h1;
  assign atLeastTwo = full | T23;
  assign T23 = 5'h2 <= T24;
  assign T24 = enq_ptr - deq_ptr;
  assign full = ptr_match & maybe_full;
  assign T25 = io_deq_valid ? T26 : deq_ptr;
  assign T26 = deq_ptr + 5'h1;
  HellaFlowQueue_ram ram (
    .CLK(clk),
    .W0A(enq_ptr),
    .W0E(do_enq),
    .W0I(T28),
    .R1A(T25),
    .R1E(T3),
    .R1O(T2)
  );
  assign T28 = T29;
  assign T29 = {io_enq_bits_data, io_enq_bits_tag};
  assign T30 = T3 ? T25 : ram_addr;
  assign io_deq_bits_data = T31;
  assign T31 = empty ? io_enq_bits_data : T32;
  assign T32 = T2[8'h84:3'h5];
  assign io_deq_valid = T33;
  assign T33 = empty ? io_enq_valid : ram_out_valid;
  assign io_enq_ready = T34;
  assign T34 = full ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T13) begin
      maybe_full <= do_enq;
    end
    if(reset) begin
      deq_ptr <= 5'h0;
    end else if(do_deq) begin
      deq_ptr <= T18;
    end
    if(reset) begin
      enq_ptr <= 5'h0;
    end else if(do_enq) begin
      enq_ptr <= T21;
    end
    if(T3) begin
      ram_addr <= T25;
    end
    ram_out_valid <= T3;
  end
endmodule

module Queue_5(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
);

  wire[4:0] T0;
  wire[132:0] T1;
  reg [132:0] ram [0:0];
  wire[132:0] T2;
  wire[132:0] T3;
  wire[132:0] T4;
  wire do_enq;
  wire[127:0] T5;
  wire T6;
  wire empty;
  reg  maybe_full;
  wire T7;
  wire T8;
  wire T9;
  wire do_deq;
  wire T10;
  wire T11;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {5{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_tag = T0;
  assign T0 = T1[3'h4:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {io_enq_bits_data, io_enq_bits_tag};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_data = T5;
  assign T5 = T1[8'h84:3'h5];
  assign io_deq_valid = T6;
  assign T6 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T10;
  assign T10 = T11 | io_deq_ready;
  assign T11 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module HellaQueue(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input [4:0] io_enq_bits_tag,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data,
    output[4:0] io_deq_bits_tag
    //output[5:0] io_count
);

  wire[4:0] fq_io_deq_bits_tag;
  wire[127:0] fq_io_deq_bits_data;
  wire fq_io_deq_valid;
  wire Queue_io_enq_ready;
  wire[4:0] Queue_io_deq_bits_tag;
  wire[127:0] Queue_io_deq_bits_data;
  wire Queue_io_deq_valid;
  wire fq_io_enq_ready;


  assign io_deq_bits_tag = Queue_io_deq_bits_tag;
  assign io_deq_bits_data = Queue_io_deq_bits_data;
  assign io_deq_valid = Queue_io_deq_valid;
  assign io_enq_ready = fq_io_enq_ready;
  HellaFlowQueue fq(.clk(clk), .reset(reset),
       .io_enq_ready( fq_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_data( io_enq_bits_data ),
       .io_enq_bits_tag( io_enq_bits_tag ),
       .io_deq_ready( Queue_io_enq_ready ),
       .io_deq_valid( fq_io_deq_valid ),
       .io_deq_bits_data( fq_io_deq_bits_data ),
       .io_deq_bits_tag( fq_io_deq_bits_tag )
       //.io_count(  )
  );
  Queue_5 Queue(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_io_enq_ready ),
       .io_enq_valid( fq_io_deq_valid ),
       .io_enq_bits_data( fq_io_deq_bits_data ),
       .io_enq_bits_tag( fq_io_deq_bits_tag ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( Queue_io_deq_valid ),
       .io_deq_bits_data( Queue_io_deq_bits_data ),
       .io_deq_bits_tag( Queue_io_deq_bits_tag )
  );
endmodule

module DRAMSideLLCNull(input clk, input reset,
    output io_cpu_req_cmd_ready,
    input  io_cpu_req_cmd_valid,
    input [25:0] io_cpu_req_cmd_bits_addr,
    input [4:0] io_cpu_req_cmd_bits_tag,
    input  io_cpu_req_cmd_bits_rw,
    output io_cpu_req_data_ready,
    input  io_cpu_req_data_valid,
    input [127:0] io_cpu_req_data_bits_data,
    input  io_cpu_resp_ready,
    output io_cpu_resp_valid,
    output[127:0] io_cpu_resp_bits_data,
    output[4:0] io_cpu_resp_bits_tag,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
);

  wire T0;
  wire cmdq_mask;
  wire T1;
  reg [5:0] count;
  wire[5:0] T2;
  wire[5:0] T3;
  wire[5:0] T4;
  wire[5:0] T5;
  wire[5:0] T6;
  wire T7;
  wire T8;
  wire dec;
  wire T9;
  wire T10;
  wire T11;
  wire inc;
  wire T12;
  wire resp_dataq_io_deq_valid;
  wire[5:0] T13;
  wire T14;
  wire T15;
  wire[5:0] T16;
  wire T17;
  wire[4:0] resp_dataq_io_deq_bits_tag;
  wire[127:0] resp_dataq_io_deq_bits_data;
  wire T18;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    count = {1{$random}};
  end
`endif

  assign io_mem_req_data_bits_data = io_cpu_req_data_bits_data;
  assign io_mem_req_data_valid = io_cpu_req_data_valid;
  assign io_mem_req_cmd_bits_rw = io_cpu_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = io_cpu_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = io_cpu_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = T0;
  assign T0 = io_cpu_req_cmd_valid & cmdq_mask;
  assign cmdq_mask = io_cpu_req_cmd_bits_rw | T1;
  assign T1 = 6'h4 <= count;
  assign T2 = reset ? 6'h20 : T3;
  assign T3 = T17 ? T16 : T4;
  assign T4 = T14 ? T13 : T5;
  assign T5 = T7 ? T6 : count;
  assign T6 = count + 6'h1;
  assign T7 = inc & T8;
  assign T8 = dec ^ 1'h1;
  assign dec = T9;
  assign T9 = T11 & T10;
  assign T10 = io_mem_req_cmd_bits_rw ^ 1'h1;
  assign T11 = io_mem_req_cmd_ready & io_mem_req_cmd_valid;
  assign inc = T12;
  assign T12 = io_cpu_resp_ready & resp_dataq_io_deq_valid;
  assign T13 = count - 6'h4;
  assign T14 = T15 & dec;
  assign T15 = inc ^ 1'h1;
  assign T16 = count - 6'h3;
  assign T17 = inc & dec;
  assign io_cpu_resp_bits_tag = resp_dataq_io_deq_bits_tag;
  assign io_cpu_resp_bits_data = resp_dataq_io_deq_bits_data;
  assign io_cpu_resp_valid = resp_dataq_io_deq_valid;
  assign io_cpu_req_data_ready = io_mem_req_data_ready;
  assign io_cpu_req_cmd_ready = T18;
  assign T18 = io_mem_req_cmd_ready & cmdq_mask;
  HellaQueue resp_dataq(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_mem_resp_valid ),
       .io_enq_bits_data( io_mem_resp_bits_data ),
       .io_enq_bits_tag( io_mem_resp_bits_tag ),
       .io_deq_ready( io_cpu_resp_ready ),
       .io_deq_valid( resp_dataq_io_deq_valid ),
       .io_deq_bits_data( resp_dataq_io_deq_bits_data ),
       .io_deq_bits_tag( resp_dataq_io_deq_bits_tag )
       //.io_count(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      count <= 6'h20;
    end else if(T17) begin
      count <= T16;
    end else if(T14) begin
      count <= T13;
    end else if(T7) begin
      count <= T6;
    end
  end
endmodule

module Queue_6(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [25:0] io_enq_bits_addr,
    input [4:0] io_enq_bits_tag,
    input  io_enq_bits_rw,
    input  io_deq_ready,
    output io_deq_valid,
    output[25:0] io_deq_bits_addr,
    output[4:0] io_deq_bits_tag,
    output io_deq_bits_rw
);

  wire T0;
  wire[31:0] T1;
  reg [31:0] ram [1:0];
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[5:0] T5;
  wire do_enq;
  reg  R6;
  wire T7;
  wire T8;
  wire T9;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  wire do_deq;
  wire[4:0] T14;
  wire[25:0] T15;
  wire T16;
  wire empty;
  wire T17;
  reg  maybe_full;
  wire T18;
  wire T19;
  wire T20;
  wire ptr_match;
  wire T21;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R10 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_rw = T0;
  assign T0 = T1[1'h0:1'h0];
  assign T1 = ram[R10];
  assign T3 = T4;
  assign T4 = {io_enq_bits_addr, T5};
  assign T5 = {io_enq_bits_tag, io_enq_bits_rw};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_enq ? T9 : R6;
  assign T9 = R6 + 1'h1;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_deq ? T13 : R10;
  assign T13 = R10 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_tag = T14;
  assign T14 = T1[3'h5:1'h1];
  assign io_deq_bits_addr = T15;
  assign T15 = T1[5'h1f:3'h6];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign T18 = reset ? 1'h0 : T19;
  assign T19 = T20 ? do_enq : maybe_full;
  assign T20 = do_enq != do_deq;
  assign ptr_match = R6 == R10;
  assign io_enq_ready = T21;
  assign T21 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T9;
    end
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_deq) begin
      R10 <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T20) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_7(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [127:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output[127:0] io_deq_bits_data
);

  wire[127:0] T0;
  wire[127:0] T1;
  reg [127:0] ram [3:0];
  wire[127:0] T2;
  wire do_enq;
  reg [1:0] R3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  reg [1:0] R7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire do_deq;
  wire T11;
  wire empty;
  wire T12;
  reg  maybe_full;
  wire T13;
  wire T14;
  wire T15;
  wire ptr_match;
  wire T16;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      ram[initvar] = {4{$random}};
    R3 = {1{$random}};
    R7 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[7'h7f:1'h0];
  assign T1 = ram[R7];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T4 = reset ? 2'h0 : T5;
  assign T5 = do_enq ? T6 : R3;
  assign T6 = R3 + 2'h1;
  assign T8 = reset ? 2'h0 : T9;
  assign T9 = do_deq ? T10 : R7;
  assign T10 = R7 + 2'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T11;
  assign T11 = empty ^ 1'h1;
  assign empty = ptr_match & T12;
  assign T12 = maybe_full ^ 1'h1;
  assign T13 = reset ? 1'h0 : T14;
  assign T14 = T15 ? do_enq : maybe_full;
  assign T15 = do_enq != do_deq;
  assign ptr_match = R3 == R7;
  assign io_enq_ready = T16;
  assign T16 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R3] <= io_enq_bits_data;
    if(reset) begin
      R3 <= 2'h0;
    end else if(do_enq) begin
      R3 <= T6;
    end
    if(reset) begin
      R7 <= 2'h0;
    end else if(do_deq) begin
      R7 <= T10;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T15) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module OuterMemorySystem(input clk, input reset,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_acquire_ready,
    input  io_htif_acquire_valid,
    input [1:0] io_htif_acquire_bits_header_src,
    input [1:0] io_htif_acquire_bits_header_dst,
    input [25:0] io_htif_acquire_bits_payload_addr,
    input [1:0] io_htif_acquire_bits_payload_client_xact_id,
    input [511:0] io_htif_acquire_bits_payload_data,
    input [2:0] io_htif_acquire_bits_payload_a_type,
    input [5:0] io_htif_acquire_bits_payload_write_mask,
    input [2:0] io_htif_acquire_bits_payload_subword_addr,
    input [3:0] io_htif_acquire_bits_payload_atomic_opcode,
    input  io_htif_grant_ready,
    output io_htif_grant_valid,
    output[1:0] io_htif_grant_bits_header_src,
    output[1:0] io_htif_grant_bits_header_dst,
    output[511:0] io_htif_grant_bits_payload_data,
    output[1:0] io_htif_grant_bits_payload_client_xact_id,
    output[2:0] io_htif_grant_bits_payload_master_xact_id,
    output[3:0] io_htif_grant_bits_payload_g_type,
    output io_htif_finish_ready,
    input  io_htif_finish_valid,
    input [1:0] io_htif_finish_bits_header_src,
    input [1:0] io_htif_finish_bits_header_dst,
    input [2:0] io_htif_finish_bits_payload_master_xact_id,
    input  io_htif_probe_ready,
    output io_htif_probe_valid,
    output[1:0] io_htif_probe_bits_header_src,
    output[1:0] io_htif_probe_bits_header_dst,
    output[25:0] io_htif_probe_bits_payload_addr,
    output[2:0] io_htif_probe_bits_payload_master_xact_id,
    output[1:0] io_htif_probe_bits_payload_p_type,
    output io_htif_release_ready,
    input  io_htif_release_valid,
    input [1:0] io_htif_release_bits_header_src,
    input [1:0] io_htif_release_bits_header_dst,
    input [25:0] io_htif_release_bits_payload_addr,
    input [1:0] io_htif_release_bits_payload_client_xact_id,
    input [2:0] io_htif_release_bits_payload_master_xact_id,
    input [511:0] io_htif_release_bits_payload_data,
    input [2:0] io_htif_release_bits_payload_r_type,
    input  io_incoherent_1,
    input  io_incoherent_0,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire llc_io_cpu_req_data_ready;
  wire[127:0] conv_io_mem_req_data_bits_data;
  wire conv_io_mem_req_data_valid;
  wire llc_io_cpu_req_cmd_ready;
  wire conv_io_mem_req_cmd_bits_rw;
  wire[4:0] conv_io_mem_req_cmd_bits_tag;
  wire[25:0] conv_io_mem_req_cmd_bits_addr;
  wire conv_io_mem_req_cmd_valid;
  wire conv_io_mem_resp_ready;
  wire[127:0] Queue_1_io_deq_bits_data;
  wire Queue_1_io_deq_valid;
  wire Queue_0_io_deq_bits_rw;
  wire[4:0] Queue_0_io_deq_bits_tag;
  wire[25:0] Queue_0_io_deq_bits_addr;
  wire Queue_0_io_deq_valid;
  wire[4:0] llc_io_cpu_resp_bits_tag;
  wire[127:0] llc_io_cpu_resp_bits_data;
  wire llc_io_cpu_resp_valid;
  wire Queue_1_io_enq_ready;
  wire Queue_0_io_enq_ready;
  wire[2:0] L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_dst;
  wire[1:0] L2CoherenceAgent_io_outer_finish_bits_header_src;
  wire L2CoherenceAgent_io_outer_finish_valid;
  wire L2CoherenceAgent_io_outer_grant_ready;
  wire[3:0] L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr;
  wire[5:0] L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask;
  wire[2:0] L2CoherenceAgent_io_outer_acquire_bits_payload_a_type;
  wire[511:0] L2CoherenceAgent_io_outer_acquire_bits_payload_data;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id;
  wire[25:0] L2CoherenceAgent_io_outer_acquire_bits_payload_addr;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_dst;
  wire[1:0] L2CoherenceAgent_io_outer_acquire_bits_header_src;
  wire L2CoherenceAgent_io_outer_acquire_valid;
  wire[3:0] conv_io_uncached_grant_bits_payload_g_type;
  wire[2:0] conv_io_uncached_grant_bits_payload_master_xact_id;
  wire[1:0] conv_io_uncached_grant_bits_payload_client_xact_id;
  wire[511:0] conv_io_uncached_grant_bits_payload_data;
  wire conv_io_uncached_grant_valid;
  wire conv_io_uncached_acquire_ready;
  wire[2:0] net_io_masters_0_release_bits_payload_r_type;
  wire[511:0] net_io_masters_0_release_bits_payload_data;
  wire[2:0] net_io_masters_0_release_bits_payload_master_xact_id;
  wire[1:0] net_io_masters_0_release_bits_payload_client_xact_id;
  wire[25:0] net_io_masters_0_release_bits_payload_addr;
  wire[1:0] net_io_masters_0_release_bits_header_dst;
  wire[1:0] net_io_masters_0_release_bits_header_src;
  wire net_io_masters_0_release_valid;
  wire net_io_masters_0_probe_ready;
  wire[2:0] net_io_masters_0_finish_bits_payload_master_xact_id;
  wire[1:0] net_io_masters_0_finish_bits_header_dst;
  wire[1:0] net_io_masters_0_finish_bits_header_src;
  wire net_io_masters_0_finish_valid;
  wire net_io_masters_0_grant_ready;
  wire[3:0] net_io_masters_0_acquire_bits_payload_atomic_opcode;
  wire[2:0] net_io_masters_0_acquire_bits_payload_subword_addr;
  wire[5:0] net_io_masters_0_acquire_bits_payload_write_mask;
  wire[2:0] net_io_masters_0_acquire_bits_payload_a_type;
  wire[511:0] net_io_masters_0_acquire_bits_payload_data;
  wire[1:0] net_io_masters_0_acquire_bits_payload_client_xact_id;
  wire[25:0] net_io_masters_0_acquire_bits_payload_addr;
  wire[1:0] net_io_masters_0_acquire_bits_header_dst;
  wire[1:0] net_io_masters_0_acquire_bits_header_src;
  wire net_io_masters_0_acquire_valid;
  wire L2CoherenceAgent_io_inner_release_ready;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_payload_p_type;
  wire[2:0] L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id;
  wire[25:0] L2CoherenceAgent_io_inner_probe_bits_payload_addr;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_dst;
  wire[1:0] L2CoherenceAgent_io_inner_probe_bits_header_src;
  wire L2CoherenceAgent_io_inner_probe_valid;
  wire L2CoherenceAgent_io_inner_finish_ready;
  wire[3:0] L2CoherenceAgent_io_inner_grant_bits_payload_g_type;
  wire[2:0] L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id;
  wire[511:0] L2CoherenceAgent_io_inner_grant_bits_payload_data;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_dst;
  wire[1:0] L2CoherenceAgent_io_inner_grant_bits_header_src;
  wire L2CoherenceAgent_io_inner_grant_valid;
  wire L2CoherenceAgent_io_inner_acquire_ready;
  wire[127:0] llc_io_mem_req_data_bits_data;
  wire llc_io_mem_req_data_valid;
  wire llc_io_mem_req_cmd_bits_rw;
  wire[4:0] llc_io_mem_req_cmd_bits_tag;
  wire[25:0] llc_io_mem_req_cmd_bits_addr;
  wire llc_io_mem_req_cmd_valid;
  wire net_io_clients_1_release_ready;
  wire[1:0] net_io_clients_1_probe_bits_payload_p_type;
  wire[2:0] net_io_clients_1_probe_bits_payload_master_xact_id;
  wire[25:0] net_io_clients_1_probe_bits_payload_addr;
  wire[1:0] net_io_clients_1_probe_bits_header_dst;
  wire[1:0] net_io_clients_1_probe_bits_header_src;
  wire net_io_clients_1_probe_valid;
  wire net_io_clients_1_finish_ready;
  wire[3:0] net_io_clients_1_grant_bits_payload_g_type;
  wire[2:0] net_io_clients_1_grant_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_1_grant_bits_payload_client_xact_id;
  wire[511:0] net_io_clients_1_grant_bits_payload_data;
  wire[1:0] net_io_clients_1_grant_bits_header_dst;
  wire[1:0] net_io_clients_1_grant_bits_header_src;
  wire net_io_clients_1_grant_valid;
  wire net_io_clients_1_acquire_ready;
  wire net_io_clients_0_release_ready;
  wire[1:0] net_io_clients_0_probe_bits_payload_p_type;
  wire[2:0] net_io_clients_0_probe_bits_payload_master_xact_id;
  wire[25:0] net_io_clients_0_probe_bits_payload_addr;
  wire[1:0] net_io_clients_0_probe_bits_header_dst;
  wire[1:0] net_io_clients_0_probe_bits_header_src;
  wire net_io_clients_0_probe_valid;
  wire net_io_clients_0_finish_ready;
  wire[3:0] net_io_clients_0_grant_bits_payload_g_type;
  wire[2:0] net_io_clients_0_grant_bits_payload_master_xact_id;
  wire[1:0] net_io_clients_0_grant_bits_payload_client_xact_id;
  wire[511:0] net_io_clients_0_grant_bits_payload_data;
  wire[1:0] net_io_clients_0_grant_bits_header_dst;
  wire[1:0] net_io_clients_0_grant_bits_header_src;
  wire net_io_clients_0_grant_valid;
  wire net_io_clients_0_acquire_ready;


  assign io_mem_req_data_bits_data = llc_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = llc_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = llc_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = llc_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = llc_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = llc_io_mem_req_cmd_valid;
  assign io_htif_release_ready = net_io_clients_1_release_ready;
  assign io_htif_probe_bits_payload_p_type = net_io_clients_1_probe_bits_payload_p_type;
  assign io_htif_probe_bits_payload_master_xact_id = net_io_clients_1_probe_bits_payload_master_xact_id;
  assign io_htif_probe_bits_payload_addr = net_io_clients_1_probe_bits_payload_addr;
  assign io_htif_probe_bits_header_dst = net_io_clients_1_probe_bits_header_dst;
  assign io_htif_probe_bits_header_src = net_io_clients_1_probe_bits_header_src;
  assign io_htif_probe_valid = net_io_clients_1_probe_valid;
  assign io_htif_finish_ready = net_io_clients_1_finish_ready;
  assign io_htif_grant_bits_payload_g_type = net_io_clients_1_grant_bits_payload_g_type;
  assign io_htif_grant_bits_payload_master_xact_id = net_io_clients_1_grant_bits_payload_master_xact_id;
  assign io_htif_grant_bits_payload_client_xact_id = net_io_clients_1_grant_bits_payload_client_xact_id;
  assign io_htif_grant_bits_payload_data = net_io_clients_1_grant_bits_payload_data;
  assign io_htif_grant_bits_header_dst = net_io_clients_1_grant_bits_header_dst;
  assign io_htif_grant_bits_header_src = net_io_clients_1_grant_bits_header_src;
  assign io_htif_grant_valid = net_io_clients_1_grant_valid;
  assign io_htif_acquire_ready = net_io_clients_1_acquire_ready;
  assign io_tiles_0_release_ready = net_io_clients_0_release_ready;
  assign io_tiles_0_probe_bits_payload_p_type = net_io_clients_0_probe_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = net_io_clients_0_probe_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = net_io_clients_0_probe_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = net_io_clients_0_probe_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = net_io_clients_0_probe_bits_header_src;
  assign io_tiles_0_probe_valid = net_io_clients_0_probe_valid;
  assign io_tiles_0_finish_ready = net_io_clients_0_finish_ready;
  assign io_tiles_0_grant_bits_payload_g_type = net_io_clients_0_grant_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = net_io_clients_0_grant_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = net_io_clients_0_grant_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = net_io_clients_0_grant_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = net_io_clients_0_grant_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = net_io_clients_0_grant_bits_header_src;
  assign io_tiles_0_grant_valid = net_io_clients_0_grant_valid;
  assign io_tiles_0_acquire_ready = net_io_clients_0_acquire_ready;
  RocketChipCrossbarNetwork net(.clk(clk), .reset(reset),
       .io_clients_1_acquire_ready( net_io_clients_1_acquire_ready ),
       .io_clients_1_acquire_valid( io_htif_acquire_valid ),
       .io_clients_1_acquire_bits_header_src( io_htif_acquire_bits_header_src ),
       .io_clients_1_acquire_bits_header_dst( io_htif_acquire_bits_header_dst ),
       .io_clients_1_acquire_bits_payload_addr( io_htif_acquire_bits_payload_addr ),
       .io_clients_1_acquire_bits_payload_client_xact_id( io_htif_acquire_bits_payload_client_xact_id ),
       .io_clients_1_acquire_bits_payload_data( io_htif_acquire_bits_payload_data ),
       .io_clients_1_acquire_bits_payload_a_type( io_htif_acquire_bits_payload_a_type ),
       .io_clients_1_acquire_bits_payload_write_mask( io_htif_acquire_bits_payload_write_mask ),
       .io_clients_1_acquire_bits_payload_subword_addr( io_htif_acquire_bits_payload_subword_addr ),
       .io_clients_1_acquire_bits_payload_atomic_opcode( io_htif_acquire_bits_payload_atomic_opcode ),
       .io_clients_1_grant_ready( io_htif_grant_ready ),
       .io_clients_1_grant_valid( net_io_clients_1_grant_valid ),
       .io_clients_1_grant_bits_header_src( net_io_clients_1_grant_bits_header_src ),
       .io_clients_1_grant_bits_header_dst( net_io_clients_1_grant_bits_header_dst ),
       .io_clients_1_grant_bits_payload_data( net_io_clients_1_grant_bits_payload_data ),
       .io_clients_1_grant_bits_payload_client_xact_id( net_io_clients_1_grant_bits_payload_client_xact_id ),
       .io_clients_1_grant_bits_payload_master_xact_id( net_io_clients_1_grant_bits_payload_master_xact_id ),
       .io_clients_1_grant_bits_payload_g_type( net_io_clients_1_grant_bits_payload_g_type ),
       .io_clients_1_finish_ready( net_io_clients_1_finish_ready ),
       .io_clients_1_finish_valid( io_htif_finish_valid ),
       .io_clients_1_finish_bits_header_src( io_htif_finish_bits_header_src ),
       .io_clients_1_finish_bits_header_dst( io_htif_finish_bits_header_dst ),
       .io_clients_1_finish_bits_payload_master_xact_id( io_htif_finish_bits_payload_master_xact_id ),
       .io_clients_1_probe_ready( io_htif_probe_ready ),
       .io_clients_1_probe_valid( net_io_clients_1_probe_valid ),
       .io_clients_1_probe_bits_header_src( net_io_clients_1_probe_bits_header_src ),
       .io_clients_1_probe_bits_header_dst( net_io_clients_1_probe_bits_header_dst ),
       .io_clients_1_probe_bits_payload_addr( net_io_clients_1_probe_bits_payload_addr ),
       .io_clients_1_probe_bits_payload_master_xact_id( net_io_clients_1_probe_bits_payload_master_xact_id ),
       .io_clients_1_probe_bits_payload_p_type( net_io_clients_1_probe_bits_payload_p_type ),
       .io_clients_1_release_ready( net_io_clients_1_release_ready ),
       .io_clients_1_release_valid( io_htif_release_valid ),
       .io_clients_1_release_bits_header_src( io_htif_release_bits_header_src ),
       .io_clients_1_release_bits_header_dst( io_htif_release_bits_header_dst ),
       .io_clients_1_release_bits_payload_addr( io_htif_release_bits_payload_addr ),
       .io_clients_1_release_bits_payload_client_xact_id( io_htif_release_bits_payload_client_xact_id ),
       .io_clients_1_release_bits_payload_master_xact_id( io_htif_release_bits_payload_master_xact_id ),
       .io_clients_1_release_bits_payload_data( io_htif_release_bits_payload_data ),
       .io_clients_1_release_bits_payload_r_type( io_htif_release_bits_payload_r_type ),
       .io_clients_0_acquire_ready( net_io_clients_0_acquire_ready ),
       .io_clients_0_acquire_valid( io_tiles_0_acquire_valid ),
       .io_clients_0_acquire_bits_header_src( io_tiles_0_acquire_bits_header_src ),
       .io_clients_0_acquire_bits_header_dst( io_tiles_0_acquire_bits_header_dst ),
       .io_clients_0_acquire_bits_payload_addr( io_tiles_0_acquire_bits_payload_addr ),
       .io_clients_0_acquire_bits_payload_client_xact_id( io_tiles_0_acquire_bits_payload_client_xact_id ),
       .io_clients_0_acquire_bits_payload_data( io_tiles_0_acquire_bits_payload_data ),
       .io_clients_0_acquire_bits_payload_a_type( io_tiles_0_acquire_bits_payload_a_type ),
       .io_clients_0_acquire_bits_payload_write_mask( io_tiles_0_acquire_bits_payload_write_mask ),
       .io_clients_0_acquire_bits_payload_subword_addr( io_tiles_0_acquire_bits_payload_subword_addr ),
       .io_clients_0_acquire_bits_payload_atomic_opcode( io_tiles_0_acquire_bits_payload_atomic_opcode ),
       .io_clients_0_grant_ready( io_tiles_0_grant_ready ),
       .io_clients_0_grant_valid( net_io_clients_0_grant_valid ),
       .io_clients_0_grant_bits_header_src( net_io_clients_0_grant_bits_header_src ),
       .io_clients_0_grant_bits_header_dst( net_io_clients_0_grant_bits_header_dst ),
       .io_clients_0_grant_bits_payload_data( net_io_clients_0_grant_bits_payload_data ),
       .io_clients_0_grant_bits_payload_client_xact_id( net_io_clients_0_grant_bits_payload_client_xact_id ),
       .io_clients_0_grant_bits_payload_master_xact_id( net_io_clients_0_grant_bits_payload_master_xact_id ),
       .io_clients_0_grant_bits_payload_g_type( net_io_clients_0_grant_bits_payload_g_type ),
       .io_clients_0_finish_ready( net_io_clients_0_finish_ready ),
       .io_clients_0_finish_valid( io_tiles_0_finish_valid ),
       .io_clients_0_finish_bits_header_src( io_tiles_0_finish_bits_header_src ),
       .io_clients_0_finish_bits_header_dst( io_tiles_0_finish_bits_header_dst ),
       .io_clients_0_finish_bits_payload_master_xact_id( io_tiles_0_finish_bits_payload_master_xact_id ),
       .io_clients_0_probe_ready( io_tiles_0_probe_ready ),
       .io_clients_0_probe_valid( net_io_clients_0_probe_valid ),
       .io_clients_0_probe_bits_header_src( net_io_clients_0_probe_bits_header_src ),
       .io_clients_0_probe_bits_header_dst( net_io_clients_0_probe_bits_header_dst ),
       .io_clients_0_probe_bits_payload_addr( net_io_clients_0_probe_bits_payload_addr ),
       .io_clients_0_probe_bits_payload_master_xact_id( net_io_clients_0_probe_bits_payload_master_xact_id ),
       .io_clients_0_probe_bits_payload_p_type( net_io_clients_0_probe_bits_payload_p_type ),
       .io_clients_0_release_ready( net_io_clients_0_release_ready ),
       .io_clients_0_release_valid( io_tiles_0_release_valid ),
       .io_clients_0_release_bits_header_src( io_tiles_0_release_bits_header_src ),
       .io_clients_0_release_bits_header_dst( io_tiles_0_release_bits_header_dst ),
       .io_clients_0_release_bits_payload_addr( io_tiles_0_release_bits_payload_addr ),
       .io_clients_0_release_bits_payload_client_xact_id( io_tiles_0_release_bits_payload_client_xact_id ),
       .io_clients_0_release_bits_payload_master_xact_id( io_tiles_0_release_bits_payload_master_xact_id ),
       .io_clients_0_release_bits_payload_data( io_tiles_0_release_bits_payload_data ),
       .io_clients_0_release_bits_payload_r_type( io_tiles_0_release_bits_payload_r_type ),
       .io_masters_0_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_masters_0_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_masters_0_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_masters_0_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_masters_0_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_masters_0_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_masters_0_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_masters_0_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_masters_0_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_masters_0_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_masters_0_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_masters_0_grant_ready( net_io_masters_0_grant_ready ),
       .io_masters_0_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_masters_0_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_masters_0_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_masters_0_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_masters_0_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_masters_0_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_masters_0_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_masters_0_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_masters_0_finish_valid( net_io_masters_0_finish_valid ),
       .io_masters_0_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_masters_0_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_masters_0_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_masters_0_probe_ready( net_io_masters_0_probe_ready ),
       .io_masters_0_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_masters_0_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_masters_0_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_masters_0_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_masters_0_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_masters_0_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_masters_0_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_masters_0_release_valid( net_io_masters_0_release_valid ),
       .io_masters_0_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_masters_0_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_masters_0_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_masters_0_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_masters_0_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_masters_0_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_masters_0_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type )
  );
  L2CoherenceAgent L2CoherenceAgent(.clk(clk), .reset(reset),
       .io_inner_acquire_ready( L2CoherenceAgent_io_inner_acquire_ready ),
       .io_inner_acquire_valid( net_io_masters_0_acquire_valid ),
       .io_inner_acquire_bits_header_src( net_io_masters_0_acquire_bits_header_src ),
       .io_inner_acquire_bits_header_dst( net_io_masters_0_acquire_bits_header_dst ),
       .io_inner_acquire_bits_payload_addr( net_io_masters_0_acquire_bits_payload_addr ),
       .io_inner_acquire_bits_payload_client_xact_id( net_io_masters_0_acquire_bits_payload_client_xact_id ),
       .io_inner_acquire_bits_payload_data( net_io_masters_0_acquire_bits_payload_data ),
       .io_inner_acquire_bits_payload_a_type( net_io_masters_0_acquire_bits_payload_a_type ),
       .io_inner_acquire_bits_payload_write_mask( net_io_masters_0_acquire_bits_payload_write_mask ),
       .io_inner_acquire_bits_payload_subword_addr( net_io_masters_0_acquire_bits_payload_subword_addr ),
       .io_inner_acquire_bits_payload_atomic_opcode( net_io_masters_0_acquire_bits_payload_atomic_opcode ),
       .io_inner_grant_ready( net_io_masters_0_grant_ready ),
       .io_inner_grant_valid( L2CoherenceAgent_io_inner_grant_valid ),
       .io_inner_grant_bits_header_src( L2CoherenceAgent_io_inner_grant_bits_header_src ),
       .io_inner_grant_bits_header_dst( L2CoherenceAgent_io_inner_grant_bits_header_dst ),
       .io_inner_grant_bits_payload_data( L2CoherenceAgent_io_inner_grant_bits_payload_data ),
       .io_inner_grant_bits_payload_client_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_client_xact_id ),
       .io_inner_grant_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_grant_bits_payload_master_xact_id ),
       .io_inner_grant_bits_payload_g_type( L2CoherenceAgent_io_inner_grant_bits_payload_g_type ),
       .io_inner_finish_ready( L2CoherenceAgent_io_inner_finish_ready ),
       .io_inner_finish_valid( net_io_masters_0_finish_valid ),
       .io_inner_finish_bits_header_src( net_io_masters_0_finish_bits_header_src ),
       .io_inner_finish_bits_header_dst( net_io_masters_0_finish_bits_header_dst ),
       .io_inner_finish_bits_payload_master_xact_id( net_io_masters_0_finish_bits_payload_master_xact_id ),
       .io_inner_probe_ready( net_io_masters_0_probe_ready ),
       .io_inner_probe_valid( L2CoherenceAgent_io_inner_probe_valid ),
       .io_inner_probe_bits_header_src( L2CoherenceAgent_io_inner_probe_bits_header_src ),
       .io_inner_probe_bits_header_dst( L2CoherenceAgent_io_inner_probe_bits_header_dst ),
       .io_inner_probe_bits_payload_addr( L2CoherenceAgent_io_inner_probe_bits_payload_addr ),
       .io_inner_probe_bits_payload_master_xact_id( L2CoherenceAgent_io_inner_probe_bits_payload_master_xact_id ),
       .io_inner_probe_bits_payload_p_type( L2CoherenceAgent_io_inner_probe_bits_payload_p_type ),
       .io_inner_release_ready( L2CoherenceAgent_io_inner_release_ready ),
       .io_inner_release_valid( net_io_masters_0_release_valid ),
       .io_inner_release_bits_header_src( net_io_masters_0_release_bits_header_src ),
       .io_inner_release_bits_header_dst( net_io_masters_0_release_bits_header_dst ),
       .io_inner_release_bits_payload_addr( net_io_masters_0_release_bits_payload_addr ),
       .io_inner_release_bits_payload_client_xact_id( net_io_masters_0_release_bits_payload_client_xact_id ),
       .io_inner_release_bits_payload_master_xact_id( net_io_masters_0_release_bits_payload_master_xact_id ),
       .io_inner_release_bits_payload_data( net_io_masters_0_release_bits_payload_data ),
       .io_inner_release_bits_payload_r_type( net_io_masters_0_release_bits_payload_r_type ),
       .io_outer_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_outer_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_outer_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_outer_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_outer_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_outer_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_outer_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_outer_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_outer_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_outer_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_outer_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_outer_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_outer_grant_valid( conv_io_uncached_grant_valid ),
       //.io_outer_grant_bits_header_src(  )
       //.io_outer_grant_bits_header_dst(  )
       .io_outer_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_outer_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_outer_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_outer_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_outer_finish_ready(  )
       .io_outer_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_outer_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_outer_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_outer_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_incoherent_1( io_incoherent_1 ),
       .io_incoherent_0( io_incoherent_0 )
  );
  `ifndef SYNTHESIS
    assign L2CoherenceAgent.io_outer_grant_bits_header_src = {1{$random}};
    assign L2CoherenceAgent.io_outer_grant_bits_header_dst = {1{$random}};
    assign L2CoherenceAgent.io_outer_finish_ready = {1{$random}};
  `endif
  MemIOUncachedTileLinkIOConverter conv(.clk(clk), .reset(reset),
       .io_uncached_acquire_ready( conv_io_uncached_acquire_ready ),
       .io_uncached_acquire_valid( L2CoherenceAgent_io_outer_acquire_valid ),
       .io_uncached_acquire_bits_header_src( L2CoherenceAgent_io_outer_acquire_bits_header_src ),
       .io_uncached_acquire_bits_header_dst( L2CoherenceAgent_io_outer_acquire_bits_header_dst ),
       .io_uncached_acquire_bits_payload_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_addr ),
       .io_uncached_acquire_bits_payload_client_xact_id( L2CoherenceAgent_io_outer_acquire_bits_payload_client_xact_id ),
       .io_uncached_acquire_bits_payload_data( L2CoherenceAgent_io_outer_acquire_bits_payload_data ),
       .io_uncached_acquire_bits_payload_a_type( L2CoherenceAgent_io_outer_acquire_bits_payload_a_type ),
       .io_uncached_acquire_bits_payload_write_mask( L2CoherenceAgent_io_outer_acquire_bits_payload_write_mask ),
       .io_uncached_acquire_bits_payload_subword_addr( L2CoherenceAgent_io_outer_acquire_bits_payload_subword_addr ),
       .io_uncached_acquire_bits_payload_atomic_opcode( L2CoherenceAgent_io_outer_acquire_bits_payload_atomic_opcode ),
       .io_uncached_grant_ready( L2CoherenceAgent_io_outer_grant_ready ),
       .io_uncached_grant_valid( conv_io_uncached_grant_valid ),
       //.io_uncached_grant_bits_header_src(  )
       //.io_uncached_grant_bits_header_dst(  )
       .io_uncached_grant_bits_payload_data( conv_io_uncached_grant_bits_payload_data ),
       .io_uncached_grant_bits_payload_client_xact_id( conv_io_uncached_grant_bits_payload_client_xact_id ),
       .io_uncached_grant_bits_payload_master_xact_id( conv_io_uncached_grant_bits_payload_master_xact_id ),
       .io_uncached_grant_bits_payload_g_type( conv_io_uncached_grant_bits_payload_g_type ),
       //.io_uncached_finish_ready(  )
       .io_uncached_finish_valid( L2CoherenceAgent_io_outer_finish_valid ),
       .io_uncached_finish_bits_header_src( L2CoherenceAgent_io_outer_finish_bits_header_src ),
       .io_uncached_finish_bits_header_dst( L2CoherenceAgent_io_outer_finish_bits_header_dst ),
       .io_uncached_finish_bits_payload_master_xact_id( L2CoherenceAgent_io_outer_finish_bits_payload_master_xact_id ),
       .io_mem_req_cmd_ready( Queue_0_io_enq_ready ),
       .io_mem_req_cmd_valid( conv_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( Queue_1_io_enq_ready ),
       .io_mem_req_data_valid( conv_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( conv_io_mem_req_data_bits_data ),
       .io_mem_resp_ready( conv_io_mem_resp_ready ),
       .io_mem_resp_valid( llc_io_cpu_resp_valid ),
       .io_mem_resp_bits_data( llc_io_cpu_resp_bits_data ),
       .io_mem_resp_bits_tag( llc_io_cpu_resp_bits_tag )
  );
  DRAMSideLLCNull llc(.clk(clk), .reset(reset),
       .io_cpu_req_cmd_ready( llc_io_cpu_req_cmd_ready ),
       .io_cpu_req_cmd_valid( Queue_0_io_deq_valid ),
       .io_cpu_req_cmd_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_cpu_req_cmd_bits_tag( Queue_0_io_deq_bits_tag ),
       .io_cpu_req_cmd_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_cpu_req_data_ready( llc_io_cpu_req_data_ready ),
       .io_cpu_req_data_valid( Queue_1_io_deq_valid ),
       .io_cpu_req_data_bits_data( Queue_1_io_deq_bits_data ),
       .io_cpu_resp_ready( conv_io_mem_resp_ready ),
       .io_cpu_resp_valid( llc_io_cpu_resp_valid ),
       .io_cpu_resp_bits_data( llc_io_cpu_resp_bits_data ),
       .io_cpu_resp_bits_tag( llc_io_cpu_resp_bits_tag ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( llc_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( llc_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( llc_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( llc_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( llc_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( llc_io_mem_req_data_bits_data ),
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
  );
  Queue_6 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_cmd_valid ),
       .io_enq_bits_addr( conv_io_mem_req_cmd_bits_addr ),
       .io_enq_bits_tag( conv_io_mem_req_cmd_bits_tag ),
       .io_enq_bits_rw( conv_io_mem_req_cmd_bits_rw ),
       .io_deq_ready( llc_io_cpu_req_cmd_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_tag( Queue_0_io_deq_bits_tag ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw )
  );
  Queue_7 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( conv_io_mem_req_data_valid ),
       .io_enq_bits_data( conv_io_mem_req_data_bits_data ),
       .io_deq_ready( llc_io_cpu_req_data_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_data( Queue_1_io_deq_bits_data )
  );
endmodule

module Queue_8(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_a_type,
    input [5:0] io_enq_bits_payload_write_mask,
    input [2:0] io_enq_bits_payload_subword_addr,
    input [3:0] io_enq_bits_payload_atomic_opcode,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_a_type,
    output[5:0] io_deq_bits_payload_write_mask,
    output[2:0] io_deq_bits_payload_subword_addr,
    output[3:0] io_deq_bits_payload_atomic_opcode
);

  wire[3:0] T0;
  wire[559:0] T1;
  reg [559:0] ram [1:0];
  wire[559:0] T2;
  wire[559:0] T3;
  wire[559:0] T4;
  wire[527:0] T5;
  wire[12:0] T6;
  wire[6:0] T7;
  wire[514:0] T8;
  wire[31:0] T9;
  wire[27:0] T10;
  wire[3:0] T11;
  wire do_enq;
  reg  R12;
  wire T13;
  wire T14;
  wire T15;
  reg  R16;
  wire T17;
  wire T18;
  wire T19;
  wire do_deq;
  wire[2:0] T20;
  wire[5:0] T21;
  wire[2:0] T22;
  wire[511:0] T23;
  wire[1:0] T24;
  wire[25:0] T25;
  wire[1:0] T26;
  wire[1:0] T27;
  wire T28;
  wire empty;
  wire T29;
  reg  maybe_full;
  wire T30;
  wire T31;
  wire T32;
  wire ptr_match;
  wire T33;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R12 = {1{$random}};
    R16 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_atomic_opcode = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[R16];
  assign T3 = T4;
  assign T4 = {T9, T5};
  assign T5 = {T8, T6};
  assign T6 = {io_enq_bits_payload_write_mask, T7};
  assign T7 = {io_enq_bits_payload_subword_addr, io_enq_bits_payload_atomic_opcode};
  assign T8 = {io_enq_bits_payload_data, io_enq_bits_payload_a_type};
  assign T9 = {T11, T10};
  assign T10 = {io_enq_bits_payload_addr, io_enq_bits_payload_client_xact_id};
  assign T11 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T13 = reset ? 1'h0 : T14;
  assign T14 = do_enq ? T15 : R12;
  assign T15 = R12 + 1'h1;
  assign T17 = reset ? 1'h0 : T18;
  assign T18 = do_deq ? T19 : R16;
  assign T19 = R16 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_subword_addr = T20;
  assign T20 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_write_mask = T21;
  assign T21 = T1[4'hc:3'h7];
  assign io_deq_bits_payload_a_type = T22;
  assign T22 = T1[4'hf:4'hd];
  assign io_deq_bits_payload_data = T23;
  assign T23 = T1[10'h20f:5'h10];
  assign io_deq_bits_payload_client_xact_id = T24;
  assign T24 = T1[10'h211:10'h210];
  assign io_deq_bits_payload_addr = T25;
  assign T25 = T1[10'h22b:10'h212];
  assign io_deq_bits_header_dst = T26;
  assign T26 = T1[10'h22d:10'h22c];
  assign io_deq_bits_header_src = T27;
  assign T27 = T1[10'h22f:10'h22e];
  assign io_deq_valid = T28;
  assign T28 = empty ^ 1'h1;
  assign empty = ptr_match & T29;
  assign T29 = maybe_full ^ 1'h1;
  assign T30 = reset ? 1'h0 : T31;
  assign T31 = T32 ? do_enq : maybe_full;
  assign T32 = do_enq != do_deq;
  assign ptr_match = R12 == R16;
  assign io_enq_ready = T33;
  assign T33 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R12] <= T3;
    if(reset) begin
      R12 <= 1'h0;
    end else if(do_enq) begin
      R12 <= T15;
    end
    if(reset) begin
      R16 <= 1'h0;
    end else if(do_deq) begin
      R16 <= T19;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T32) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_9(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [511:0] io_enq_bits_payload_data,
    input [2:0] io_enq_bits_payload_r_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[511:0] io_deq_bits_payload_data,
    output[2:0] io_deq_bits_payload_r_type
);

  wire[2:0] T0;
  wire[549:0] T1;
  reg [549:0] ram [1:0];
  wire[549:0] T2;
  wire[549:0] T3;
  wire[549:0] T4;
  wire[519:0] T5;
  wire[514:0] T6;
  wire[4:0] T7;
  wire[29:0] T8;
  wire[27:0] T9;
  wire do_enq;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  reg  R14;
  wire T15;
  wire T16;
  wire T17;
  wire do_deq;
  wire[511:0] T18;
  wire[2:0] T19;
  wire[1:0] T20;
  wire[25:0] T21;
  wire[1:0] T22;
  wire[1:0] T23;
  wire T24;
  wire empty;
  wire T25;
  reg  maybe_full;
  wire T26;
  wire T27;
  wire T28;
  wire ptr_match;
  wire T29;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {18{$random}};
    R10 = {1{$random}};
    R14 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_r_type = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R14];
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_enq_bits_payload_data, io_enq_bits_payload_r_type};
  assign T7 = {io_enq_bits_payload_client_xact_id, io_enq_bits_payload_master_xact_id};
  assign T8 = {io_enq_bits_header_src, T9};
  assign T9 = {io_enq_bits_header_dst, io_enq_bits_payload_addr};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_enq ? T13 : R10;
  assign T13 = R10 + 1'h1;
  assign T15 = reset ? 1'h0 : T16;
  assign T16 = do_deq ? T17 : R14;
  assign T17 = R14 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_data = T18;
  assign T18 = T1[10'h202:2'h3];
  assign io_deq_bits_payload_master_xact_id = T19;
  assign T19 = T1[10'h205:10'h203];
  assign io_deq_bits_payload_client_xact_id = T20;
  assign T20 = T1[10'h207:10'h206];
  assign io_deq_bits_payload_addr = T21;
  assign T21 = T1[10'h221:10'h208];
  assign io_deq_bits_header_dst = T22;
  assign T22 = T1[10'h223:10'h222];
  assign io_deq_bits_header_src = T23;
  assign T23 = T1[10'h225:10'h224];
  assign io_deq_valid = T24;
  assign T24 = empty ^ 1'h1;
  assign empty = ptr_match & T25;
  assign T25 = maybe_full ^ 1'h1;
  assign T26 = reset ? 1'h0 : T27;
  assign T27 = T28 ? do_enq : maybe_full;
  assign T28 = do_enq != do_deq;
  assign ptr_match = R10 == R14;
  assign io_enq_ready = T29;
  assign T29 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R10] <= T3;
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_enq) begin
      R10 <= T13;
    end
    if(reset) begin
      R14 <= 1'h0;
    end else if(do_deq) begin
      R14 <= T17;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T28) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_10(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[2:0] io_deq_bits_payload_master_xact_id
);

  wire[2:0] T0;
  wire[6:0] T1;
  reg [6:0] ram [1:0];
  wire[6:0] T2;
  wire[6:0] T3;
  wire[6:0] T4;
  wire[4:0] T5;
  wire do_enq;
  reg  R6;
  wire T7;
  wire T8;
  wire T9;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  wire do_deq;
  wire[1:0] T14;
  wire[1:0] T15;
  wire T16;
  wire empty;
  wire T17;
  reg  maybe_full;
  wire T18;
  wire T19;
  wire T20;
  wire ptr_match;
  wire T21;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R6 = {1{$random}};
    R10 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_master_xact_id = T0;
  assign T0 = T1[2'h2:1'h0];
  assign T1 = ram[R10];
  assign T3 = T4;
  assign T4 = {io_enq_bits_header_src, T5};
  assign T5 = {io_enq_bits_header_dst, io_enq_bits_payload_master_xact_id};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_enq ? T9 : R6;
  assign T9 = R6 + 1'h1;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_deq ? T13 : R10;
  assign T13 = R10 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_header_dst = T14;
  assign T14 = T1[3'h4:2'h3];
  assign io_deq_bits_header_src = T15;
  assign T15 = T1[3'h6:3'h5];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign T18 = reset ? 1'h0 : T19;
  assign T19 = T20 ? do_enq : maybe_full;
  assign T20 = do_enq != do_deq;
  assign ptr_match = R6 == R10;
  assign io_enq_ready = T21;
  assign T21 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T9;
    end
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_deq) begin
      R10 <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T20) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_11(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [511:0] io_enq_bits_payload_data,
    input [1:0] io_enq_bits_payload_client_xact_id,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [3:0] io_enq_bits_payload_g_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[511:0] io_deq_bits_payload_data,
    output[1:0] io_deq_bits_payload_client_xact_id,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[3:0] io_deq_bits_payload_g_type
);

  wire[3:0] T0;
  wire[524:0] T1;
  reg [524:0] ram [0:0];
  wire[524:0] T2;
  wire[524:0] T3;
  wire[524:0] T4;
  wire[8:0] T5;
  wire[6:0] T6;
  wire[515:0] T7;
  wire[513:0] T8;
  wire do_enq;
  wire[2:0] T9;
  wire[1:0] T10;
  wire[511:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire empty;
  reg  maybe_full;
  wire T15;
  wire T16;
  wire T17;
  wire do_deq;
  wire T18;
  wire T19;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 1; initvar = initvar+1)
      ram[initvar] = {17{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_g_type = T0;
  assign T0 = T1[2'h3:1'h0];
  assign T1 = ram[1'h0];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_client_xact_id, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_g_type};
  assign T7 = {io_enq_bits_header_src, T8};
  assign T8 = {io_enq_bits_header_dst, io_enq_bits_payload_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_deq_bits_payload_master_xact_id = T9;
  assign T9 = T1[3'h6:3'h4];
  assign io_deq_bits_payload_client_xact_id = T10;
  assign T10 = T1[4'h8:3'h7];
  assign io_deq_bits_payload_data = T11;
  assign T11 = T1[10'h208:4'h9];
  assign io_deq_bits_header_dst = T12;
  assign T12 = T1[10'h20a:10'h209];
  assign io_deq_bits_header_src = T13;
  assign T13 = T1[10'h20c:10'h20b];
  assign io_deq_valid = T14;
  assign T14 = empty ^ 1'h1;
  assign empty = maybe_full ^ 1'h1;
  assign T15 = reset ? 1'h0 : T16;
  assign T16 = T17 ? do_enq : maybe_full;
  assign T17 = do_enq != do_deq;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_enq_ready = T18;
  assign T18 = T19 | io_deq_ready;
  assign T19 = maybe_full ^ 1'h1;

  always @(posedge clk) begin
    if (do_enq)
      ram[1'h0] <= T3;
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T17) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_12(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [1:0] io_enq_bits_header_src,
    input [1:0] io_enq_bits_header_dst,
    input [25:0] io_enq_bits_payload_addr,
    input [2:0] io_enq_bits_payload_master_xact_id,
    input [1:0] io_enq_bits_payload_p_type,
    input  io_deq_ready,
    output io_deq_valid,
    output[1:0] io_deq_bits_header_src,
    output[1:0] io_deq_bits_header_dst,
    output[25:0] io_deq_bits_payload_addr,
    output[2:0] io_deq_bits_payload_master_xact_id,
    output[1:0] io_deq_bits_payload_p_type
);

  wire[1:0] T0;
  wire[34:0] T1;
  reg [34:0] ram [1:0];
  wire[34:0] T2;
  wire[34:0] T3;
  wire[34:0] T4;
  wire[30:0] T5;
  wire[4:0] T6;
  wire[3:0] T7;
  wire do_enq;
  reg  R8;
  wire T9;
  wire T10;
  wire T11;
  reg  R12;
  wire T13;
  wire T14;
  wire T15;
  wire do_deq;
  wire[2:0] T16;
  wire[25:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire T20;
  wire empty;
  wire T21;
  reg  maybe_full;
  wire T22;
  wire T23;
  wire T24;
  wire ptr_match;
  wire T25;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R8 = {1{$random}};
    R12 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_payload_p_type = T0;
  assign T0 = T1[1'h1:1'h0];
  assign T1 = ram[R12];
  assign T3 = T4;
  assign T4 = {T7, T5};
  assign T5 = {io_enq_bits_payload_addr, T6};
  assign T6 = {io_enq_bits_payload_master_xact_id, io_enq_bits_payload_p_type};
  assign T7 = {io_enq_bits_header_src, io_enq_bits_header_dst};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T9 = reset ? 1'h0 : T10;
  assign T10 = do_enq ? T11 : R8;
  assign T11 = R8 + 1'h1;
  assign T13 = reset ? 1'h0 : T14;
  assign T14 = do_deq ? T15 : R12;
  assign T15 = R12 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_payload_master_xact_id = T16;
  assign T16 = T1[3'h4:2'h2];
  assign io_deq_bits_payload_addr = T17;
  assign T17 = T1[5'h1e:3'h5];
  assign io_deq_bits_header_dst = T18;
  assign T18 = T1[6'h20:5'h1f];
  assign io_deq_bits_header_src = T19;
  assign T19 = T1[6'h22:6'h21];
  assign io_deq_valid = T20;
  assign T20 = empty ^ 1'h1;
  assign empty = ptr_match & T21;
  assign T21 = maybe_full ^ 1'h1;
  assign T22 = reset ? 1'h0 : T23;
  assign T23 = T24 ? do_enq : maybe_full;
  assign T24 = do_enq != do_deq;
  assign ptr_match = R8 == R12;
  assign io_enq_ready = T25;
  assign T25 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R8] <= T3;
    if(reset) begin
      R8 <= 1'h0;
    end else if(do_enq) begin
      R8 <= T11;
    end
    if(reset) begin
      R12 <= 1'h0;
    end else if(do_deq) begin
      R12 <= T15;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T24) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Uncore(input clk, input reset,
    //output io_host_clk
    //output io_host_clk_edge
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    //output io_mem_resp_ready
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    output io_tiles_0_acquire_ready,
    input  io_tiles_0_acquire_valid,
    input [1:0] io_tiles_0_acquire_bits_header_src,
    input [1:0] io_tiles_0_acquire_bits_header_dst,
    input [25:0] io_tiles_0_acquire_bits_payload_addr,
    input [1:0] io_tiles_0_acquire_bits_payload_client_xact_id,
    input [511:0] io_tiles_0_acquire_bits_payload_data,
    input [2:0] io_tiles_0_acquire_bits_payload_a_type,
    input [5:0] io_tiles_0_acquire_bits_payload_write_mask,
    input [2:0] io_tiles_0_acquire_bits_payload_subword_addr,
    input [3:0] io_tiles_0_acquire_bits_payload_atomic_opcode,
    input  io_tiles_0_grant_ready,
    output io_tiles_0_grant_valid,
    output[1:0] io_tiles_0_grant_bits_header_src,
    output[1:0] io_tiles_0_grant_bits_header_dst,
    output[511:0] io_tiles_0_grant_bits_payload_data,
    output[1:0] io_tiles_0_grant_bits_payload_client_xact_id,
    output[2:0] io_tiles_0_grant_bits_payload_master_xact_id,
    output[3:0] io_tiles_0_grant_bits_payload_g_type,
    output io_tiles_0_finish_ready,
    input  io_tiles_0_finish_valid,
    input [1:0] io_tiles_0_finish_bits_header_src,
    input [1:0] io_tiles_0_finish_bits_header_dst,
    input [2:0] io_tiles_0_finish_bits_payload_master_xact_id,
    input  io_tiles_0_probe_ready,
    output io_tiles_0_probe_valid,
    output[1:0] io_tiles_0_probe_bits_header_src,
    output[1:0] io_tiles_0_probe_bits_header_dst,
    output[25:0] io_tiles_0_probe_bits_payload_addr,
    output[2:0] io_tiles_0_probe_bits_payload_master_xact_id,
    output[1:0] io_tiles_0_probe_bits_payload_p_type,
    output io_tiles_0_release_ready,
    input  io_tiles_0_release_valid,
    input [1:0] io_tiles_0_release_bits_header_src,
    input [1:0] io_tiles_0_release_bits_header_dst,
    input [25:0] io_tiles_0_release_bits_payload_addr,
    input [1:0] io_tiles_0_release_bits_payload_client_xact_id,
    input [2:0] io_tiles_0_release_bits_payload_master_xact_id,
    input [511:0] io_tiles_0_release_bits_payload_data,
    input [2:0] io_tiles_0_release_bits_payload_r_type,
    output io_htif_0_reset,
    //output io_htif_0_id
    input  io_htif_0_pcr_req_ready,
    output io_htif_0_pcr_req_valid,
    output io_htif_0_pcr_req_bits_rw,
    output[4:0] io_htif_0_pcr_req_bits_addr,
    output[63:0] io_htif_0_pcr_req_bits_data,
    output io_htif_0_pcr_rep_ready,
    input  io_htif_0_pcr_rep_valid,
    input [63:0] io_htif_0_pcr_rep_bits,
    output io_htif_0_ipi_req_ready,
    input  io_htif_0_ipi_req_valid,
    input  io_htif_0_ipi_req_bits,
    input  io_htif_0_ipi_rep_ready,
    output io_htif_0_ipi_rep_valid,
    output io_htif_0_ipi_rep_bits,
    input  io_htif_0_debug_stats_pcr,
    input  io_incoherent_0
    //input  io_mem_backup_req_ready
    //output io_mem_backup_req_valid
    //output[15:0] io_mem_backup_req_bits
    //input  io_mem_backup_resp_valid
    //input [15:0] io_mem_backup_resp_bits
    //input  io_mem_backup_en
);

  wire htif_io_mem_probe_ready;
  wire[1:0] outmemsys_io_htif_probe_bits_payload_p_type;
  wire[2:0] outmemsys_io_htif_probe_bits_payload_master_xact_id;
  wire[25:0] outmemsys_io_htif_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_htif_probe_bits_header_dst;
  wire[1:0] outmemsys_io_htif_probe_bits_header_src;
  wire outmemsys_io_htif_probe_valid;
  wire htif_io_mem_grant_ready;
  wire[3:0] outmemsys_io_htif_grant_bits_payload_g_type;
  wire[2:0] outmemsys_io_htif_grant_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_htif_grant_bits_payload_client_xact_id;
  wire[511:0] outmemsys_io_htif_grant_bits_payload_data;
  wire[1:0] outmemsys_io_htif_grant_bits_header_dst;
  wire[1:0] outmemsys_io_htif_grant_bits_header_src;
  wire outmemsys_io_htif_grant_valid;
  wire outmemsys_io_htif_finish_ready;
  wire[2:0] T0;
  wire[2:0] htif_io_mem_finish_bits_payload_master_xact_id;
  wire[1:0] T1;
  wire[1:0] htif_io_mem_finish_bits_header_dst;
  wire[1:0] T2;
  wire T3;
  wire htif_io_mem_finish_valid;
  wire outmemsys_io_htif_release_ready;
  wire[2:0] T4;
  wire[2:0] htif_io_mem_release_bits_payload_r_type;
  wire[511:0] T5;
  wire[511:0] htif_io_mem_release_bits_payload_data;
  wire[2:0] T6;
  wire[2:0] htif_io_mem_release_bits_payload_master_xact_id;
  wire[1:0] T7;
  wire[1:0] htif_io_mem_release_bits_payload_client_xact_id;
  wire[25:0] T8;
  wire[25:0] htif_io_mem_release_bits_payload_addr;
  wire[1:0] T9;
  wire[1:0] T10;
  wire T11;
  wire htif_io_mem_release_valid;
  wire outmemsys_io_htif_acquire_ready;
  wire[3:0] T12;
  wire[3:0] htif_io_mem_acquire_bits_payload_atomic_opcode;
  wire[2:0] T13;
  wire[2:0] htif_io_mem_acquire_bits_payload_subword_addr;
  wire[5:0] T14;
  wire[5:0] htif_io_mem_acquire_bits_payload_write_mask;
  wire[2:0] T15;
  wire[2:0] htif_io_mem_acquire_bits_payload_a_type;
  wire[511:0] T16;
  wire[511:0] htif_io_mem_acquire_bits_payload_data;
  wire[1:0] T17;
  wire[1:0] htif_io_mem_acquire_bits_payload_client_xact_id;
  wire[25:0] T18;
  wire[25:0] htif_io_mem_acquire_bits_payload_addr;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire htif_io_mem_acquire_valid;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_payload_p_type;
  wire[2:0] outmemsys_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[25:0] outmemsys_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_dst;
  wire[1:0] outmemsys_io_tiles_0_probe_bits_header_src;
  wire outmemsys_io_tiles_0_probe_valid;
  wire[3:0] outmemsys_io_tiles_0_grant_bits_payload_g_type;
  wire[2:0] outmemsys_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[511:0] outmemsys_io_tiles_0_grant_bits_payload_data;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_dst;
  wire[1:0] outmemsys_io_tiles_0_grant_bits_header_src;
  wire outmemsys_io_tiles_0_grant_valid;
  wire outmemsys_io_tiles_0_finish_ready;
  wire[2:0] T22;
  wire[1:0] T23;
  wire[1:0] T24;
  wire T25;
  wire outmemsys_io_tiles_0_release_ready;
  wire[2:0] T26;
  wire[511:0] T27;
  wire[2:0] T28;
  wire[1:0] T29;
  wire[25:0] T30;
  wire[1:0] T31;
  wire[1:0] T32;
  wire T33;
  wire outmemsys_io_tiles_0_acquire_ready;
  wire[3:0] T34;
  wire[2:0] T35;
  wire[5:0] T36;
  wire[2:0] T37;
  wire[511:0] T38;
  wire[1:0] T39;
  wire[25:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire[2:0] Queue_6_io_deq_bits_payload_r_type;
  wire[511:0] Queue_6_io_deq_bits_payload_data;
  wire[2:0] Queue_6_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_6_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_6_io_deq_bits_payload_addr;
  wire[1:0] Queue_6_io_deq_bits_header_dst;
  wire[1:0] Queue_6_io_deq_bits_header_src;
  wire Queue_6_io_deq_valid;
  wire Queue_9_io_enq_ready;
  wire[2:0] Queue_7_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_7_io_deq_bits_header_dst;
  wire[1:0] Queue_7_io_deq_bits_header_src;
  wire Queue_7_io_deq_valid;
  wire Queue_8_io_enq_ready;
  wire[3:0] Queue_5_io_deq_bits_payload_atomic_opcode;
  wire[2:0] Queue_5_io_deq_bits_payload_subword_addr;
  wire[5:0] Queue_5_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_5_io_deq_bits_payload_a_type;
  wire[511:0] Queue_5_io_deq_bits_payload_data;
  wire[1:0] Queue_5_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_5_io_deq_bits_payload_addr;
  wire[1:0] Queue_5_io_deq_bits_header_dst;
  wire[1:0] Queue_5_io_deq_bits_header_src;
  wire Queue_5_io_deq_valid;
  wire[2:0] Queue_1_io_deq_bits_payload_r_type;
  wire[511:0] Queue_1_io_deq_bits_payload_data;
  wire[2:0] Queue_1_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_1_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_1_io_deq_bits_payload_addr;
  wire[1:0] Queue_1_io_deq_bits_header_dst;
  wire[1:0] Queue_1_io_deq_bits_header_src;
  wire Queue_1_io_deq_valid;
  wire Queue_4_io_enq_ready;
  wire[2:0] Queue_2_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_2_io_deq_bits_header_dst;
  wire[1:0] Queue_2_io_deq_bits_header_src;
  wire Queue_2_io_deq_valid;
  wire Queue_3_io_enq_ready;
  wire[3:0] Queue_0_io_deq_bits_payload_atomic_opcode;
  wire[2:0] Queue_0_io_deq_bits_payload_subword_addr;
  wire[5:0] Queue_0_io_deq_bits_payload_write_mask;
  wire[2:0] Queue_0_io_deq_bits_payload_a_type;
  wire[511:0] Queue_0_io_deq_bits_payload_data;
  wire[1:0] Queue_0_io_deq_bits_payload_client_xact_id;
  wire[25:0] Queue_0_io_deq_bits_payload_addr;
  wire[1:0] Queue_0_io_deq_bits_header_dst;
  wire[1:0] Queue_0_io_deq_bits_header_src;
  wire Queue_0_io_deq_valid;
  wire T44;
  wire Queue_6_io_enq_ready;
  wire[1:0] Queue_9_io_deq_bits_payload_p_type;
  wire[2:0] Queue_9_io_deq_bits_payload_master_xact_id;
  wire[25:0] Queue_9_io_deq_bits_payload_addr;
  wire[1:0] Queue_9_io_deq_bits_header_dst;
  wire[1:0] Queue_9_io_deq_bits_header_src;
  wire Queue_9_io_deq_valid;
  wire T45;
  wire Queue_7_io_enq_ready;
  wire[3:0] Queue_8_io_deq_bits_payload_g_type;
  wire[2:0] Queue_8_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_8_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_8_io_deq_bits_payload_data;
  wire[1:0] Queue_8_io_deq_bits_header_dst;
  wire[1:0] Queue_8_io_deq_bits_header_src;
  wire Queue_8_io_deq_valid;
  wire T46;
  wire Queue_5_io_enq_ready;
  wire htif_io_cpu_0_ipi_rep_valid;
  wire htif_io_cpu_0_ipi_req_ready;
  wire htif_io_cpu_0_pcr_rep_ready;
  wire[63:0] htif_io_cpu_0_pcr_req_bits_data;
  wire[4:0] htif_io_cpu_0_pcr_req_bits_addr;
  wire htif_io_cpu_0_pcr_req_bits_rw;
  wire htif_io_cpu_0_pcr_req_valid;
  wire htif_io_cpu_0_reset;
  wire T47;
  wire Queue_1_io_enq_ready;
  wire[1:0] Queue_4_io_deq_bits_payload_p_type;
  wire[2:0] Queue_4_io_deq_bits_payload_master_xact_id;
  wire[25:0] Queue_4_io_deq_bits_payload_addr;
  wire[1:0] Queue_4_io_deq_bits_header_dst;
  wire[1:0] Queue_4_io_deq_bits_header_src;
  wire Queue_4_io_deq_valid;
  wire T48;
  wire Queue_2_io_enq_ready;
  wire[3:0] Queue_3_io_deq_bits_payload_g_type;
  wire[2:0] Queue_3_io_deq_bits_payload_master_xact_id;
  wire[1:0] Queue_3_io_deq_bits_payload_client_xact_id;
  wire[511:0] Queue_3_io_deq_bits_payload_data;
  wire[1:0] Queue_3_io_deq_bits_header_dst;
  wire[1:0] Queue_3_io_deq_bits_header_src;
  wire Queue_3_io_deq_valid;
  wire T49;
  wire Queue_0_io_enq_ready;
  wire[127:0] outmemsys_io_mem_req_data_bits_data;
  wire outmemsys_io_mem_req_data_valid;
  wire outmemsys_io_mem_req_cmd_bits_rw;
  wire[4:0] outmemsys_io_mem_req_cmd_bits_tag;
  wire[25:0] outmemsys_io_mem_req_cmd_bits_addr;
  wire outmemsys_io_mem_req_cmd_valid;
  wire htif_io_host_debug_stats_pcr;
  wire[15:0] htif_io_host_out_bits;
  wire htif_io_host_out_valid;
  wire htif_io_host_in_ready;


  assign T0 = htif_io_mem_finish_bits_payload_master_xact_id;
  assign T1 = htif_io_mem_finish_bits_header_dst;
  assign T2 = 2'h1;
  assign T3 = htif_io_mem_finish_valid;
  assign T4 = htif_io_mem_release_bits_payload_r_type;
  assign T5 = htif_io_mem_release_bits_payload_data;
  assign T6 = htif_io_mem_release_bits_payload_master_xact_id;
  assign T7 = htif_io_mem_release_bits_payload_client_xact_id;
  assign T8 = htif_io_mem_release_bits_payload_addr;
  assign T9 = 2'h0;
  assign T10 = 2'h1;
  assign T11 = htif_io_mem_release_valid;
  assign T12 = htif_io_mem_acquire_bits_payload_atomic_opcode;
  assign T13 = htif_io_mem_acquire_bits_payload_subword_addr;
  assign T14 = htif_io_mem_acquire_bits_payload_write_mask;
  assign T15 = htif_io_mem_acquire_bits_payload_a_type;
  assign T16 = htif_io_mem_acquire_bits_payload_data;
  assign T17 = htif_io_mem_acquire_bits_payload_client_xact_id;
  assign T18 = htif_io_mem_acquire_bits_payload_addr;
  assign T19 = 2'h0;
  assign T20 = 2'h1;
  assign T21 = htif_io_mem_acquire_valid;
  assign T22 = io_tiles_0_finish_bits_payload_master_xact_id;
  assign T23 = io_tiles_0_finish_bits_header_dst;
  assign T24 = 2'h0;
  assign T25 = io_tiles_0_finish_valid;
  assign T26 = io_tiles_0_release_bits_payload_r_type;
  assign T27 = io_tiles_0_release_bits_payload_data;
  assign T28 = io_tiles_0_release_bits_payload_master_xact_id;
  assign T29 = io_tiles_0_release_bits_payload_client_xact_id;
  assign T30 = io_tiles_0_release_bits_payload_addr;
  assign T31 = 2'h0;
  assign T32 = 2'h0;
  assign T33 = io_tiles_0_release_valid;
  assign T34 = io_tiles_0_acquire_bits_payload_atomic_opcode;
  assign T35 = io_tiles_0_acquire_bits_payload_subword_addr;
  assign T36 = io_tiles_0_acquire_bits_payload_write_mask;
  assign T37 = io_tiles_0_acquire_bits_payload_a_type;
  assign T38 = io_tiles_0_acquire_bits_payload_data;
  assign T39 = io_tiles_0_acquire_bits_payload_client_xact_id;
  assign T40 = io_tiles_0_acquire_bits_payload_addr;
  assign T41 = 2'h0;
  assign T42 = 2'h0;
  assign T43 = io_tiles_0_acquire_valid;
  assign T44 = Queue_6_io_enq_ready;
  assign T45 = Queue_7_io_enq_ready;
  assign T46 = Queue_5_io_enq_ready;
  assign io_htif_0_ipi_rep_valid = htif_io_cpu_0_ipi_rep_valid;
  assign io_htif_0_ipi_req_ready = htif_io_cpu_0_ipi_req_ready;
  assign io_htif_0_pcr_rep_ready = htif_io_cpu_0_pcr_rep_ready;
  assign io_htif_0_pcr_req_bits_data = htif_io_cpu_0_pcr_req_bits_data;
  assign io_htif_0_pcr_req_bits_addr = htif_io_cpu_0_pcr_req_bits_addr;
  assign io_htif_0_pcr_req_bits_rw = htif_io_cpu_0_pcr_req_bits_rw;
  assign io_htif_0_pcr_req_valid = htif_io_cpu_0_pcr_req_valid;
  assign io_htif_0_reset = htif_io_cpu_0_reset;
  assign io_tiles_0_release_ready = T47;
  assign T47 = Queue_1_io_enq_ready;
  assign io_tiles_0_probe_bits_payload_p_type = Queue_4_io_deq_bits_payload_p_type;
  assign io_tiles_0_probe_bits_payload_master_xact_id = Queue_4_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_probe_bits_payload_addr = Queue_4_io_deq_bits_payload_addr;
  assign io_tiles_0_probe_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_tiles_0_probe_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_tiles_0_probe_valid = Queue_4_io_deq_valid;
  assign io_tiles_0_finish_ready = T48;
  assign T48 = Queue_2_io_enq_ready;
  assign io_tiles_0_grant_bits_payload_g_type = Queue_3_io_deq_bits_payload_g_type;
  assign io_tiles_0_grant_bits_payload_master_xact_id = Queue_3_io_deq_bits_payload_master_xact_id;
  assign io_tiles_0_grant_bits_payload_client_xact_id = Queue_3_io_deq_bits_payload_client_xact_id;
  assign io_tiles_0_grant_bits_payload_data = Queue_3_io_deq_bits_payload_data;
  assign io_tiles_0_grant_bits_header_dst = Queue_3_io_deq_bits_header_dst;
  assign io_tiles_0_grant_bits_header_src = Queue_3_io_deq_bits_header_src;
  assign io_tiles_0_grant_valid = Queue_3_io_deq_valid;
  assign io_tiles_0_acquire_ready = T49;
  assign T49 = Queue_0_io_enq_ready;
  assign io_mem_req_data_bits_data = outmemsys_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = outmemsys_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = outmemsys_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = outmemsys_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = outmemsys_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = outmemsys_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = htif_io_host_debug_stats_pcr;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_in_ready = htif_io_host_in_ready;
  HTIF htif(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( htif_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( htif_io_host_out_valid ),
       .io_host_out_bits( htif_io_host_out_bits ),
       .io_host_debug_stats_pcr( htif_io_host_debug_stats_pcr ),
       .io_cpu_0_reset( htif_io_cpu_0_reset ),
       //.io_cpu_0_id(  )
       .io_cpu_0_pcr_req_ready( io_htif_0_pcr_req_ready ),
       .io_cpu_0_pcr_req_valid( htif_io_cpu_0_pcr_req_valid ),
       .io_cpu_0_pcr_req_bits_rw( htif_io_cpu_0_pcr_req_bits_rw ),
       .io_cpu_0_pcr_req_bits_addr( htif_io_cpu_0_pcr_req_bits_addr ),
       .io_cpu_0_pcr_req_bits_data( htif_io_cpu_0_pcr_req_bits_data ),
       .io_cpu_0_pcr_rep_ready( htif_io_cpu_0_pcr_rep_ready ),
       .io_cpu_0_pcr_rep_valid( io_htif_0_pcr_rep_valid ),
       .io_cpu_0_pcr_rep_bits( io_htif_0_pcr_rep_bits ),
       .io_cpu_0_ipi_req_ready( htif_io_cpu_0_ipi_req_ready ),
       .io_cpu_0_ipi_req_valid( io_htif_0_ipi_req_valid ),
       .io_cpu_0_ipi_req_bits( io_htif_0_ipi_req_bits ),
       .io_cpu_0_ipi_rep_ready( io_htif_0_ipi_rep_ready ),
       .io_cpu_0_ipi_rep_valid( htif_io_cpu_0_ipi_rep_valid ),
       //.io_cpu_0_ipi_rep_bits(  )
       .io_cpu_0_debug_stats_pcr( io_htif_0_debug_stats_pcr ),
       .io_mem_acquire_ready( T46 ),
       .io_mem_acquire_valid( htif_io_mem_acquire_valid ),
       //.io_mem_acquire_bits_header_src(  )
       //.io_mem_acquire_bits_header_dst(  )
       .io_mem_acquire_bits_payload_addr( htif_io_mem_acquire_bits_payload_addr ),
       .io_mem_acquire_bits_payload_client_xact_id( htif_io_mem_acquire_bits_payload_client_xact_id ),
       .io_mem_acquire_bits_payload_data( htif_io_mem_acquire_bits_payload_data ),
       .io_mem_acquire_bits_payload_a_type( htif_io_mem_acquire_bits_payload_a_type ),
       .io_mem_acquire_bits_payload_write_mask( htif_io_mem_acquire_bits_payload_write_mask ),
       .io_mem_acquire_bits_payload_subword_addr( htif_io_mem_acquire_bits_payload_subword_addr ),
       .io_mem_acquire_bits_payload_atomic_opcode( htif_io_mem_acquire_bits_payload_atomic_opcode ),
       .io_mem_grant_ready( htif_io_mem_grant_ready ),
       .io_mem_grant_valid( Queue_8_io_deq_valid ),
       .io_mem_grant_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_mem_grant_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_mem_grant_bits_payload_data( Queue_8_io_deq_bits_payload_data ),
       .io_mem_grant_bits_payload_client_xact_id( Queue_8_io_deq_bits_payload_client_xact_id ),
       .io_mem_grant_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_mem_grant_bits_payload_g_type( Queue_8_io_deq_bits_payload_g_type ),
       .io_mem_finish_ready( T45 ),
       .io_mem_finish_valid( htif_io_mem_finish_valid ),
       //.io_mem_finish_bits_header_src(  )
       .io_mem_finish_bits_header_dst( htif_io_mem_finish_bits_header_dst ),
       .io_mem_finish_bits_payload_master_xact_id( htif_io_mem_finish_bits_payload_master_xact_id ),
       .io_mem_probe_ready( htif_io_mem_probe_ready ),
       .io_mem_probe_valid( Queue_9_io_deq_valid ),
       .io_mem_probe_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_mem_probe_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_mem_probe_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_mem_probe_bits_payload_master_xact_id( Queue_9_io_deq_bits_payload_master_xact_id ),
       .io_mem_probe_bits_payload_p_type( Queue_9_io_deq_bits_payload_p_type ),
       .io_mem_release_ready( T44 ),
       .io_mem_release_valid( htif_io_mem_release_valid ),
       //.io_mem_release_bits_header_src(  )
       //.io_mem_release_bits_header_dst(  )
       .io_mem_release_bits_payload_addr( htif_io_mem_release_bits_payload_addr ),
       .io_mem_release_bits_payload_client_xact_id( htif_io_mem_release_bits_payload_client_xact_id ),
       .io_mem_release_bits_payload_master_xact_id( htif_io_mem_release_bits_payload_master_xact_id ),
       .io_mem_release_bits_payload_data( htif_io_mem_release_bits_payload_data ),
       .io_mem_release_bits_payload_r_type( htif_io_mem_release_bits_payload_r_type )
       //.io_scr_rdata_63(  )
       //.io_scr_rdata_62(  )
       //.io_scr_rdata_61(  )
       //.io_scr_rdata_60(  )
       //.io_scr_rdata_59(  )
       //.io_scr_rdata_58(  )
       //.io_scr_rdata_57(  )
       //.io_scr_rdata_56(  )
       //.io_scr_rdata_55(  )
       //.io_scr_rdata_54(  )
       //.io_scr_rdata_53(  )
       //.io_scr_rdata_52(  )
       //.io_scr_rdata_51(  )
       //.io_scr_rdata_50(  )
       //.io_scr_rdata_49(  )
       //.io_scr_rdata_48(  )
       //.io_scr_rdata_47(  )
       //.io_scr_rdata_46(  )
       //.io_scr_rdata_45(  )
       //.io_scr_rdata_44(  )
       //.io_scr_rdata_43(  )
       //.io_scr_rdata_42(  )
       //.io_scr_rdata_41(  )
       //.io_scr_rdata_40(  )
       //.io_scr_rdata_39(  )
       //.io_scr_rdata_38(  )
       //.io_scr_rdata_37(  )
       //.io_scr_rdata_36(  )
       //.io_scr_rdata_35(  )
       //.io_scr_rdata_34(  )
       //.io_scr_rdata_33(  )
       //.io_scr_rdata_32(  )
       //.io_scr_rdata_31(  )
       //.io_scr_rdata_30(  )
       //.io_scr_rdata_29(  )
       //.io_scr_rdata_28(  )
       //.io_scr_rdata_27(  )
       //.io_scr_rdata_26(  )
       //.io_scr_rdata_25(  )
       //.io_scr_rdata_24(  )
       //.io_scr_rdata_23(  )
       //.io_scr_rdata_22(  )
       //.io_scr_rdata_21(  )
       //.io_scr_rdata_20(  )
       //.io_scr_rdata_19(  )
       //.io_scr_rdata_18(  )
       //.io_scr_rdata_17(  )
       //.io_scr_rdata_16(  )
       //.io_scr_rdata_15(  )
       //.io_scr_rdata_14(  )
       //.io_scr_rdata_13(  )
       //.io_scr_rdata_12(  )
       //.io_scr_rdata_11(  )
       //.io_scr_rdata_10(  )
       //.io_scr_rdata_9(  )
       //.io_scr_rdata_8(  )
       //.io_scr_rdata_7(  )
       //.io_scr_rdata_6(  )
       //.io_scr_rdata_5(  )
       //.io_scr_rdata_4(  )
       //.io_scr_rdata_3(  )
       //.io_scr_rdata_2(  )
       //.io_scr_rdata_1(  )
       //.io_scr_rdata_0(  )
       //.io_scr_wen(  )
       //.io_scr_waddr(  )
       //.io_scr_wdata(  )
  );
  `ifndef SYNTHESIS
    assign htif.io_mem_release_bits_payload_addr = {1{$random}};
    assign htif.io_mem_release_bits_payload_client_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_master_xact_id = {1{$random}};
    assign htif.io_mem_release_bits_payload_data = {16{$random}};
    assign htif.io_mem_release_bits_payload_r_type = {1{$random}};
    assign htif.io_scr_rdata_63 = {2{$random}};
    assign htif.io_scr_rdata_62 = {2{$random}};
    assign htif.io_scr_rdata_61 = {2{$random}};
    assign htif.io_scr_rdata_60 = {2{$random}};
    assign htif.io_scr_rdata_59 = {2{$random}};
    assign htif.io_scr_rdata_58 = {2{$random}};
    assign htif.io_scr_rdata_57 = {2{$random}};
    assign htif.io_scr_rdata_56 = {2{$random}};
    assign htif.io_scr_rdata_55 = {2{$random}};
    assign htif.io_scr_rdata_54 = {2{$random}};
    assign htif.io_scr_rdata_53 = {2{$random}};
    assign htif.io_scr_rdata_52 = {2{$random}};
    assign htif.io_scr_rdata_51 = {2{$random}};
    assign htif.io_scr_rdata_50 = {2{$random}};
    assign htif.io_scr_rdata_49 = {2{$random}};
    assign htif.io_scr_rdata_48 = {2{$random}};
    assign htif.io_scr_rdata_47 = {2{$random}};
    assign htif.io_scr_rdata_46 = {2{$random}};
    assign htif.io_scr_rdata_45 = {2{$random}};
    assign htif.io_scr_rdata_44 = {2{$random}};
    assign htif.io_scr_rdata_43 = {2{$random}};
    assign htif.io_scr_rdata_42 = {2{$random}};
    assign htif.io_scr_rdata_41 = {2{$random}};
    assign htif.io_scr_rdata_40 = {2{$random}};
    assign htif.io_scr_rdata_39 = {2{$random}};
    assign htif.io_scr_rdata_38 = {2{$random}};
    assign htif.io_scr_rdata_37 = {2{$random}};
    assign htif.io_scr_rdata_36 = {2{$random}};
    assign htif.io_scr_rdata_35 = {2{$random}};
    assign htif.io_scr_rdata_34 = {2{$random}};
    assign htif.io_scr_rdata_33 = {2{$random}};
    assign htif.io_scr_rdata_32 = {2{$random}};
    assign htif.io_scr_rdata_31 = {2{$random}};
    assign htif.io_scr_rdata_30 = {2{$random}};
    assign htif.io_scr_rdata_29 = {2{$random}};
    assign htif.io_scr_rdata_28 = {2{$random}};
    assign htif.io_scr_rdata_27 = {2{$random}};
    assign htif.io_scr_rdata_26 = {2{$random}};
    assign htif.io_scr_rdata_25 = {2{$random}};
    assign htif.io_scr_rdata_24 = {2{$random}};
    assign htif.io_scr_rdata_23 = {2{$random}};
    assign htif.io_scr_rdata_22 = {2{$random}};
    assign htif.io_scr_rdata_21 = {2{$random}};
    assign htif.io_scr_rdata_20 = {2{$random}};
    assign htif.io_scr_rdata_19 = {2{$random}};
    assign htif.io_scr_rdata_18 = {2{$random}};
    assign htif.io_scr_rdata_17 = {2{$random}};
    assign htif.io_scr_rdata_16 = {2{$random}};
    assign htif.io_scr_rdata_15 = {2{$random}};
    assign htif.io_scr_rdata_14 = {2{$random}};
    assign htif.io_scr_rdata_13 = {2{$random}};
    assign htif.io_scr_rdata_12 = {2{$random}};
    assign htif.io_scr_rdata_11 = {2{$random}};
    assign htif.io_scr_rdata_10 = {2{$random}};
    assign htif.io_scr_rdata_9 = {2{$random}};
    assign htif.io_scr_rdata_8 = {2{$random}};
    assign htif.io_scr_rdata_7 = {2{$random}};
    assign htif.io_scr_rdata_6 = {2{$random}};
    assign htif.io_scr_rdata_5 = {2{$random}};
    assign htif.io_scr_rdata_4 = {2{$random}};
    assign htif.io_scr_rdata_3 = {2{$random}};
    assign htif.io_scr_rdata_2 = {2{$random}};
  `endif
  OuterMemorySystem outmemsys(.clk(clk), .reset(reset),
       .io_tiles_0_acquire_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Queue_0_io_deq_valid ),
       .io_tiles_0_acquire_bits_header_src( Queue_0_io_deq_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Queue_0_io_deq_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Queue_0_io_deq_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Queue_0_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Queue_0_io_deq_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Queue_0_io_deq_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Queue_0_io_deq_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Queue_0_io_deq_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Queue_0_io_deq_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Queue_3_io_enq_ready ),
       .io_tiles_0_grant_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Queue_2_io_deq_valid ),
       .io_tiles_0_finish_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Queue_2_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Queue_4_io_enq_ready ),
       .io_tiles_0_probe_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( outmemsys_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Queue_1_io_deq_valid ),
       .io_tiles_0_release_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Queue_1_io_deq_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Queue_1_io_deq_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Queue_1_io_deq_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Queue_1_io_deq_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Queue_1_io_deq_bits_payload_r_type ),
       .io_htif_acquire_ready( outmemsys_io_htif_acquire_ready ),
       .io_htif_acquire_valid( Queue_5_io_deq_valid ),
       .io_htif_acquire_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_htif_acquire_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_htif_acquire_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_htif_acquire_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_htif_acquire_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_htif_acquire_bits_payload_a_type( Queue_5_io_deq_bits_payload_a_type ),
       .io_htif_acquire_bits_payload_write_mask( Queue_5_io_deq_bits_payload_write_mask ),
       .io_htif_acquire_bits_payload_subword_addr( Queue_5_io_deq_bits_payload_subword_addr ),
       .io_htif_acquire_bits_payload_atomic_opcode( Queue_5_io_deq_bits_payload_atomic_opcode ),
       .io_htif_grant_ready( Queue_8_io_enq_ready ),
       .io_htif_grant_valid( outmemsys_io_htif_grant_valid ),
       .io_htif_grant_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_htif_grant_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_htif_grant_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_htif_grant_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_htif_grant_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_htif_grant_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_htif_finish_ready( outmemsys_io_htif_finish_ready ),
       .io_htif_finish_valid( Queue_7_io_deq_valid ),
       .io_htif_finish_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_htif_finish_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_htif_finish_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id ),
       .io_htif_probe_ready( Queue_9_io_enq_ready ),
       .io_htif_probe_valid( outmemsys_io_htif_probe_valid ),
       .io_htif_probe_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_htif_probe_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_htif_probe_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_htif_probe_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_htif_probe_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_htif_release_ready( outmemsys_io_htif_release_ready ),
       .io_htif_release_valid( Queue_6_io_deq_valid ),
       .io_htif_release_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_htif_release_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_htif_release_bits_payload_addr( Queue_6_io_deq_bits_payload_addr ),
       .io_htif_release_bits_payload_client_xact_id( Queue_6_io_deq_bits_payload_client_xact_id ),
       .io_htif_release_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_htif_release_bits_payload_data( Queue_6_io_deq_bits_payload_data ),
       .io_htif_release_bits_payload_r_type( Queue_6_io_deq_bits_payload_r_type ),
       .io_incoherent_1( 1'h1 ),
       .io_incoherent_0( io_incoherent_0 ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( outmemsys_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( outmemsys_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( outmemsys_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( outmemsys_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( outmemsys_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( outmemsys_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  Queue_8 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( T43 ),
       .io_enq_bits_header_src( T42 ),
       .io_enq_bits_header_dst( T41 ),
       .io_enq_bits_payload_addr( T40 ),
       .io_enq_bits_payload_client_xact_id( T39 ),
       .io_enq_bits_payload_data( T38 ),
       .io_enq_bits_payload_a_type( T37 ),
       .io_enq_bits_payload_write_mask( T36 ),
       .io_enq_bits_payload_subword_addr( T35 ),
       .io_enq_bits_payload_atomic_opcode( T34 ),
       .io_deq_ready( outmemsys_io_tiles_0_acquire_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_header_src( Queue_0_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_0_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_0_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_0_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_0_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_0_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_0_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_0_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_0_io_deq_bits_payload_atomic_opcode )
  );
  Queue_9 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( T33 ),
       .io_enq_bits_header_src( T32 ),
       .io_enq_bits_header_dst( T31 ),
       .io_enq_bits_payload_addr( T30 ),
       .io_enq_bits_payload_client_xact_id( T29 ),
       .io_enq_bits_payload_master_xact_id( T28 ),
       .io_enq_bits_payload_data( T27 ),
       .io_enq_bits_payload_r_type( T26 ),
       .io_deq_ready( outmemsys_io_tiles_0_release_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits_header_src( Queue_1_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_1_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_1_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_1_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_1_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_1_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_1_io_deq_bits_payload_r_type )
  );
  Queue_10 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( T25 ),
       .io_enq_bits_header_src( T24 ),
       .io_enq_bits_header_dst( T23 ),
       .io_enq_bits_payload_master_xact_id( T22 ),
       .io_deq_ready( outmemsys_io_tiles_0_finish_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits_header_src( Queue_2_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_2_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_2_io_deq_bits_payload_master_xact_id )
  );
  Queue_11 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_tiles_0_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_tiles_0_grant_bits_payload_g_type ),
       .io_deq_ready( io_tiles_0_grant_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits_header_src( Queue_3_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_3_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_3_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_3_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_3_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_3_io_deq_bits_payload_g_type )
  );
  Queue_12 Queue_4(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_4_io_enq_ready ),
       .io_enq_valid( outmemsys_io_tiles_0_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_tiles_0_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_tiles_0_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_tiles_0_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_tiles_0_probe_bits_payload_p_type ),
       .io_deq_ready( io_tiles_0_probe_ready ),
       .io_deq_valid( Queue_4_io_deq_valid ),
       .io_deq_bits_header_src( Queue_4_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_4_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_4_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_4_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_4_io_deq_bits_payload_p_type )
  );
  Queue_8 Queue_5(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_5_io_enq_ready ),
       .io_enq_valid( T21 ),
       .io_enq_bits_header_src( T20 ),
       .io_enq_bits_header_dst( T19 ),
       .io_enq_bits_payload_addr( T18 ),
       .io_enq_bits_payload_client_xact_id( T17 ),
       .io_enq_bits_payload_data( T16 ),
       .io_enq_bits_payload_a_type( T15 ),
       .io_enq_bits_payload_write_mask( T14 ),
       .io_enq_bits_payload_subword_addr( T13 ),
       .io_enq_bits_payload_atomic_opcode( T12 ),
       .io_deq_ready( outmemsys_io_htif_acquire_ready ),
       .io_deq_valid( Queue_5_io_deq_valid ),
       .io_deq_bits_header_src( Queue_5_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_5_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_5_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_5_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_data( Queue_5_io_deq_bits_payload_data ),
       .io_deq_bits_payload_a_type( Queue_5_io_deq_bits_payload_a_type ),
       .io_deq_bits_payload_write_mask( Queue_5_io_deq_bits_payload_write_mask ),
       .io_deq_bits_payload_subword_addr( Queue_5_io_deq_bits_payload_subword_addr ),
       .io_deq_bits_payload_atomic_opcode( Queue_5_io_deq_bits_payload_atomic_opcode )
  );
  Queue_9 Queue_6(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_6_io_enq_ready ),
       .io_enq_valid( T11 ),
       .io_enq_bits_header_src( T10 ),
       .io_enq_bits_header_dst( T9 ),
       .io_enq_bits_payload_addr( T8 ),
       .io_enq_bits_payload_client_xact_id( T7 ),
       .io_enq_bits_payload_master_xact_id( T6 ),
       .io_enq_bits_payload_data( T5 ),
       .io_enq_bits_payload_r_type( T4 ),
       .io_deq_ready( outmemsys_io_htif_release_ready ),
       .io_deq_valid( Queue_6_io_deq_valid ),
       .io_deq_bits_header_src( Queue_6_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_6_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_6_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_client_xact_id( Queue_6_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_6_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_data( Queue_6_io_deq_bits_payload_data ),
       .io_deq_bits_payload_r_type( Queue_6_io_deq_bits_payload_r_type )
  );
  Queue_10 Queue_7(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_7_io_enq_ready ),
       .io_enq_valid( T3 ),
       .io_enq_bits_header_src( T2 ),
       .io_enq_bits_header_dst( T1 ),
       .io_enq_bits_payload_master_xact_id( T0 ),
       .io_deq_ready( outmemsys_io_htif_finish_ready ),
       .io_deq_valid( Queue_7_io_deq_valid ),
       .io_deq_bits_header_src( Queue_7_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_7_io_deq_bits_header_dst ),
       .io_deq_bits_payload_master_xact_id( Queue_7_io_deq_bits_payload_master_xact_id )
  );
  Queue_11 Queue_8(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_8_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_grant_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_grant_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_grant_bits_header_dst ),
       .io_enq_bits_payload_data( outmemsys_io_htif_grant_bits_payload_data ),
       .io_enq_bits_payload_client_xact_id( outmemsys_io_htif_grant_bits_payload_client_xact_id ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_grant_bits_payload_master_xact_id ),
       .io_enq_bits_payload_g_type( outmemsys_io_htif_grant_bits_payload_g_type ),
       .io_deq_ready( htif_io_mem_grant_ready ),
       .io_deq_valid( Queue_8_io_deq_valid ),
       .io_deq_bits_header_src( Queue_8_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_8_io_deq_bits_header_dst ),
       .io_deq_bits_payload_data( Queue_8_io_deq_bits_payload_data ),
       .io_deq_bits_payload_client_xact_id( Queue_8_io_deq_bits_payload_client_xact_id ),
       .io_deq_bits_payload_master_xact_id( Queue_8_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_g_type( Queue_8_io_deq_bits_payload_g_type )
  );
  Queue_12 Queue_9(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_9_io_enq_ready ),
       .io_enq_valid( outmemsys_io_htif_probe_valid ),
       .io_enq_bits_header_src( outmemsys_io_htif_probe_bits_header_src ),
       .io_enq_bits_header_dst( outmemsys_io_htif_probe_bits_header_dst ),
       .io_enq_bits_payload_addr( outmemsys_io_htif_probe_bits_payload_addr ),
       .io_enq_bits_payload_master_xact_id( outmemsys_io_htif_probe_bits_payload_master_xact_id ),
       .io_enq_bits_payload_p_type( outmemsys_io_htif_probe_bits_payload_p_type ),
       .io_deq_ready( htif_io_mem_probe_ready ),
       .io_deq_valid( Queue_9_io_deq_valid ),
       .io_deq_bits_header_src( Queue_9_io_deq_bits_header_src ),
       .io_deq_bits_header_dst( Queue_9_io_deq_bits_header_dst ),
       .io_deq_bits_payload_addr( Queue_9_io_deq_bits_payload_addr ),
       .io_deq_bits_payload_master_xact_id( Queue_9_io_deq_bits_payload_master_xact_id ),
       .io_deq_bits_payload_p_type( Queue_9_io_deq_bits_payload_p_type )
  );
endmodule

module Queue_13(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits_rw,
    input [4:0] io_enq_bits_addr,
    input [63:0] io_enq_bits_data,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits_rw,
    output[4:0] io_deq_bits_addr,
    output[63:0] io_deq_bits_data
);

  wire[63:0] T0;
  wire[69:0] T1;
  reg [69:0] ram [1:0];
  wire[69:0] T2;
  wire[69:0] T3;
  wire[69:0] T4;
  wire[68:0] T5;
  wire do_enq;
  reg  R6;
  wire T7;
  wire T8;
  wire T9;
  reg  R10;
  wire T11;
  wire T12;
  wire T13;
  wire do_deq;
  wire[4:0] T14;
  wire T15;
  wire T16;
  wire empty;
  wire T17;
  reg  maybe_full;
  wire T18;
  wire T19;
  wire T20;
  wire ptr_match;
  wire T21;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {3{$random}};
    R6 = {1{$random}};
    R10 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits_data = T0;
  assign T0 = T1[6'h3f:1'h0];
  assign T1 = ram[R10];
  assign T3 = T4;
  assign T4 = {io_enq_bits_rw, T5};
  assign T5 = {io_enq_bits_addr, io_enq_bits_data};
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_enq ? T9 : R6;
  assign T9 = R6 + 1'h1;
  assign T11 = reset ? 1'h0 : T12;
  assign T12 = do_deq ? T13 : R10;
  assign T13 = R10 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_bits_addr = T14;
  assign T14 = T1[7'h44:7'h40];
  assign io_deq_bits_rw = T15;
  assign T15 = T1[7'h45:7'h45];
  assign io_deq_valid = T16;
  assign T16 = empty ^ 1'h1;
  assign empty = ptr_match & T17;
  assign T17 = maybe_full ^ 1'h1;
  assign T18 = reset ? 1'h0 : T19;
  assign T19 = T20 ? do_enq : maybe_full;
  assign T20 = do_enq != do_deq;
  assign ptr_match = R6 == R10;
  assign io_enq_ready = T21;
  assign T21 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R6] <= T3;
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_enq) begin
      R6 <= T9;
    end
    if(reset) begin
      R10 <= 1'h0;
    end else if(do_deq) begin
      R10 <= T13;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T20) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_14(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [63:0] io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output[63:0] io_deq_bits
);

  wire[63:0] T0;
  reg [63:0] ram [1:0];
  wire[63:0] T1;
  wire do_enq;
  reg  R2;
  wire T3;
  wire T4;
  wire T5;
  reg  R6;
  wire T7;
  wire T8;
  wire T9;
  wire do_deq;
  wire T10;
  wire empty;
  wire T11;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire ptr_match;
  wire T15;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {2{$random}};
    R2 = {1{$random}};
    R6 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R6];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T3 = reset ? 1'h0 : T4;
  assign T4 = do_enq ? T5 : R2;
  assign T5 = R2 + 1'h1;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_deq ? T9 : R6;
  assign T9 = R6 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T10;
  assign T10 = empty ^ 1'h1;
  assign empty = ptr_match & T11;
  assign T11 = maybe_full ^ 1'h1;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign ptr_match = R2 == R6;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T5;
    end
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_deq) begin
      R6 <= T9;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Queue_15(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input  io_enq_bits,
    input  io_deq_ready,
    output io_deq_valid,
    output io_deq_bits
);

  wire T0;
  reg [0:0] ram [1:0];
  wire T1;
  wire do_enq;
  reg  R2;
  wire T3;
  wire T4;
  wire T5;
  reg  R6;
  wire T7;
  wire T8;
  wire T9;
  wire do_deq;
  wire T10;
  wire empty;
  wire T11;
  reg  maybe_full;
  wire T12;
  wire T13;
  wire T14;
  wire ptr_match;
  wire T15;
  wire full;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      ram[initvar] = {1{$random}};
    R2 = {1{$random}};
    R6 = {1{$random}};
    maybe_full = {1{$random}};
  end
`endif

  assign io_deq_bits = T0;
  assign T0 = ram[R6];
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T3 = reset ? 1'h0 : T4;
  assign T4 = do_enq ? T5 : R2;
  assign T5 = R2 + 1'h1;
  assign T7 = reset ? 1'h0 : T8;
  assign T8 = do_deq ? T9 : R6;
  assign T9 = R6 + 1'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign io_deq_valid = T10;
  assign T10 = empty ^ 1'h1;
  assign empty = ptr_match & T11;
  assign T11 = maybe_full ^ 1'h1;
  assign T12 = reset ? 1'h0 : T13;
  assign T13 = T14 ? do_enq : maybe_full;
  assign T14 = do_enq != do_deq;
  assign ptr_match = R2 == R6;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if (do_enq)
      ram[R2] <= io_enq_bits;
    if(reset) begin
      R2 <= 1'h0;
    end else if(do_enq) begin
      R2 <= T5;
    end
    if(reset) begin
      R6 <= 1'h0;
    end else if(do_deq) begin
      R6 <= T9;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T14) begin
      maybe_full <= do_enq;
    end
  end
endmodule

module Top(input clk, input reset,
    output io_host_clk,
    output io_host_clk_edge,
    output io_host_in_ready,
    input  io_host_in_valid,
    input [15:0] io_host_in_bits,
    input  io_host_out_ready,
    output io_host_out_valid,
    output[15:0] io_host_out_bits,
    output io_host_debug_stats_pcr,
    input  io_mem_req_cmd_ready,
    output io_mem_req_cmd_valid,
    output[25:0] io_mem_req_cmd_bits_addr,
    output[4:0] io_mem_req_cmd_bits_tag,
    output io_mem_req_cmd_bits_rw,
    input  io_mem_req_data_ready,
    output io_mem_req_data_valid,
    output[127:0] io_mem_req_data_bits_data,
    output io_mem_resp_ready,
    input  io_mem_resp_valid,
    input [127:0] io_mem_resp_bits_data,
    input [4:0] io_mem_resp_bits_tag,
    input  io_mem_backup_en,
    output io_in_mem_ready,
    input  io_in_mem_valid,
    input  io_out_mem_ready,
    output io_out_mem_valid
);

  wire resetSigs_0;
  wire uncore_io_htif_0_reset;
  wire Tile_io_host_ipi_rep_ready;
  wire uncore_io_htif_0_ipi_rep_bits;
  wire uncore_io_htif_0_ipi_rep_valid;
  wire uncore_io_htif_0_ipi_req_ready;
  wire Tile_io_host_ipi_req_bits;
  wire Tile_io_host_ipi_req_valid;
  wire uncore_io_htif_0_pcr_rep_ready;
  wire[63:0] Tile_io_host_pcr_rep_bits;
  wire Tile_io_host_pcr_rep_valid;
  wire Tile_io_host_pcr_req_ready;
  wire[63:0] uncore_io_htif_0_pcr_req_bits_data;
  wire[4:0] uncore_io_htif_0_pcr_req_bits_addr;
  wire uncore_io_htif_0_pcr_req_bits_rw;
  wire uncore_io_htif_0_pcr_req_valid;
  wire Tile_io_host_debug_stats_pcr;
  wire Queue_3_io_enq_ready;
  wire Queue_2_io_deq_bits;
  wire Queue_2_io_deq_valid;
  wire[63:0] Queue_1_io_deq_bits;
  wire Queue_1_io_deq_valid;
  wire Queue_0_io_enq_ready;
  wire[2:0] Tile_io_tilelink_release_bits_payload_r_type;
  wire[511:0] Tile_io_tilelink_release_bits_payload_data;
  wire[2:0] Tile_io_tilelink_release_bits_payload_master_xact_id;
  wire[1:0] Tile_io_tilelink_release_bits_payload_client_xact_id;
  wire[25:0] Tile_io_tilelink_release_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_release_bits_header_dst;
  wire[1:0] Tile_io_tilelink_release_bits_header_src;
  wire Tile_io_tilelink_release_valid;
  wire Tile_io_tilelink_probe_ready;
  wire[2:0] Tile_io_tilelink_finish_bits_payload_master_xact_id;
  wire[1:0] Tile_io_tilelink_finish_bits_header_dst;
  wire[1:0] Tile_io_tilelink_finish_bits_header_src;
  wire Tile_io_tilelink_finish_valid;
  wire Tile_io_tilelink_grant_ready;
  wire[3:0] Tile_io_tilelink_acquire_bits_payload_atomic_opcode;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_subword_addr;
  wire[5:0] Tile_io_tilelink_acquire_bits_payload_write_mask;
  wire[2:0] Tile_io_tilelink_acquire_bits_payload_a_type;
  wire[511:0] Tile_io_tilelink_acquire_bits_payload_data;
  wire[1:0] Tile_io_tilelink_acquire_bits_payload_client_xact_id;
  wire[25:0] Tile_io_tilelink_acquire_bits_payload_addr;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_dst;
  wire[1:0] Tile_io_tilelink_acquire_bits_header_src;
  wire Tile_io_tilelink_acquire_valid;
  wire Queue_3_io_deq_bits;
  wire Queue_3_io_deq_valid;
  wire Queue_2_io_enq_ready;
  wire Queue_1_io_enq_ready;
  wire[63:0] Queue_0_io_deq_bits_data;
  wire[4:0] Queue_0_io_deq_bits_addr;
  wire Queue_0_io_deq_bits_rw;
  wire Queue_0_io_deq_valid;
  reg  R0;
  reg  R1;
  wire uncore_io_tiles_0_release_ready;
  wire[1:0] uncore_io_tiles_0_probe_bits_payload_p_type;
  wire[2:0] uncore_io_tiles_0_probe_bits_payload_master_xact_id;
  wire[25:0] uncore_io_tiles_0_probe_bits_payload_addr;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_dst;
  wire[1:0] uncore_io_tiles_0_probe_bits_header_src;
  wire uncore_io_tiles_0_probe_valid;
  wire uncore_io_tiles_0_finish_ready;
  wire[3:0] uncore_io_tiles_0_grant_bits_payload_g_type;
  wire[2:0] uncore_io_tiles_0_grant_bits_payload_master_xact_id;
  wire[1:0] uncore_io_tiles_0_grant_bits_payload_client_xact_id;
  wire[511:0] uncore_io_tiles_0_grant_bits_payload_data;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_dst;
  wire[1:0] uncore_io_tiles_0_grant_bits_header_src;
  wire uncore_io_tiles_0_grant_valid;
  wire uncore_io_tiles_0_acquire_ready;
  wire[127:0] uncore_io_mem_req_data_bits_data;
  wire uncore_io_mem_req_data_valid;
  wire uncore_io_mem_req_cmd_bits_rw;
  wire[4:0] uncore_io_mem_req_cmd_bits_tag;
  wire[25:0] uncore_io_mem_req_cmd_bits_addr;
  wire uncore_io_mem_req_cmd_valid;
  wire uncore_io_host_debug_stats_pcr;
  wire[15:0] uncore_io_host_out_bits;
  wire uncore_io_host_out_valid;
  wire uncore_io_host_in_ready;

`ifndef SYNTHESIS
  integer initvar;
  initial begin
    #0.002;
    R0 = {1{$random}};
    R1 = {1{$random}};
  end
`endif

  assign resetSigs_0 = uncore_io_htif_0_reset;
  assign io_mem_req_data_bits_data = uncore_io_mem_req_data_bits_data;
  assign io_mem_req_data_valid = uncore_io_mem_req_data_valid;
  assign io_mem_req_cmd_bits_rw = uncore_io_mem_req_cmd_bits_rw;
  assign io_mem_req_cmd_bits_tag = uncore_io_mem_req_cmd_bits_tag;
  assign io_mem_req_cmd_bits_addr = uncore_io_mem_req_cmd_bits_addr;
  assign io_mem_req_cmd_valid = uncore_io_mem_req_cmd_valid;
  assign io_host_debug_stats_pcr = uncore_io_host_debug_stats_pcr;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_in_ready = uncore_io_host_in_ready;
  Tile Tile(.clk(clk), .reset(resetSigs_0),
       .io_tilelink_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tilelink_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tilelink_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tilelink_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tilelink_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tilelink_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tilelink_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tilelink_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tilelink_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tilelink_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tilelink_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tilelink_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tilelink_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tilelink_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tilelink_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tilelink_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tilelink_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tilelink_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tilelink_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tilelink_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tilelink_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tilelink_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tilelink_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tilelink_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tilelink_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tilelink_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tilelink_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tilelink_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tilelink_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tilelink_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tilelink_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tilelink_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tilelink_release_valid( Tile_io_tilelink_release_valid ),
       .io_tilelink_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tilelink_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tilelink_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tilelink_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tilelink_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tilelink_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tilelink_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_host_reset( R0 ),
       .io_host_id( 1'h0 ),
       .io_host_pcr_req_ready( Tile_io_host_pcr_req_ready ),
       .io_host_pcr_req_valid( Queue_0_io_deq_valid ),
       .io_host_pcr_req_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_host_pcr_req_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_host_pcr_req_bits_data( Queue_0_io_deq_bits_data ),
       .io_host_pcr_rep_ready( Queue_1_io_enq_ready ),
       .io_host_pcr_rep_valid( Tile_io_host_pcr_rep_valid ),
       .io_host_pcr_rep_bits( Tile_io_host_pcr_rep_bits ),
       .io_host_ipi_req_ready( Queue_2_io_enq_ready ),
       .io_host_ipi_req_valid( Tile_io_host_ipi_req_valid ),
       .io_host_ipi_req_bits( Tile_io_host_ipi_req_bits ),
       .io_host_ipi_rep_ready( Tile_io_host_ipi_rep_ready ),
       .io_host_ipi_rep_valid( Queue_3_io_deq_valid ),
       .io_host_ipi_rep_bits( Queue_3_io_deq_bits ),
       .io_host_debug_stats_pcr( Tile_io_host_debug_stats_pcr )
  );
  Uncore uncore(.clk(clk), .reset(reset),
       //.io_host_clk(  )
       //.io_host_clk_edge(  )
       .io_host_in_ready( uncore_io_host_in_ready ),
       .io_host_in_valid( io_host_in_valid ),
       .io_host_in_bits( io_host_in_bits ),
       .io_host_out_ready( io_host_out_ready ),
       .io_host_out_valid( uncore_io_host_out_valid ),
       .io_host_out_bits( uncore_io_host_out_bits ),
       .io_host_debug_stats_pcr( uncore_io_host_debug_stats_pcr ),
       .io_mem_req_cmd_ready( io_mem_req_cmd_ready ),
       .io_mem_req_cmd_valid( uncore_io_mem_req_cmd_valid ),
       .io_mem_req_cmd_bits_addr( uncore_io_mem_req_cmd_bits_addr ),
       .io_mem_req_cmd_bits_tag( uncore_io_mem_req_cmd_bits_tag ),
       .io_mem_req_cmd_bits_rw( uncore_io_mem_req_cmd_bits_rw ),
       .io_mem_req_data_ready( io_mem_req_data_ready ),
       .io_mem_req_data_valid( uncore_io_mem_req_data_valid ),
       .io_mem_req_data_bits_data( uncore_io_mem_req_data_bits_data ),
       //.io_mem_resp_ready(  )
       .io_mem_resp_valid( io_mem_resp_valid ),
       .io_mem_resp_bits_data( io_mem_resp_bits_data ),
       .io_mem_resp_bits_tag( io_mem_resp_bits_tag ),
       .io_tiles_0_acquire_ready( uncore_io_tiles_0_acquire_ready ),
       .io_tiles_0_acquire_valid( Tile_io_tilelink_acquire_valid ),
       .io_tiles_0_acquire_bits_header_src( Tile_io_tilelink_acquire_bits_header_src ),
       .io_tiles_0_acquire_bits_header_dst( Tile_io_tilelink_acquire_bits_header_dst ),
       .io_tiles_0_acquire_bits_payload_addr( Tile_io_tilelink_acquire_bits_payload_addr ),
       .io_tiles_0_acquire_bits_payload_client_xact_id( Tile_io_tilelink_acquire_bits_payload_client_xact_id ),
       .io_tiles_0_acquire_bits_payload_data( Tile_io_tilelink_acquire_bits_payload_data ),
       .io_tiles_0_acquire_bits_payload_a_type( Tile_io_tilelink_acquire_bits_payload_a_type ),
       .io_tiles_0_acquire_bits_payload_write_mask( Tile_io_tilelink_acquire_bits_payload_write_mask ),
       .io_tiles_0_acquire_bits_payload_subword_addr( Tile_io_tilelink_acquire_bits_payload_subword_addr ),
       .io_tiles_0_acquire_bits_payload_atomic_opcode( Tile_io_tilelink_acquire_bits_payload_atomic_opcode ),
       .io_tiles_0_grant_ready( Tile_io_tilelink_grant_ready ),
       .io_tiles_0_grant_valid( uncore_io_tiles_0_grant_valid ),
       .io_tiles_0_grant_bits_header_src( uncore_io_tiles_0_grant_bits_header_src ),
       .io_tiles_0_grant_bits_header_dst( uncore_io_tiles_0_grant_bits_header_dst ),
       .io_tiles_0_grant_bits_payload_data( uncore_io_tiles_0_grant_bits_payload_data ),
       .io_tiles_0_grant_bits_payload_client_xact_id( uncore_io_tiles_0_grant_bits_payload_client_xact_id ),
       .io_tiles_0_grant_bits_payload_master_xact_id( uncore_io_tiles_0_grant_bits_payload_master_xact_id ),
       .io_tiles_0_grant_bits_payload_g_type( uncore_io_tiles_0_grant_bits_payload_g_type ),
       .io_tiles_0_finish_ready( uncore_io_tiles_0_finish_ready ),
       .io_tiles_0_finish_valid( Tile_io_tilelink_finish_valid ),
       .io_tiles_0_finish_bits_header_src( Tile_io_tilelink_finish_bits_header_src ),
       .io_tiles_0_finish_bits_header_dst( Tile_io_tilelink_finish_bits_header_dst ),
       .io_tiles_0_finish_bits_payload_master_xact_id( Tile_io_tilelink_finish_bits_payload_master_xact_id ),
       .io_tiles_0_probe_ready( Tile_io_tilelink_probe_ready ),
       .io_tiles_0_probe_valid( uncore_io_tiles_0_probe_valid ),
       .io_tiles_0_probe_bits_header_src( uncore_io_tiles_0_probe_bits_header_src ),
       .io_tiles_0_probe_bits_header_dst( uncore_io_tiles_0_probe_bits_header_dst ),
       .io_tiles_0_probe_bits_payload_addr( uncore_io_tiles_0_probe_bits_payload_addr ),
       .io_tiles_0_probe_bits_payload_master_xact_id( uncore_io_tiles_0_probe_bits_payload_master_xact_id ),
       .io_tiles_0_probe_bits_payload_p_type( uncore_io_tiles_0_probe_bits_payload_p_type ),
       .io_tiles_0_release_ready( uncore_io_tiles_0_release_ready ),
       .io_tiles_0_release_valid( Tile_io_tilelink_release_valid ),
       .io_tiles_0_release_bits_header_src( Tile_io_tilelink_release_bits_header_src ),
       .io_tiles_0_release_bits_header_dst( Tile_io_tilelink_release_bits_header_dst ),
       .io_tiles_0_release_bits_payload_addr( Tile_io_tilelink_release_bits_payload_addr ),
       .io_tiles_0_release_bits_payload_client_xact_id( Tile_io_tilelink_release_bits_payload_client_xact_id ),
       .io_tiles_0_release_bits_payload_master_xact_id( Tile_io_tilelink_release_bits_payload_master_xact_id ),
       .io_tiles_0_release_bits_payload_data( Tile_io_tilelink_release_bits_payload_data ),
       .io_tiles_0_release_bits_payload_r_type( Tile_io_tilelink_release_bits_payload_r_type ),
       .io_htif_0_reset( uncore_io_htif_0_reset ),
       //.io_htif_0_id(  )
       .io_htif_0_pcr_req_ready( Queue_0_io_enq_ready ),
       .io_htif_0_pcr_req_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_htif_0_pcr_req_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_htif_0_pcr_req_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_htif_0_pcr_req_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_htif_0_pcr_rep_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_htif_0_pcr_rep_valid( Queue_1_io_deq_valid ),
       .io_htif_0_pcr_rep_bits( Queue_1_io_deq_bits ),
       .io_htif_0_ipi_req_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_htif_0_ipi_req_valid( Queue_2_io_deq_valid ),
       .io_htif_0_ipi_req_bits( Queue_2_io_deq_bits ),
       .io_htif_0_ipi_rep_ready( Queue_3_io_enq_ready ),
       .io_htif_0_ipi_rep_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_htif_0_ipi_rep_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_htif_0_debug_stats_pcr( Tile_io_host_debug_stats_pcr ),
       .io_incoherent_0( uncore_io_htif_0_reset )
       //.io_mem_backup_req_ready(  )
       //.io_mem_backup_req_valid(  )
       //.io_mem_backup_req_bits(  )
       //.io_mem_backup_resp_valid(  )
       //.io_mem_backup_resp_bits(  )
       //.io_mem_backup_en(  )
  );
  `ifndef SYNTHESIS
    assign uncore.io_htif_0_ipi_rep_bits = {1{$random}};
  `endif
  Queue_13 Queue_0(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_0_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_pcr_req_valid ),
       .io_enq_bits_rw( uncore_io_htif_0_pcr_req_bits_rw ),
       .io_enq_bits_addr( uncore_io_htif_0_pcr_req_bits_addr ),
       .io_enq_bits_data( uncore_io_htif_0_pcr_req_bits_data ),
       .io_deq_ready( Tile_io_host_pcr_req_ready ),
       .io_deq_valid( Queue_0_io_deq_valid ),
       .io_deq_bits_rw( Queue_0_io_deq_bits_rw ),
       .io_deq_bits_addr( Queue_0_io_deq_bits_addr ),
       .io_deq_bits_data( Queue_0_io_deq_bits_data )
  );
  Queue_14 Queue_1(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_1_io_enq_ready ),
       .io_enq_valid( Tile_io_host_pcr_rep_valid ),
       .io_enq_bits( Tile_io_host_pcr_rep_bits ),
       .io_deq_ready( uncore_io_htif_0_pcr_rep_ready ),
       .io_deq_valid( Queue_1_io_deq_valid ),
       .io_deq_bits( Queue_1_io_deq_bits )
  );
  Queue_15 Queue_2(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_2_io_enq_ready ),
       .io_enq_valid( Tile_io_host_ipi_req_valid ),
       .io_enq_bits( Tile_io_host_ipi_req_bits ),
       .io_deq_ready( uncore_io_htif_0_ipi_req_ready ),
       .io_deq_valid( Queue_2_io_deq_valid ),
       .io_deq_bits( Queue_2_io_deq_bits )
  );
  Queue_15 Queue_3(.clk(clk), .reset(reset),
       .io_enq_ready( Queue_3_io_enq_ready ),
       .io_enq_valid( uncore_io_htif_0_ipi_rep_valid ),
       .io_enq_bits( uncore_io_htif_0_ipi_rep_bits ),
       .io_deq_ready( Tile_io_host_ipi_rep_ready ),
       .io_deq_valid( Queue_3_io_deq_valid ),
       .io_deq_bits( Queue_3_io_deq_bits )
  );

  always @(posedge clk) begin
    R0 <= R1;
    R1 <= uncore_io_htif_0_reset;
  end
endmodule

module DataArray_T2(
  input CLK,
  input RST,
  input init,
  input [7:0] W0A,
  input W0E,
  input [127:0] W0I,
  input [127:0] W0M,
  input [7:0] R1A,
  input R1E,
  output [127:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<2; i=i+64) begin
    for (j=1; j<64; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][63:0] <= W0I[63:0];
  if (W0E && W0M[64]) ram[W0A][127:64] <= W0I[127:64];
end
assign R1O = ram[reg_R1A];

endmodule


module MetadataArray_tag_arr(
  input CLK,
  input RST,
  input init,
  input [5:0] W0A,
  input W0E,
  input [21:0] W0I,
  input [21:0] W0M,
  input [5:0] R1A,
  input R1E,
  output [21:0] R1O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+22) begin
    for (j=1; j<22; j=j+1) begin
      if (W0M[i] != W0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [21:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_R1A;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
  if (W0E && W0M[0]) ram[W0A][21:0] <= W0I[21:0];
end
assign R1O = ram[reg_R1A];

endmodule


module ICache_tag_array(
  input CLK,
  input RST,
  input init,
  input [5:0] RW0A,
  input RW0E,
  input RW0W,
  input [19:0] RW0M,
  input [19:0] RW0I,
  output [19:0] RW0O
);

`ifndef SYNTHESIS
integer i;
integer j;
always @(posedge CLK) begin
  for (i=0; i<1; i=i+20) begin
    for (j=1; j<20; j=j+1) begin
      if (RW0M[i] != RW0M[i+j]) begin
        $fwrite(32'h80000002, "ASSERTION FAILED: write mask granularity\n");
        $finish;
      end
    end
  end
end
`endif

reg [19:0] ram [63:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 64; initvar = initvar+1)
        ram[initvar] = {1 {$random}};
    end
  `endif
  reg [5:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W && RW0M[0]) ram[RW0A][19:0] <= RW0I[19:0];
end
assign RW0O = ram[reg_RW0A];

endmodule


module ICache_T121(
  input CLK,
  input RST,
  input init,
  input [7:0] RW0A,
  input RW0E,
  input RW0W,
  input [127:0] RW0I,
  output [127:0] RW0O
);

reg [127:0] ram [255:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 256; initvar = initvar+1)
        ram[initvar] = {4 {$random}};
    end
  `endif
  reg [7:0] reg_RW0A;
always @(posedge CLK) begin
  if (RW0E && !RW0W) reg_RW0A <= RW0A;
  if (RW0E && RW0W) ram[RW0A] <= RW0I;
end
assign RW0O = ram[reg_RW0A];

endmodule


module HellaFlowQueue_ram(
  input CLK,
  input RST,
  input init,
  input [4:0] W0A,
  input W0E,
  input [132:0] W0I,
  input [4:0] R1A,
  input R1E,
  output [132:0] R1O
);

reg [132:0] ram [31:0];
  `ifndef SYNTHESIS
    integer initvar;
    initial begin
      #0.002;
      for (initvar = 0; initvar < 32; initvar = initvar+1)
        ram[initvar] = {5 {$random}};
    end
  `endif
  reg [4:0] reg_R1A;
  reg [4:0] latch_W0A;
  reg [132:0] latch_W0I;
  reg latch_W0E;
always @(posedge CLK) begin
  if (R1E) reg_R1A <= R1A;
end
assign R1O = ram[reg_R1A];
  always @(*) begin
    if (!CLK && W0E) latch_W0A <= W0A;
    if (!CLK && W0E) latch_W0I <= W0I;
    if (!CLK) latch_W0E <= W0E;
  end
  always @(*)
    if (CLK && latch_W0E)
      ram[latch_W0A] <= latch_W0I;

endmodule


